
library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

package CONV_PACK_rmedt_square is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_rmedt_square;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_inc_3 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_0_DW01_inc_3;

architecture SYN_cla of KSA_0_DW01_inc_3 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U2 : XOR2X1 port map( A => n3, B => A(6), Y => SUM(6));
   U3 : XOR2X1 port map( A => n5, B => A(4), Y => SUM(4));
   U4 : AND2X2 port map( A => A(1), B => A(0), Y => n1);
   U5 : XOR2X1 port map( A => n1, B => A(2), Y => SUM(2));
   U6 : XNOR2X1 port map( A => A(7), B => n2, Y => SUM(7));
   U7 : NAND2X1 port map( A => A(6), B => n3, Y => n2);
   U8 : INVX2 port map( A => n4, Y => n3);
   U9 : NAND3X1 port map( A => A(4), B => A(5), C => n5, Y => n4);
   U10 : XNOR2X1 port map( A => A(5), B => n6, Y => SUM(5));
   U11 : NAND2X1 port map( A => A(4), B => n5, Y => n6);
   U12 : INVX2 port map( A => n7, Y => n5);
   U13 : NAND3X1 port map( A => A(2), B => A(3), C => n1, Y => n7);
   U14 : XNOR2X1 port map( A => A(3), B => n8, Y => SUM(3));
   U15 : NAND2X1 port map( A => A(2), B => n1, Y => n8);
   U16 : XOR2X1 port map( A => A(1), B => A(0), Y => SUM(1));
   U17 : INVX2 port map( A => A(0), Y => SUM(0));

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_add_9 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_0_DW01_add_9;

architecture SYN_cla of KSA_0_DW01_add_9 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59 : 
      std_logic;

begin
   
   U2 : INVX2 port map( A => n17, Y => n1);
   U3 : INVX1 port map( A => n5, Y => n21);
   U4 : AND2X2 port map( A => n27, B => n11, Y => n2);
   U5 : NAND2X1 port map( A => n3, B => n37, Y => n15);
   U6 : AND2X2 port map( A => n38, B => n39, Y => n3);
   U7 : AND2X2 port map( A => B(0), B => A(0), Y => n4);
   U8 : OAI21X1 port map( A => B(6), B => A(6), C => n11, Y => n5);
   U9 : OR2X2 port map( A => A(6), B => B(6), Y => n12);
   U10 : INVX2 port map( A => n37, Y => n34);
   U11 : INVX2 port map( A => n59, Y => SUM(0));
   U12 : XOR2X1 port map( A => n6, B => n7, Y => SUM(7));
   U13 : XOR2X1 port map( A => B(7), B => A(7), Y => n7);
   U14 : NAND3X1 port map( A => n8, B => n9, C => n10, Y => n6);
   U15 : NAND3X1 port map( A => n11, B => n12, C => n13, Y => n10);
   U16 : NAND3X1 port map( A => n14, B => n11, C => n15, Y => n9);
   U17 : AOI21X1 port map( A => n16, B => n17, C => n18, Y => n14);
   U18 : NAND2X1 port map( A => n19, B => n20, Y => n18);
   U19 : INVX2 port map( A => B(6), Y => n17);
   U20 : INVX2 port map( A => A(6), Y => n16);
   U21 : AOI21X1 port map( A => n21, B => n22, C => n23, Y => n8);
   U22 : NAND2X1 port map( A => n24, B => n25, Y => n23);
   U23 : OAI21X1 port map( A => A(6), B => B(6), C => n26, Y => n25);
   U24 : INVX2 port map( A => n27, Y => n26);
   U25 : XOR2X1 port map( A => n28, B => n29, Y => SUM(6));
   U26 : INVX2 port map( A => n30, Y => n29);
   U27 : OAI21X1 port map( A => n1, B => A(6), C => n24, Y => n30);
   U28 : NAND2X1 port map( A => B(6), B => A(6), Y => n24);
   U29 : NAND3X1 port map( A => n27, B => n31, C => n32, Y => n28);
   U30 : OAI21X1 port map( A => n33, B => n34, C => n35, Y => n32);
   U31 : AND2X2 port map( A => n36, B => n11, Y => n35);
   U32 : NAND2X1 port map( A => n38, B => n39, Y => n33);
   U33 : AOI22X1 port map( A => n22, B => n11, C => n13, D => n11, Y => n31);
   U34 : INVX2 port map( A => n40, Y => n13);
   U35 : INVX2 port map( A => n41, Y => n22);
   U36 : XNOR2X1 port map( A => n42, B => n2, Y => SUM(5));
   U37 : OR2X2 port map( A => A(5), B => B(5), Y => n11);
   U38 : NAND2X1 port map( A => B(5), B => A(5), Y => n27);
   U39 : AOI21X1 port map( A => n36, B => n15, C => n43, Y => n42);
   U40 : NAND2X1 port map( A => n40, B => n41, Y => n43);
   U41 : NAND3X1 port map( A => A(3), B => B(3), C => n19, Y => n40);
   U42 : INVX2 port map( A => n44, Y => n36);
   U43 : OAI21X1 port map( A => A(4), B => B(4), C => n20, Y => n44);
   U44 : XNOR2X1 port map( A => n45, B => n46, Y => SUM(4));
   U45 : AND2X2 port map( A => n19, B => n41, Y => n46);
   U46 : NAND2X1 port map( A => B(4), B => A(4), Y => n41);
   U47 : OR2X2 port map( A => A(4), B => B(4), Y => n19);
   U48 : AOI21X1 port map( A => n15, B => n20, C => n47, Y => n45);
   U49 : INVX2 port map( A => n48, Y => n47);
   U50 : XNOR2X1 port map( A => n15, B => n49, Y => SUM(3));
   U51 : NAND2X1 port map( A => n20, B => n48, Y => n49);
   U52 : NAND2X1 port map( A => B(3), B => A(3), Y => n48);
   U53 : OR2X2 port map( A => A(3), B => B(3), Y => n20);
   U54 : NAND3X1 port map( A => n50, B => n51, C => n52, Y => n37);
   U55 : AND2X2 port map( A => B(0), B => A(0), Y => n52);
   U56 : NAND3X1 port map( A => A(1), B => B(1), C => n51, Y => n38);
   U57 : XOR2X1 port map( A => n53, B => n54, Y => SUM(2));
   U58 : AOI21X1 port map( A => n4, B => n50, C => n55, Y => n54);
   U59 : INVX2 port map( A => n56, Y => n55);
   U60 : NAND2X1 port map( A => n51, B => n39, Y => n53);
   U61 : NAND2X1 port map( A => B(2), B => A(2), Y => n39);
   U62 : OR2X2 port map( A => A(2), B => B(2), Y => n51);
   U63 : XNOR2X1 port map( A => n57, B => n4, Y => SUM(1));
   U64 : NAND2X1 port map( A => n50, B => n56, Y => n57);
   U65 : NAND2X1 port map( A => B(1), B => A(1), Y => n56);
   U66 : OR2X2 port map( A => A(1), B => B(1), Y => n50);
   U67 : OAI21X1 port map( A => A(0), B => B(0), C => n58, Y => n59);
   U68 : NAND2X1 port map( A => B(0), B => A(0), Y => n58);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_inc_3 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_1_DW01_inc_3;

architecture SYN_cla of KSA_1_DW01_inc_3 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U2 : XOR2X1 port map( A => n5, B => A(4), Y => SUM(4));
   U3 : XOR2X1 port map( A => n1, B => A(2), Y => SUM(2));
   U4 : XOR2X1 port map( A => n3, B => A(6), Y => SUM(6));
   U5 : AND2X2 port map( A => A(1), B => A(0), Y => n1);
   U6 : XNOR2X1 port map( A => A(7), B => n2, Y => SUM(7));
   U7 : NAND2X1 port map( A => A(6), B => n3, Y => n2);
   U8 : INVX2 port map( A => n4, Y => n3);
   U9 : NAND3X1 port map( A => A(4), B => A(5), C => n5, Y => n4);
   U10 : XNOR2X1 port map( A => A(5), B => n6, Y => SUM(5));
   U11 : NAND2X1 port map( A => A(4), B => n5, Y => n6);
   U12 : INVX2 port map( A => n7, Y => n5);
   U13 : NAND3X1 port map( A => A(2), B => A(3), C => n1, Y => n7);
   U14 : XNOR2X1 port map( A => A(3), B => n8, Y => SUM(3));
   U15 : NAND2X1 port map( A => A(2), B => n1, Y => n8);
   U16 : XOR2X1 port map( A => A(1), B => A(0), Y => SUM(1));
   U17 : INVX2 port map( A => A(0), Y => SUM(0));

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_add_9 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_1_DW01_add_9;

architecture SYN_cla of KSA_1_DW01_add_9 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61 : std_logic;

begin
   
   U2 : NAND2X1 port map( A => n5, B => n39, Y => n1);
   U3 : NAND2X1 port map( A => n5, B => n39, Y => n2);
   U4 : INVX1 port map( A => n19, Y => n3);
   U5 : INVX1 port map( A => B(6), Y => n19);
   U6 : INVX1 port map( A => n7, Y => n23);
   U7 : AND2X2 port map( A => n29, B => n13, Y => n4);
   U8 : NAND2X1 port map( A => n5, B => n39, Y => n17);
   U9 : AND2X2 port map( A => n40, B => n41, Y => n5);
   U10 : AND2X2 port map( A => B(0), B => A(0), Y => n6);
   U11 : OAI21X1 port map( A => B(6), B => A(6), C => n13, Y => n7);
   U12 : OR2X2 port map( A => B(6), B => A(6), Y => n14);
   U13 : INVX2 port map( A => n39, Y => n36);
   U14 : INVX2 port map( A => n61, Y => SUM(0));
   U15 : XOR2X1 port map( A => n8, B => n9, Y => SUM(7));
   U16 : XOR2X1 port map( A => B(7), B => A(7), Y => n9);
   U17 : NAND3X1 port map( A => n10, B => n11, C => n12, Y => n8);
   U18 : NAND3X1 port map( A => n13, B => n14, C => n15, Y => n12);
   U19 : NAND3X1 port map( A => n16, B => n13, C => n17, Y => n11);
   U20 : AOI21X1 port map( A => n18, B => n19, C => n20, Y => n16);
   U21 : NAND2X1 port map( A => n21, B => n22, Y => n20);
   U22 : INVX2 port map( A => A(6), Y => n18);
   U23 : AOI21X1 port map( A => n23, B => n24, C => n25, Y => n10);
   U24 : NAND2X1 port map( A => n26, B => n27, Y => n25);
   U25 : OAI21X1 port map( A => A(6), B => B(6), C => n28, Y => n27);
   U26 : INVX2 port map( A => n29, Y => n28);
   U27 : XOR2X1 port map( A => n30, B => n31, Y => SUM(6));
   U28 : INVX2 port map( A => n32, Y => n31);
   U29 : OAI21X1 port map( A => n3, B => A(6), C => n26, Y => n32);
   U30 : NAND2X1 port map( A => B(6), B => A(6), Y => n26);
   U31 : NAND3X1 port map( A => n29, B => n33, C => n34, Y => n30);
   U32 : OAI21X1 port map( A => n35, B => n36, C => n37, Y => n34);
   U33 : AND2X2 port map( A => n38, B => n13, Y => n37);
   U34 : NAND2X1 port map( A => n40, B => n41, Y => n35);
   U35 : AOI22X1 port map( A => n24, B => n13, C => n15, D => n13, Y => n33);
   U36 : INVX2 port map( A => n42, Y => n15);
   U37 : INVX2 port map( A => n43, Y => n24);
   U38 : XNOR2X1 port map( A => n44, B => n4, Y => SUM(5));
   U39 : OR2X2 port map( A => A(5), B => B(5), Y => n13);
   U40 : NAND2X1 port map( A => B(5), B => A(5), Y => n29);
   U41 : AOI21X1 port map( A => n38, B => n1, C => n45, Y => n44);
   U42 : NAND2X1 port map( A => n42, B => n43, Y => n45);
   U43 : NAND3X1 port map( A => A(3), B => B(3), C => n21, Y => n42);
   U44 : INVX2 port map( A => n46, Y => n38);
   U45 : OAI21X1 port map( A => A(4), B => B(4), C => n22, Y => n46);
   U46 : XNOR2X1 port map( A => n47, B => n48, Y => SUM(4));
   U47 : AND2X2 port map( A => n21, B => n43, Y => n48);
   U48 : NAND2X1 port map( A => B(4), B => A(4), Y => n43);
   U49 : OR2X2 port map( A => A(4), B => B(4), Y => n21);
   U50 : AOI21X1 port map( A => n2, B => n22, C => n49, Y => n47);
   U51 : INVX2 port map( A => n50, Y => n49);
   U52 : XNOR2X1 port map( A => n17, B => n51, Y => SUM(3));
   U53 : NAND2X1 port map( A => n22, B => n50, Y => n51);
   U54 : NAND2X1 port map( A => B(3), B => A(3), Y => n50);
   U55 : OR2X2 port map( A => A(3), B => B(3), Y => n22);
   U56 : NAND3X1 port map( A => n52, B => n53, C => n54, Y => n39);
   U57 : AND2X2 port map( A => B(0), B => A(0), Y => n54);
   U58 : NAND3X1 port map( A => A(1), B => B(1), C => n53, Y => n40);
   U59 : XOR2X1 port map( A => n55, B => n56, Y => SUM(2));
   U60 : AOI21X1 port map( A => n6, B => n52, C => n57, Y => n56);
   U61 : INVX2 port map( A => n58, Y => n57);
   U62 : NAND2X1 port map( A => n53, B => n41, Y => n55);
   U63 : NAND2X1 port map( A => B(2), B => A(2), Y => n41);
   U64 : OR2X2 port map( A => A(2), B => B(2), Y => n53);
   U65 : XNOR2X1 port map( A => n59, B => n6, Y => SUM(1));
   U66 : NAND2X1 port map( A => n52, B => n58, Y => n59);
   U67 : NAND2X1 port map( A => B(1), B => A(1), Y => n58);
   U68 : OR2X2 port map( A => A(1), B => B(1), Y => n52);
   U69 : OAI21X1 port map( A => A(0), B => B(0), C => n60, Y => n61);
   U70 : NAND2X1 port map( A => B(0), B => A(0), Y => n60);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_add_8 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_0_DW01_add_8;

architecture SYN_cla of KSA_0_DW01_add_8 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49 : std_logic;

begin
   
   U2 : OAI21X1 port map( A => n17, B => n18, C => n19, Y => n1);
   U3 : XNOR2X1 port map( A => n6, B => n10, Y => SUM(6));
   U4 : XNOR2X1 port map( A => n27, B => n2, Y => SUM(4));
   U5 : NAND2X1 port map( A => n21, B => n23, Y => n2);
   U6 : XOR2X1 port map( A => n48, B => n47, Y => SUM(1));
   U7 : XOR2X1 port map( A => n35, B => n36, Y => SUM(3));
   U8 : AND2X2 port map( A => n33, B => n31, Y => n3);
   U9 : INVX2 port map( A => n39, Y => n38);
   U10 : NAND2X1 port map( A => n45, B => n42, Y => n43);
   U11 : INVX2 port map( A => n49, Y => SUM(0));
   U12 : XNOR2X1 port map( A => n4, B => n5, Y => SUM(7));
   U13 : XOR2X1 port map( A => B(7), B => A(7), Y => n5);
   U14 : AOI21X1 port map( A => n6, B => n7, C => n8, Y => n4);
   U15 : INVX2 port map( A => n9, Y => n8);
   U16 : NAND2X1 port map( A => n7, B => n9, Y => n10);
   U17 : NAND2X1 port map( A => B(6), B => A(6), Y => n9);
   U18 : OR2X2 port map( A => A(6), B => B(6), Y => n7);
   U19 : OAI21X1 port map( A => n11, B => n12, C => n13, Y => n6);
   U20 : INVX2 port map( A => n14, Y => n12);
   U21 : INVX2 port map( A => n15, Y => n11);
   U22 : XNOR2X1 port map( A => n16, B => n1, Y => SUM(5));
   U23 : OAI21X1 port map( A => n17, B => n18, C => n19, Y => n14);
   U24 : AOI21X1 port map( A => n20, B => n21, C => n22, Y => n19);
   U25 : INVX2 port map( A => n23, Y => n22);
   U26 : NAND2X1 port map( A => n24, B => n25, Y => n20);
   U27 : NAND3X1 port map( A => n26, B => n21, C => n3, Y => n18);
   U28 : NAND2X1 port map( A => n13, B => n15, Y => n16);
   U29 : OR2X2 port map( A => A(5), B => B(5), Y => n15);
   U30 : NAND2X1 port map( A => B(5), B => A(5), Y => n13);
   U31 : NAND2X1 port map( A => B(4), B => A(4), Y => n23);
   U32 : OR2X2 port map( A => A(4), B => B(4), Y => n21);
   U33 : OAI21X1 port map( A => n17, B => n28, C => n29, Y => n27);
   U34 : AND2X2 port map( A => n24, B => n25, Y => n29);
   U35 : NAND2X1 port map( A => n30, B => n31, Y => n24);
   U36 : INVX2 port map( A => n32, Y => n30);
   U37 : NAND2X1 port map( A => n3, B => n26, Y => n28);
   U38 : AOI21X1 port map( A => B(0), B => A(0), C => n34, Y => n17);
   U39 : NAND2X1 port map( A => n25, B => n31, Y => n36);
   U40 : OR2X2 port map( A => A(3), B => B(3), Y => n31);
   U41 : NAND2X1 port map( A => B(3), B => A(3), Y => n25);
   U42 : NOR2X1 port map( A => n37, B => n38, Y => n35);
   U43 : NAND3X1 port map( A => n26, B => n33, C => n40, Y => n39);
   U44 : AND2X2 port map( A => B(0), B => A(0), Y => n40);
   U45 : NAND2X1 port map( A => n41, B => n32, Y => n37);
   U46 : NAND2X1 port map( A => n34, B => n33, Y => n41);
   U47 : INVX2 port map( A => n42, Y => n34);
   U48 : XNOR2X1 port map( A => n43, B => n44, Y => SUM(2));
   U49 : NAND2X1 port map( A => n33, B => n32, Y => n44);
   U50 : NAND2X1 port map( A => B(2), B => A(2), Y => n32);
   U51 : OR2X2 port map( A => A(2), B => B(2), Y => n33);
   U52 : NAND2X1 port map( A => n46, B => n26, Y => n45);
   U53 : AND2X2 port map( A => A(0), B => B(0), Y => n46);
   U54 : NAND2X1 port map( A => n42, B => n26, Y => n47);
   U55 : OR2X2 port map( A => A(1), B => B(1), Y => n26);
   U56 : NAND2X1 port map( A => B(1), B => A(1), Y => n42);
   U57 : OAI21X1 port map( A => A(0), B => B(0), C => n48, Y => n49);
   U58 : NAND2X1 port map( A => B(0), B => A(0), Y => n48);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_add_8 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_1_DW01_add_8;

architecture SYN_cla of KSA_1_DW01_add_8 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49 : std_logic;

begin
   
   U2 : BUFX2 port map( A => n6, Y => n1);
   U3 : XNOR2X1 port map( A => n6, B => n10, Y => SUM(6));
   U4 : XNOR2X1 port map( A => n27, B => n2, Y => SUM(4));
   U5 : NAND2X1 port map( A => n21, B => n23, Y => n2);
   U6 : XOR2X1 port map( A => n48, B => n47, Y => SUM(1));
   U7 : XOR2X1 port map( A => n35, B => n36, Y => SUM(3));
   U8 : AND2X2 port map( A => n33, B => n31, Y => n3);
   U9 : INVX2 port map( A => n39, Y => n38);
   U10 : NAND2X1 port map( A => n45, B => n42, Y => n43);
   U11 : INVX2 port map( A => n49, Y => SUM(0));
   U12 : XNOR2X1 port map( A => n4, B => n5, Y => SUM(7));
   U13 : XOR2X1 port map( A => B(7), B => A(7), Y => n5);
   U14 : AOI21X1 port map( A => n1, B => n7, C => n8, Y => n4);
   U15 : INVX2 port map( A => n9, Y => n8);
   U16 : NAND2X1 port map( A => n7, B => n9, Y => n10);
   U17 : NAND2X1 port map( A => B(6), B => A(6), Y => n9);
   U18 : OR2X2 port map( A => A(6), B => B(6), Y => n7);
   U19 : OAI21X1 port map( A => n11, B => n12, C => n13, Y => n6);
   U20 : INVX2 port map( A => n14, Y => n12);
   U21 : INVX2 port map( A => n15, Y => n11);
   U22 : XNOR2X1 port map( A => n14, B => n16, Y => SUM(5));
   U23 : OAI21X1 port map( A => n17, B => n18, C => n19, Y => n14);
   U24 : AOI21X1 port map( A => n20, B => n21, C => n22, Y => n19);
   U25 : INVX2 port map( A => n23, Y => n22);
   U26 : NAND2X1 port map( A => n24, B => n25, Y => n20);
   U27 : NAND3X1 port map( A => n26, B => n21, C => n3, Y => n18);
   U28 : NAND2X1 port map( A => n13, B => n15, Y => n16);
   U29 : OR2X2 port map( A => A(5), B => B(5), Y => n15);
   U30 : NAND2X1 port map( A => B(5), B => A(5), Y => n13);
   U31 : NAND2X1 port map( A => B(4), B => A(4), Y => n23);
   U32 : OR2X2 port map( A => A(4), B => B(4), Y => n21);
   U33 : OAI21X1 port map( A => n17, B => n28, C => n29, Y => n27);
   U34 : AND2X2 port map( A => n24, B => n25, Y => n29);
   U35 : NAND2X1 port map( A => n30, B => n31, Y => n24);
   U36 : INVX2 port map( A => n32, Y => n30);
   U37 : NAND2X1 port map( A => n3, B => n26, Y => n28);
   U38 : AOI21X1 port map( A => B(0), B => A(0), C => n34, Y => n17);
   U39 : NAND2X1 port map( A => n25, B => n31, Y => n36);
   U40 : OR2X2 port map( A => A(3), B => B(3), Y => n31);
   U41 : NAND2X1 port map( A => B(3), B => A(3), Y => n25);
   U42 : NOR2X1 port map( A => n37, B => n38, Y => n35);
   U43 : NAND3X1 port map( A => n26, B => n33, C => n40, Y => n39);
   U44 : AND2X2 port map( A => B(0), B => A(0), Y => n40);
   U45 : NAND2X1 port map( A => n41, B => n32, Y => n37);
   U46 : NAND2X1 port map( A => n34, B => n33, Y => n41);
   U47 : INVX2 port map( A => n42, Y => n34);
   U48 : XNOR2X1 port map( A => n43, B => n44, Y => SUM(2));
   U49 : NAND2X1 port map( A => n33, B => n32, Y => n44);
   U50 : NAND2X1 port map( A => B(2), B => A(2), Y => n32);
   U51 : OR2X2 port map( A => A(2), B => B(2), Y => n33);
   U52 : NAND2X1 port map( A => n46, B => n26, Y => n45);
   U53 : AND2X2 port map( A => A(0), B => B(0), Y => n46);
   U54 : NAND2X1 port map( A => n42, B => n26, Y => n47);
   U55 : OR2X2 port map( A => A(1), B => B(1), Y => n26);
   U56 : NAND2X1 port map( A => B(1), B => A(1), Y => n42);
   U57 : OAI21X1 port map( A => A(0), B => B(0), C => n48, Y => n49);
   U58 : NAND2X1 port map( A => B(0), B => A(0), Y => n48);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity keyreg_1_DW01_add_1 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end keyreg_1_DW01_add_1;

architecture SYN_cla of keyreg_1_DW01_add_1 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41 : std_logic;

begin
   
   U2 : AND2X2 port map( A => n21, B => n17, Y => n1);
   U3 : XNOR2X1 port map( A => n32, B => n33, Y => SUM(3));
   U4 : XOR2X1 port map( A => n27, B => n2, Y => SUM(2));
   U5 : NAND2X1 port map( A => n31, B => n30, Y => n2);
   U6 : NAND2X1 port map( A => n35, B => n36, Y => n22);
   U7 : INVX2 port map( A => n41, Y => SUM(0));
   U8 : XNOR2X1 port map( A => n3, B => n4, Y => SUM(7));
   U9 : XOR2X1 port map( A => B(7), B => A(7), Y => n4);
   U10 : AOI21X1 port map( A => n5, B => n6, C => n7, Y => n3);
   U11 : NAND2X1 port map( A => n8, B => n9, Y => n7);
   U12 : NAND2X1 port map( A => n10, B => n11, Y => n8);
   U13 : AND2X2 port map( A => n12, B => n11, Y => n5);
   U14 : XNOR2X1 port map( A => n13, B => n14, Y => SUM(6));
   U15 : AND2X2 port map( A => n11, B => n9, Y => n14);
   U16 : NAND2X1 port map( A => B(6), B => A(6), Y => n9);
   U17 : OR2X2 port map( A => A(6), B => B(6), Y => n11);
   U18 : AOI21X1 port map( A => n6, B => n12, C => n10, Y => n13);
   U19 : INVX2 port map( A => n15, Y => n10);
   U20 : XNOR2X1 port map( A => n6, B => n16, Y => SUM(5));
   U21 : NAND2X1 port map( A => n12, B => n15, Y => n16);
   U22 : NAND2X1 port map( A => B(5), B => A(5), Y => n15);
   U23 : OR2X2 port map( A => A(5), B => B(5), Y => n12);
   U24 : NAND3X1 port map( A => n17, B => n18, C => n19, Y => n6);
   U25 : NAND3X1 port map( A => n20, B => n21, C => n22, Y => n19);
   U26 : INVX2 port map( A => n23, Y => n20);
   U27 : NAND3X1 port map( A => n24, B => n21, C => n25, Y => n18);
   U28 : XOR2X1 port map( A => n26, B => n1, Y => SUM(4));
   U29 : NAND2X1 port map( A => B(4), B => A(4), Y => n17);
   U30 : OR2X2 port map( A => A(4), B => B(4), Y => n21);
   U31 : OAI21X1 port map( A => n27, B => n23, C => n28, Y => n26);
   U32 : NAND2X1 port map( A => n24, B => n25, Y => n28);
   U33 : NAND2X1 port map( A => n29, B => n30, Y => n25);
   U34 : NAND2X1 port map( A => n31, B => n24, Y => n23);
   U35 : NAND2X1 port map( A => n24, B => n29, Y => n33);
   U36 : NAND2X1 port map( A => B(3), B => A(3), Y => n29);
   U37 : OR2X2 port map( A => A(3), B => B(3), Y => n24);
   U38 : NAND2X1 port map( A => n30, B => n34, Y => n32);
   U39 : NAND2X1 port map( A => n22, B => n31, Y => n34);
   U40 : NAND2X1 port map( A => B(2), B => A(2), Y => n30);
   U41 : OR2X2 port map( A => A(2), B => B(2), Y => n31);
   U42 : INVX2 port map( A => n22, Y => n27);
   U43 : NAND2X1 port map( A => n38, B => n37, Y => n35);
   U44 : AND2X2 port map( A => A(0), B => B(0), Y => n38);
   U45 : XOR2X1 port map( A => n39, B => n40, Y => SUM(1));
   U46 : NAND2X1 port map( A => n37, B => n36, Y => n39);
   U47 : NAND2X1 port map( A => B(1), B => A(1), Y => n36);
   U48 : OR2X2 port map( A => A(1), B => B(1), Y => n37);
   U49 : OAI21X1 port map( A => A(0), B => B(0), C => n40, Y => n41);
   U50 : NAND2X1 port map( A => B(0), B => A(0), Y => n40);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity keyreg_0_DW01_add_1 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end keyreg_0_DW01_add_1;

architecture SYN_cla of keyreg_0_DW01_add_1 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41 : std_logic;

begin
   
   U2 : AND2X2 port map( A => n21, B => n17, Y => n1);
   U3 : XNOR2X1 port map( A => n32, B => n33, Y => SUM(3));
   U4 : XOR2X1 port map( A => n27, B => n2, Y => SUM(2));
   U5 : NAND2X1 port map( A => n31, B => n30, Y => n2);
   U6 : NAND2X1 port map( A => n35, B => n36, Y => n22);
   U7 : INVX2 port map( A => n41, Y => SUM(0));
   U8 : XNOR2X1 port map( A => n3, B => n4, Y => SUM(7));
   U9 : XOR2X1 port map( A => B(7), B => A(7), Y => n4);
   U10 : AOI21X1 port map( A => n5, B => n6, C => n7, Y => n3);
   U11 : NAND2X1 port map( A => n8, B => n9, Y => n7);
   U12 : NAND2X1 port map( A => n10, B => n11, Y => n8);
   U13 : AND2X2 port map( A => n12, B => n11, Y => n5);
   U14 : XNOR2X1 port map( A => n13, B => n14, Y => SUM(6));
   U15 : AND2X2 port map( A => n11, B => n9, Y => n14);
   U16 : NAND2X1 port map( A => B(6), B => A(6), Y => n9);
   U17 : OR2X2 port map( A => A(6), B => B(6), Y => n11);
   U18 : AOI21X1 port map( A => n6, B => n12, C => n10, Y => n13);
   U19 : INVX2 port map( A => n15, Y => n10);
   U20 : XNOR2X1 port map( A => n6, B => n16, Y => SUM(5));
   U21 : NAND2X1 port map( A => n12, B => n15, Y => n16);
   U22 : NAND2X1 port map( A => B(5), B => A(5), Y => n15);
   U23 : OR2X2 port map( A => A(5), B => B(5), Y => n12);
   U24 : NAND3X1 port map( A => n17, B => n18, C => n19, Y => n6);
   U25 : NAND3X1 port map( A => n20, B => n21, C => n22, Y => n19);
   U26 : INVX2 port map( A => n23, Y => n20);
   U27 : NAND3X1 port map( A => n24, B => n21, C => n25, Y => n18);
   U28 : XOR2X1 port map( A => n26, B => n1, Y => SUM(4));
   U29 : NAND2X1 port map( A => B(4), B => A(4), Y => n17);
   U30 : OR2X2 port map( A => A(4), B => B(4), Y => n21);
   U31 : OAI21X1 port map( A => n27, B => n23, C => n28, Y => n26);
   U32 : NAND2X1 port map( A => n24, B => n25, Y => n28);
   U33 : NAND2X1 port map( A => n29, B => n30, Y => n25);
   U34 : NAND2X1 port map( A => n31, B => n24, Y => n23);
   U35 : NAND2X1 port map( A => n24, B => n29, Y => n33);
   U36 : NAND2X1 port map( A => B(3), B => A(3), Y => n29);
   U37 : OR2X2 port map( A => A(3), B => B(3), Y => n24);
   U38 : NAND2X1 port map( A => n30, B => n34, Y => n32);
   U39 : NAND2X1 port map( A => n22, B => n31, Y => n34);
   U40 : NAND2X1 port map( A => B(2), B => A(2), Y => n30);
   U41 : OR2X2 port map( A => A(2), B => B(2), Y => n31);
   U42 : INVX2 port map( A => n22, Y => n27);
   U43 : NAND2X1 port map( A => n38, B => n37, Y => n35);
   U44 : AND2X2 port map( A => A(0), B => B(0), Y => n38);
   U45 : XOR2X1 port map( A => n39, B => n40, Y => SUM(1));
   U46 : NAND2X1 port map( A => n37, B => n36, Y => n39);
   U47 : NAND2X1 port map( A => B(1), B => A(1), Y => n36);
   U48 : OR2X2 port map( A => A(1), B => B(1), Y => n37);
   U49 : OAI21X1 port map( A => A(0), B => B(0), C => n40, Y => n41);
   U50 : NAND2X1 port map( A => B(0), B => A(0), Y => n40);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_add_7 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_1_DW01_add_7;

architecture SYN_cla of KSA_1_DW01_add_7 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40 : std_logic;

begin
   
   U2 : NAND2X1 port map( A => n35, B => n36, Y => n30);
   U3 : INVX2 port map( A => n40, Y => SUM(0));
   U4 : XNOR2X1 port map( A => n1, B => n2, Y => SUM(7));
   U5 : XOR2X1 port map( A => B(7), B => A(7), Y => n2);
   U6 : AOI21X1 port map( A => n3, B => n4, C => n5, Y => n1);
   U7 : INVX2 port map( A => n6, Y => n5);
   U8 : XNOR2X1 port map( A => n3, B => n7, Y => SUM(6));
   U9 : NAND2X1 port map( A => n4, B => n6, Y => n7);
   U10 : NAND2X1 port map( A => B(6), B => A(6), Y => n6);
   U11 : OR2X2 port map( A => A(6), B => B(6), Y => n4);
   U12 : NAND2X1 port map( A => n8, B => n9, Y => n3);
   U13 : NAND2X1 port map( A => n10, B => n11, Y => n9);
   U14 : XNOR2X1 port map( A => n10, B => n12, Y => SUM(5));
   U15 : NAND2X1 port map( A => n8, B => n11, Y => n12);
   U16 : OR2X2 port map( A => A(5), B => B(5), Y => n11);
   U17 : NAND2X1 port map( A => B(5), B => A(5), Y => n8);
   U18 : OAI21X1 port map( A => n13, B => n14, C => n15, Y => n10);
   U19 : AOI21X1 port map( A => n16, B => n17, C => n18, Y => n15);
   U20 : INVX2 port map( A => n19, Y => n18);
   U21 : INVX2 port map( A => n20, Y => n16);
   U22 : NAND2X1 port map( A => n21, B => n17, Y => n14);
   U23 : INVX2 port map( A => n22, Y => n21);
   U24 : XNOR2X1 port map( A => n23, B => n24, Y => SUM(4));
   U25 : OAI21X1 port map( A => n13, B => n22, C => n20, Y => n24);
   U26 : OAI21X1 port map( A => n25, B => n26, C => n27, Y => n20);
   U27 : INVX2 port map( A => n28, Y => n26);
   U28 : NAND2X1 port map( A => n29, B => n27, Y => n22);
   U29 : INVX2 port map( A => n30, Y => n13);
   U30 : NAND2X1 port map( A => n17, B => n19, Y => n23);
   U31 : NAND2X1 port map( A => B(4), B => A(4), Y => n19);
   U32 : OR2X2 port map( A => A(4), B => B(4), Y => n17);
   U33 : XNOR2X1 port map( A => n31, B => n32, Y => SUM(3));
   U34 : AND2X2 port map( A => n27, B => n28, Y => n32);
   U35 : NAND2X1 port map( A => B(3), B => A(3), Y => n28);
   U36 : OR2X2 port map( A => A(3), B => B(3), Y => n27);
   U37 : AOI21X1 port map( A => n30, B => n29, C => n25, Y => n31);
   U38 : INVX2 port map( A => n33, Y => n25);
   U39 : XNOR2X1 port map( A => n34, B => n30, Y => SUM(2));
   U40 : NAND3X1 port map( A => A(0), B => B(0), C => n37, Y => n36);
   U41 : NAND2X1 port map( A => n29, B => n33, Y => n34);
   U42 : NAND2X1 port map( A => B(2), B => A(2), Y => n33);
   U43 : OR2X2 port map( A => A(2), B => B(2), Y => n29);
   U44 : XOR2X1 port map( A => n38, B => n39, Y => SUM(1));
   U45 : NAND2X1 port map( A => n37, B => n35, Y => n38);
   U46 : NAND2X1 port map( A => B(1), B => A(1), Y => n35);
   U47 : OR2X2 port map( A => A(1), B => B(1), Y => n37);
   U48 : OAI21X1 port map( A => A(0), B => B(0), C => n39, Y => n40);
   U49 : NAND2X1 port map( A => B(0), B => A(0), Y => n39);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_add_6 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_1_DW01_add_6;

architecture SYN_cla of KSA_1_DW01_add_6 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38 : std_logic;

begin
   
   U2 : AND2X2 port map( A => n18, B => n14, Y => n1);
   U3 : NAND2X1 port map( A => n33, B => n34, Y => n19);
   U4 : INVX2 port map( A => n38, Y => SUM(0));
   U5 : XNOR2X1 port map( A => n2, B => n3, Y => SUM(7));
   U6 : XOR2X1 port map( A => B(7), B => A(7), Y => n3);
   U7 : AOI21X1 port map( A => n4, B => n5, C => n6, Y => n2);
   U8 : INVX2 port map( A => n7, Y => n6);
   U9 : XNOR2X1 port map( A => n4, B => n8, Y => SUM(6));
   U10 : NAND2X1 port map( A => n5, B => n7, Y => n8);
   U11 : NAND2X1 port map( A => B(6), B => A(6), Y => n7);
   U12 : OR2X2 port map( A => A(6), B => B(6), Y => n5);
   U13 : NAND2X1 port map( A => n9, B => n10, Y => n4);
   U14 : NAND2X1 port map( A => n11, B => n12, Y => n10);
   U15 : XNOR2X1 port map( A => n11, B => n13, Y => SUM(5));
   U16 : NAND2X1 port map( A => n9, B => n12, Y => n13);
   U17 : OR2X2 port map( A => A(5), B => B(5), Y => n12);
   U18 : NAND2X1 port map( A => B(5), B => A(5), Y => n9);
   U19 : NAND3X1 port map( A => n14, B => n15, C => n16, Y => n11);
   U20 : NAND3X1 port map( A => n17, B => n18, C => n19, Y => n16);
   U21 : INVX2 port map( A => n20, Y => n17);
   U22 : NAND3X1 port map( A => n21, B => n18, C => n22, Y => n15);
   U23 : XOR2X1 port map( A => n23, B => n1, Y => SUM(4));
   U24 : NAND2X1 port map( A => B(4), B => A(4), Y => n14);
   U25 : OR2X2 port map( A => A(4), B => B(4), Y => n18);
   U26 : OAI21X1 port map( A => n24, B => n20, C => n25, Y => n23);
   U27 : NAND2X1 port map( A => n21, B => n22, Y => n25);
   U28 : NAND2X1 port map( A => n26, B => n27, Y => n22);
   U29 : NAND2X1 port map( A => n28, B => n21, Y => n20);
   U30 : INVX2 port map( A => n19, Y => n24);
   U31 : XNOR2X1 port map( A => n29, B => n30, Y => SUM(3));
   U32 : AND2X2 port map( A => n21, B => n26, Y => n30);
   U33 : NAND2X1 port map( A => B(3), B => A(3), Y => n26);
   U34 : OR2X2 port map( A => A(3), B => B(3), Y => n21);
   U35 : AOI21X1 port map( A => n19, B => n28, C => n31, Y => n29);
   U36 : INVX2 port map( A => n27, Y => n31);
   U37 : XNOR2X1 port map( A => n32, B => n19, Y => SUM(2));
   U38 : NAND3X1 port map( A => A(0), B => B(0), C => n35, Y => n34);
   U39 : NAND2X1 port map( A => n28, B => n27, Y => n32);
   U40 : NAND2X1 port map( A => B(2), B => A(2), Y => n27);
   U41 : OR2X2 port map( A => A(2), B => B(2), Y => n28);
   U42 : XOR2X1 port map( A => n36, B => n37, Y => SUM(1));
   U43 : NAND2X1 port map( A => n35, B => n33, Y => n36);
   U44 : NAND2X1 port map( A => B(1), B => A(1), Y => n33);
   U45 : OR2X2 port map( A => A(1), B => B(1), Y => n35);
   U46 : OAI21X1 port map( A => A(0), B => B(0), C => n37, Y => n38);
   U47 : NAND2X1 port map( A => B(0), B => A(0), Y => n37);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_add_7 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_0_DW01_add_7;

architecture SYN_cla of KSA_0_DW01_add_7 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40 : std_logic;

begin
   
   U2 : NAND2X1 port map( A => n35, B => n36, Y => n30);
   U3 : INVX2 port map( A => n40, Y => SUM(0));
   U4 : XNOR2X1 port map( A => n1, B => n2, Y => SUM(7));
   U5 : XOR2X1 port map( A => B(7), B => A(7), Y => n2);
   U6 : AOI21X1 port map( A => n3, B => n4, C => n5, Y => n1);
   U7 : INVX2 port map( A => n6, Y => n5);
   U8 : XNOR2X1 port map( A => n3, B => n7, Y => SUM(6));
   U9 : NAND2X1 port map( A => n4, B => n6, Y => n7);
   U10 : NAND2X1 port map( A => B(6), B => A(6), Y => n6);
   U11 : OR2X2 port map( A => A(6), B => B(6), Y => n4);
   U12 : NAND2X1 port map( A => n8, B => n9, Y => n3);
   U13 : NAND2X1 port map( A => n10, B => n11, Y => n9);
   U14 : XNOR2X1 port map( A => n10, B => n12, Y => SUM(5));
   U15 : NAND2X1 port map( A => n8, B => n11, Y => n12);
   U16 : OR2X2 port map( A => A(5), B => B(5), Y => n11);
   U17 : NAND2X1 port map( A => B(5), B => A(5), Y => n8);
   U18 : OAI21X1 port map( A => n13, B => n14, C => n15, Y => n10);
   U19 : AOI21X1 port map( A => n16, B => n17, C => n18, Y => n15);
   U20 : INVX2 port map( A => n19, Y => n18);
   U21 : INVX2 port map( A => n20, Y => n16);
   U22 : NAND2X1 port map( A => n21, B => n17, Y => n14);
   U23 : INVX2 port map( A => n22, Y => n21);
   U24 : XNOR2X1 port map( A => n23, B => n24, Y => SUM(4));
   U25 : OAI21X1 port map( A => n13, B => n22, C => n20, Y => n24);
   U26 : OAI21X1 port map( A => n25, B => n26, C => n27, Y => n20);
   U27 : INVX2 port map( A => n28, Y => n26);
   U28 : NAND2X1 port map( A => n29, B => n27, Y => n22);
   U29 : INVX2 port map( A => n30, Y => n13);
   U30 : NAND2X1 port map( A => n17, B => n19, Y => n23);
   U31 : NAND2X1 port map( A => B(4), B => A(4), Y => n19);
   U32 : OR2X2 port map( A => A(4), B => B(4), Y => n17);
   U33 : XNOR2X1 port map( A => n31, B => n32, Y => SUM(3));
   U34 : AND2X2 port map( A => n27, B => n28, Y => n32);
   U35 : NAND2X1 port map( A => B(3), B => A(3), Y => n28);
   U36 : OR2X2 port map( A => A(3), B => B(3), Y => n27);
   U37 : AOI21X1 port map( A => n30, B => n29, C => n25, Y => n31);
   U38 : INVX2 port map( A => n33, Y => n25);
   U39 : XNOR2X1 port map( A => n34, B => n30, Y => SUM(2));
   U40 : NAND3X1 port map( A => A(0), B => B(0), C => n37, Y => n36);
   U41 : NAND2X1 port map( A => n29, B => n33, Y => n34);
   U42 : NAND2X1 port map( A => B(2), B => A(2), Y => n33);
   U43 : OR2X2 port map( A => A(2), B => B(2), Y => n29);
   U44 : XOR2X1 port map( A => n38, B => n39, Y => SUM(1));
   U45 : NAND2X1 port map( A => n37, B => n35, Y => n38);
   U46 : NAND2X1 port map( A => B(1), B => A(1), Y => n35);
   U47 : OR2X2 port map( A => A(1), B => B(1), Y => n37);
   U48 : OAI21X1 port map( A => A(0), B => B(0), C => n39, Y => n40);
   U49 : NAND2X1 port map( A => B(0), B => A(0), Y => n39);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_add_6 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_0_DW01_add_6;

architecture SYN_cla of KSA_0_DW01_add_6 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38 : std_logic;

begin
   
   U2 : AND2X2 port map( A => n18, B => n14, Y => n1);
   U3 : NAND2X1 port map( A => n33, B => n34, Y => n19);
   U4 : INVX2 port map( A => n38, Y => SUM(0));
   U5 : XNOR2X1 port map( A => n2, B => n3, Y => SUM(7));
   U6 : XOR2X1 port map( A => B(7), B => A(7), Y => n3);
   U7 : AOI21X1 port map( A => n4, B => n5, C => n6, Y => n2);
   U8 : INVX2 port map( A => n7, Y => n6);
   U9 : XNOR2X1 port map( A => n4, B => n8, Y => SUM(6));
   U10 : NAND2X1 port map( A => n5, B => n7, Y => n8);
   U11 : NAND2X1 port map( A => B(6), B => A(6), Y => n7);
   U12 : OR2X2 port map( A => A(6), B => B(6), Y => n5);
   U13 : NAND2X1 port map( A => n9, B => n10, Y => n4);
   U14 : NAND2X1 port map( A => n11, B => n12, Y => n10);
   U15 : XNOR2X1 port map( A => n11, B => n13, Y => SUM(5));
   U16 : NAND2X1 port map( A => n9, B => n12, Y => n13);
   U17 : OR2X2 port map( A => A(5), B => B(5), Y => n12);
   U18 : NAND2X1 port map( A => B(5), B => A(5), Y => n9);
   U19 : NAND3X1 port map( A => n14, B => n15, C => n16, Y => n11);
   U20 : NAND3X1 port map( A => n17, B => n18, C => n19, Y => n16);
   U21 : INVX2 port map( A => n20, Y => n17);
   U22 : NAND3X1 port map( A => n21, B => n18, C => n22, Y => n15);
   U23 : XOR2X1 port map( A => n23, B => n1, Y => SUM(4));
   U24 : NAND2X1 port map( A => B(4), B => A(4), Y => n14);
   U25 : OR2X2 port map( A => A(4), B => B(4), Y => n18);
   U26 : OAI21X1 port map( A => n24, B => n20, C => n25, Y => n23);
   U27 : NAND2X1 port map( A => n21, B => n22, Y => n25);
   U28 : NAND2X1 port map( A => n26, B => n27, Y => n22);
   U29 : NAND2X1 port map( A => n28, B => n21, Y => n20);
   U30 : INVX2 port map( A => n19, Y => n24);
   U31 : XNOR2X1 port map( A => n29, B => n30, Y => SUM(3));
   U32 : AND2X2 port map( A => n21, B => n26, Y => n30);
   U33 : NAND2X1 port map( A => B(3), B => A(3), Y => n26);
   U34 : OR2X2 port map( A => A(3), B => B(3), Y => n21);
   U35 : AOI21X1 port map( A => n19, B => n28, C => n31, Y => n29);
   U36 : INVX2 port map( A => n27, Y => n31);
   U37 : XNOR2X1 port map( A => n32, B => n19, Y => SUM(2));
   U38 : NAND3X1 port map( A => A(0), B => B(0), C => n35, Y => n34);
   U39 : NAND2X1 port map( A => n28, B => n27, Y => n32);
   U40 : NAND2X1 port map( A => B(2), B => A(2), Y => n27);
   U41 : OR2X2 port map( A => A(2), B => B(2), Y => n28);
   U42 : XOR2X1 port map( A => n36, B => n37, Y => SUM(1));
   U43 : NAND2X1 port map( A => n35, B => n33, Y => n36);
   U44 : NAND2X1 port map( A => B(1), B => A(1), Y => n33);
   U45 : OR2X2 port map( A => A(1), B => B(1), Y => n35);
   U46 : OAI21X1 port map( A => A(0), B => B(0), C => n37, Y => n38);
   U47 : NAND2X1 port map( A => B(0), B => A(0), Y => n37);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_inc_1 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_1_DW01_inc_1;

architecture SYN_rpl of KSA_1_DW01_inc_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_1_DW01_inc_0;

architecture SYN_rpl of KSA_1_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX1 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_timer_1_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end uart_timer_1_DW01_inc_0;

architecture SYN_rpl of uart_timer_1_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_tcu_1_DW01_inc_0 is

   port( A : in std_logic_vector (6 downto 0);  SUM : out std_logic_vector (6 
         downto 0));

end tx_tcu_1_DW01_inc_0;

architecture SYN_rpl of tx_tcu_1_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port 
      : std_logic;

begin
   
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_6_port, B => A(6), Y => SUM(6));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_inc_1 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_0_DW01_inc_1;

architecture SYN_rpl of KSA_0_DW01_inc_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_0_DW01_inc_0;

architecture SYN_rpl of KSA_0_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX1 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_timer_0_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end uart_timer_0_DW01_inc_0;

architecture SYN_rpl of uart_timer_0_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_tcu_0_DW01_inc_0 is

   port( A : in std_logic_vector (6 downto 0);  SUM : out std_logic_vector (6 
         downto 0));

end tx_tcu_0_DW01_inc_0;

architecture SYN_rpl of tx_tcu_0_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port 
      : std_logic;

begin
   
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_6_port, B => A(6), Y => SUM(6));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_timer_0 is

   port( CLK, RST, TIMER_TRIG : in std_logic;  STOP_RCVING, SHIFT_STROBE : out 
         std_logic);

end uart_timer_0;

architecture SYN_timerB of uart_timer_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component uart_timer_0_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal state_7_port, state_6_port, state_5_port, state_4_port, state_3_port,
      state_2_port, state_1_port, state_0_port, nextState_7_port, 
      nextState_6_port, nextState_5_port, nextState_4_port, nextState_3_port, 
      nextState_2_port, nextState_1_port, nextState_0_port, N26, N27, N28, N29,
      N30, N31, N32, N33, n10, n17, n19, n20, n21, n22, n23, n24, n25, n26_port
      , n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126 : std_logic;

begin
   
   nextState_reg_0_inst : DFFSR port map( D => n74, CLK => CLK, R => n17, S => 
                           n111, Q => nextState_0_port);
   nextState_reg_1_inst : DFFSR port map( D => n75, CLK => CLK, R => n17, S => 
                           n112, Q => nextState_1_port);
   nextState_reg_2_inst : DFFSR port map( D => n76, CLK => CLK, R => n17, S => 
                           n113, Q => nextState_2_port);
   nextState_reg_3_inst : DFFSR port map( D => n77, CLK => CLK, R => n17, S => 
                           n114, Q => nextState_3_port);
   nextState_reg_4_inst : DFFSR port map( D => n78, CLK => CLK, R => n17, S => 
                           n115, Q => nextState_4_port);
   nextState_reg_5_inst : DFFSR port map( D => n79, CLK => CLK, R => n17, S => 
                           n116, Q => nextState_5_port);
   nextState_reg_6_inst : DFFSR port map( D => n80, CLK => CLK, R => n17, S => 
                           n117, Q => nextState_6_port);
   STOP_RCVING_reg : DFFSR port map( D => n73, CLK => CLK, R => n17, S => n118,
                           Q => STOP_RCVING);
   state_reg_7_inst : DFFSR port map( D => nextState_7_port, CLK => CLK, R => 
                           n17, S => n119, Q => state_7_port);
   state_reg_6_inst : DFFSR port map( D => nextState_6_port, CLK => CLK, R => 
                           n17, S => n120, Q => state_6_port);
   state_reg_5_inst : DFFSR port map( D => nextState_5_port, CLK => CLK, R => 
                           n17, S => n121, Q => state_5_port);
   state_reg_4_inst : DFFSR port map( D => nextState_4_port, CLK => CLK, R => 
                           n17, S => n122, Q => state_4_port);
   state_reg_3_inst : DFFSR port map( D => nextState_3_port, CLK => CLK, R => 
                           n17, S => n123, Q => state_3_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n17, S => n124, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n17, S => n125, Q => state_1_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n17, S => n126, Q => state_0_port);
   n126 <= '1';
   n125 <= '1';
   n124 <= '1';
   n123 <= '1';
   n122 <= '1';
   n121 <= '1';
   n120 <= '1';
   n119 <= '1';
   n118 <= '1';
   n117 <= '1';
   n116 <= '1';
   n115 <= '1';
   n114 <= '1';
   n113 <= '1';
   n112 <= '1';
   n111 <= '1';
   U21 : OR2X2 port map( A => state_7_port, B => n95, Y => n96);
   U38 : OAI21X1 port map( A => n20, B => n27_port, C => n110, Y => n81);
   U39 : NAND2X1 port map( A => N33, B => n109, Y => n110);
   U40 : OAI21X1 port map( A => n26_port, B => n20, C => n108, Y => n80);
   U41 : NAND2X1 port map( A => N32, B => n109, Y => n108);
   U42 : OAI21X1 port map( A => n25, B => n20, C => n107, Y => n79);
   U43 : NAND2X1 port map( A => N31, B => n109, Y => n107);
   U44 : OAI21X1 port map( A => n20, B => n24, C => n106, Y => n78);
   U45 : NAND2X1 port map( A => N30, B => n109, Y => n106);
   U46 : OAI21X1 port map( A => n23, B => n20, C => n105, Y => n77);
   U47 : NAND2X1 port map( A => N29, B => n109, Y => n105);
   U48 : OAI21X1 port map( A => n22, B => n20, C => n104, Y => n76);
   U49 : NAND2X1 port map( A => N28, B => n109, Y => n104);
   U50 : OAI21X1 port map( A => n20, B => n21, C => n103, Y => n75);
   U51 : NAND2X1 port map( A => N27, B => n109, Y => n103);
   U52 : OAI21X1 port map( A => n19, B => n20, C => n102, Y => n74);
   U53 : NAND2X1 port map( A => N26, B => n109, Y => n102);
   U54 : NOR2X1 port map( A => n101, B => n73, Y => n109);
   U55 : NOR2X1 port map( A => n73, B => TIMER_TRIG, Y => n101);
   U56 : NOR2X1 port map( A => n100, B => n99, Y => n73);
   U57 : NAND3X1 port map( A => nextState_6_port, B => nextState_5_port, C => 
                           n98, Y => n99);
   U58 : NOR2X1 port map( A => n22, B => n23, Y => n98);
   U59 : NAND3X1 port map( A => nextState_0_port, B => n21, C => n97, Y => n100
                           );
   U60 : NOR2X1 port map( A => nextState_7_port, B => nextState_4_port, Y => 
                           n97);
   U61 : NOR2X1 port map( A => state_0_port, B => n96, Y => SHIFT_STROBE);
   U62 : AOI21X1 port map( A => n94, B => n32_port, C => n93, Y => n95);
   U63 : OAI21X1 port map( A => n33_port, B => n92, C => n91, Y => n93);
   U64 : NAND3X1 port map( A => state_6_port, B => state_1_port, C => n90, Y =>
                           n91);
   U65 : AOI21X1 port map( A => n89, B => n88, C => state_3_port, Y => n90);
   U66 : NAND3X1 port map( A => n33_port, B => n31_port, C => state_4_port, Y 
                           => n88);
   U67 : NAND3X1 port map( A => state_2_port, B => n32_port, C => state_5_port,
                           Y => n89);
   U68 : NAND2X1 port map( A => state_4_port, B => n87, Y => n92);
   U69 : OAI21X1 port map( A => state_2_port, B => n28_port, C => n86, Y => n94
                           );
   U70 : NAND3X1 port map( A => state_2_port, B => n29_port, C => n30_port, Y 
                           => n86);
   U71 : OAI22X1 port map( A => state_6_port, B => n84, C => n29_port, D => n85
                           , Y => n87);
   U72 : NAND3X1 port map( A => n34, B => n31_port, C => state_3_port, Y => n85
                           );
   U73 : AOI22X1 port map( A => n83, B => state_1_port, C => n82, D => 
                           state_5_port, Y => n84);
   U74 : XOR2X1 port map( A => n34, B => state_3_port, Y => n82);
   U75 : NOR2X1 port map( A => state_5_port, B => state_3_port, Y => n83);
   add_39 : uart_timer_0_DW01_inc_0 port map( A(7) => nextState_7_port, A(6) =>
                           nextState_6_port, A(5) => nextState_5_port, A(4) => 
                           nextState_4_port, A(3) => nextState_3_port, A(2) => 
                           nextState_2_port, A(1) => nextState_1_port, A(0) => 
                           nextState_0_port, SUM(7) => N33, SUM(6) => N32, 
                           SUM(5) => N31, SUM(4) => N30, SUM(3) => N29, SUM(2) 
                           => N28, SUM(1) => N27, SUM(0) => N26);
   nextState_reg_7_inst : DFFSR port map( D => n81, CLK => CLK, R => n17, S => 
                           n10, Q => nextState_7_port);
   n10 <= '1';
   U19 : INVX2 port map( A => RST, Y => n17);
   U22 : INVX2 port map( A => nextState_0_port, Y => n19);
   U23 : INVX2 port map( A => n101, Y => n20);
   U24 : INVX2 port map( A => nextState_1_port, Y => n21);
   U25 : INVX2 port map( A => nextState_2_port, Y => n22);
   U26 : INVX2 port map( A => nextState_3_port, Y => n23);
   U27 : INVX2 port map( A => nextState_4_port, Y => n24);
   U28 : INVX2 port map( A => nextState_5_port, Y => n25);
   U29 : INVX2 port map( A => nextState_6_port, Y => n26_port);
   U30 : INVX2 port map( A => nextState_7_port, Y => n27_port);
   U31 : INVX2 port map( A => n87, Y => n28_port);
   U32 : INVX2 port map( A => state_6_port, Y => n29_port);
   U33 : INVX2 port map( A => n85, Y => n30_port);
   U34 : INVX2 port map( A => state_5_port, Y => n31_port);
   U35 : INVX2 port map( A => state_4_port, Y => n32_port);
   U36 : INVX2 port map( A => state_2_port, Y => n33_port);
   U37 : INVX2 port map( A => state_1_port, Y => n34);

end SYN_timerB;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity keyreg_0 is

   port( CLK, RST, SBE, OE, RBUF_FULL : in std_logic;  RCV_DATA : in 
         std_logic_vector (7 downto 0);  PLAINKEY : out std_logic_vector (63 
         downto 0);  KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR : out 
         std_logic);

end keyreg_0;

architecture SYN_keyb of keyreg_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component keyreg_0_DW01_add_1
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port, 
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port, CLR_RBUFF_port, state_3_port, state_2_port, state_1_port
      , state_0_port, parityError, keyCount_3_port, keyCount_2_port, 
      keyCount_1_port, keyCount_0_port, address_7_port, address_6_port, 
      address_5_port, address_4_port, address_3_port, address_2_port, 
      address_1_port, address_0_port, currentPlainKey_63_port, 
      currentPlainKey_62_port, currentPlainKey_61_port, currentPlainKey_60_port
      , currentPlainKey_59_port, currentPlainKey_58_port, 
      currentPlainKey_57_port, currentPlainKey_56_port, currentPlainKey_55_port
      , currentPlainKey_54_port, currentPlainKey_53_port, 
      currentPlainKey_52_port, currentPlainKey_51_port, currentPlainKey_50_port
      , currentPlainKey_49_port, currentPlainKey_48_port, 
      currentPlainKey_47_port, currentPlainKey_46_port, currentPlainKey_45_port
      , currentPlainKey_44_port, currentPlainKey_43_port, 
      currentPlainKey_42_port, currentPlainKey_41_port, currentPlainKey_40_port
      , currentPlainKey_39_port, currentPlainKey_38_port, 
      currentPlainKey_37_port, currentPlainKey_36_port, currentPlainKey_35_port
      , currentPlainKey_34_port, currentPlainKey_33_port, 
      currentPlainKey_32_port, currentPlainKey_31_port, currentPlainKey_30_port
      , currentPlainKey_29_port, currentPlainKey_28_port, 
      currentPlainKey_27_port, currentPlainKey_26_port, currentPlainKey_25_port
      , currentPlainKey_24_port, currentPlainKey_23_port, 
      currentPlainKey_22_port, currentPlainKey_21_port, currentPlainKey_20_port
      , currentPlainKey_19_port, currentPlainKey_18_port, 
      currentPlainKey_17_port, currentPlainKey_16_port, currentPlainKey_15_port
      , currentPlainKey_14_port, currentPlainKey_13_port, 
      currentPlainKey_12_port, currentPlainKey_11_port, currentPlainKey_10_port
      , currentPlainKey_9_port, currentPlainKey_8_port, currentPlainKey_7_port,
      currentPlainKey_6_port, currentPlainKey_5_port, currentPlainKey_4_port, 
      currentPlainKey_3_port, currentPlainKey_2_port, currentPlainKey_1_port, 
      currentPlainKey_0_port, parityAccumulator_7_port, 
      parityAccumulator_6_port, parityAccumulator_5_port, 
      parityAccumulator_4_port, parityAccumulator_3_port, 
      parityAccumulator_2_port, parityAccumulator_1_port, 
      parityAccumulator_0_port, nextParityError, N1792, N1793, N1794, N1795, 
      N1796, N1797, N1798, N1799, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n14
      , n16, n17, n19, n20, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, 
      n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63, n65, n67, n69
      , n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95, n97, 
      n99, n101, n103, n105, n107, n109, n111, n113, n115, n117, n119, n121, 
      n123, n125, n127, n129, n131, n133, n135, n137, n139, n141, n143, n145, 
      n147, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1267, n1268, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
      n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
      n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
      n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
      n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, 
      n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
      n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
      n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
      n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
      n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
      n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
      n1790, n1791, n1792_port, n1793_port, n1794_port, n1795_port, n1796_port,
      n1797_port, n1798_port, n1799_port, n1800, n1801, n1802, n1803, n1804, 
      n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, 
      n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
      n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, 
      n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, 
      n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
      n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, 
      n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
      n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, 
      n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
      n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, 
      n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
      n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
      n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, 
      n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, 
      n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
      n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
      n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
      n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, 
      n1985, n1986, n1987, n1988, n1989, n_1020 : std_logic;

begin
   PLAINKEY <= ( PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port, 
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port );
   CLR_RBUFF <= CLR_RBUFF_port;
   
   n1989 <= '0';
   keyCount_reg_0_inst : DFFPOSX1 port map( D => n1762, CLK => CLK, Q => 
                           keyCount_0_port);
   keyCount_reg_2_inst : DFFPOSX1 port map( D => n1769, CLK => CLK, Q => 
                           keyCount_2_port);
   keyCount_reg_3_inst : DFFPOSX1 port map( D => n1763, CLK => CLK, Q => 
                           keyCount_3_port);
   state_reg_0_inst : DFFSR port map( D => n1765, CLK => CLK, R => n293, S => 
                           n1850, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => n1767, CLK => CLK, R => n290, S => 
                           n1851, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => n1766, CLK => CLK, R => n292, S => 
                           n1852, Q => state_2_port);
   state_reg_3_inst : DFFSR port map( D => n1764, CLK => CLK, R => n291, S => 
                           n1853, Q => state_3_port);
   parityAccumulator_reg_0_inst : DFFPOSX1 port map( D => n1770, CLK => CLK, Q 
                           => parityAccumulator_0_port);
   parityAccumulator_reg_1_inst : DFFPOSX1 port map( D => n1771, CLK => CLK, Q 
                           => parityAccumulator_1_port);
   parityAccumulator_reg_2_inst : DFFPOSX1 port map( D => n1772, CLK => CLK, Q 
                           => parityAccumulator_2_port);
   parityAccumulator_reg_3_inst : DFFPOSX1 port map( D => n1773, CLK => CLK, Q 
                           => parityAccumulator_3_port);
   parityAccumulator_reg_4_inst : DFFPOSX1 port map( D => n1774, CLK => CLK, Q 
                           => parityAccumulator_4_port);
   parityAccumulator_reg_5_inst : DFFPOSX1 port map( D => n1775, CLK => CLK, Q 
                           => parityAccumulator_5_port);
   parityAccumulator_reg_6_inst : DFFPOSX1 port map( D => n1776, CLK => CLK, Q 
                           => parityAccumulator_6_port);
   parityAccumulator_reg_7_inst : DFFPOSX1 port map( D => n1777, CLK => CLK, Q 
                           => parityAccumulator_7_port);
   keyCount_reg_1_inst : DFFPOSX1 port map( D => n1768, CLK => CLK, Q => 
                           keyCount_1_port);
   PARITY_ERROR_reg : DFFSR port map( D => nextParityError, CLK => CLK, R => 
                           n292, S => n1854, Q => PARITY_ERROR);
   parityError_reg : DFFSR port map( D => nextParityError, CLK => CLK, R => 
                           n292, S => n1855, Q => parityError);
   address_reg_7_inst : DFFPOSX1 port map( D => n1778, CLK => CLK, Q => 
                           address_7_port);
   address_reg_6_inst : DFFPOSX1 port map( D => n1779, CLK => CLK, Q => 
                           address_6_port);
   address_reg_5_inst : DFFPOSX1 port map( D => n1780, CLK => CLK, Q => 
                           address_5_port);
   address_reg_4_inst : DFFPOSX1 port map( D => n1781, CLK => CLK, Q => 
                           address_4_port);
   address_reg_3_inst : DFFPOSX1 port map( D => n1782, CLK => CLK, Q => 
                           address_3_port);
   address_reg_2_inst : DFFPOSX1 port map( D => n1783, CLK => CLK, Q => 
                           address_2_port);
   address_reg_1_inst : DFFPOSX1 port map( D => n1784, CLK => CLK, Q => 
                           address_1_port);
   address_reg_0_inst : DFFPOSX1 port map( D => n1785, CLK => CLK, Q => 
                           address_0_port);
   currentPlainKey_reg_63_inst : DFFPOSX1 port map( D => n1849, CLK => CLK, Q 
                           => currentPlainKey_63_port);
   currentPlainKey_reg_62_inst : DFFPOSX1 port map( D => n1848, CLK => CLK, Q 
                           => currentPlainKey_62_port);
   currentPlainKey_reg_61_inst : DFFPOSX1 port map( D => n1847, CLK => CLK, Q 
                           => currentPlainKey_61_port);
   currentPlainKey_reg_60_inst : DFFPOSX1 port map( D => n1846, CLK => CLK, Q 
                           => currentPlainKey_60_port);
   currentPlainKey_reg_59_inst : DFFPOSX1 port map( D => n1845, CLK => CLK, Q 
                           => currentPlainKey_59_port);
   currentPlainKey_reg_58_inst : DFFPOSX1 port map( D => n1844, CLK => CLK, Q 
                           => currentPlainKey_58_port);
   currentPlainKey_reg_57_inst : DFFPOSX1 port map( D => n1843, CLK => CLK, Q 
                           => currentPlainKey_57_port);
   currentPlainKey_reg_56_inst : DFFPOSX1 port map( D => n1842, CLK => CLK, Q 
                           => currentPlainKey_56_port);
   currentPlainKey_reg_55_inst : DFFPOSX1 port map( D => n1841, CLK => CLK, Q 
                           => currentPlainKey_55_port);
   currentPlainKey_reg_54_inst : DFFPOSX1 port map( D => n1840, CLK => CLK, Q 
                           => currentPlainKey_54_port);
   currentPlainKey_reg_53_inst : DFFPOSX1 port map( D => n1839, CLK => CLK, Q 
                           => currentPlainKey_53_port);
   currentPlainKey_reg_52_inst : DFFPOSX1 port map( D => n1838, CLK => CLK, Q 
                           => currentPlainKey_52_port);
   currentPlainKey_reg_51_inst : DFFPOSX1 port map( D => n1837, CLK => CLK, Q 
                           => currentPlainKey_51_port);
   currentPlainKey_reg_50_inst : DFFPOSX1 port map( D => n1836, CLK => CLK, Q 
                           => currentPlainKey_50_port);
   currentPlainKey_reg_49_inst : DFFPOSX1 port map( D => n1835, CLK => CLK, Q 
                           => currentPlainKey_49_port);
   currentPlainKey_reg_48_inst : DFFPOSX1 port map( D => n1834, CLK => CLK, Q 
                           => currentPlainKey_48_port);
   currentPlainKey_reg_47_inst : DFFPOSX1 port map( D => n1833, CLK => CLK, Q 
                           => currentPlainKey_47_port);
   currentPlainKey_reg_46_inst : DFFPOSX1 port map( D => n1832, CLK => CLK, Q 
                           => currentPlainKey_46_port);
   currentPlainKey_reg_45_inst : DFFPOSX1 port map( D => n1831, CLK => CLK, Q 
                           => currentPlainKey_45_port);
   currentPlainKey_reg_44_inst : DFFPOSX1 port map( D => n1830, CLK => CLK, Q 
                           => currentPlainKey_44_port);
   currentPlainKey_reg_43_inst : DFFPOSX1 port map( D => n1829, CLK => CLK, Q 
                           => currentPlainKey_43_port);
   currentPlainKey_reg_42_inst : DFFPOSX1 port map( D => n1828, CLK => CLK, Q 
                           => currentPlainKey_42_port);
   currentPlainKey_reg_41_inst : DFFPOSX1 port map( D => n1827, CLK => CLK, Q 
                           => currentPlainKey_41_port);
   currentPlainKey_reg_40_inst : DFFPOSX1 port map( D => n1826, CLK => CLK, Q 
                           => currentPlainKey_40_port);
   currentPlainKey_reg_39_inst : DFFPOSX1 port map( D => n1825, CLK => CLK, Q 
                           => currentPlainKey_39_port);
   currentPlainKey_reg_38_inst : DFFPOSX1 port map( D => n1824, CLK => CLK, Q 
                           => currentPlainKey_38_port);
   currentPlainKey_reg_37_inst : DFFPOSX1 port map( D => n1823, CLK => CLK, Q 
                           => currentPlainKey_37_port);
   currentPlainKey_reg_36_inst : DFFPOSX1 port map( D => n1822, CLK => CLK, Q 
                           => currentPlainKey_36_port);
   currentPlainKey_reg_35_inst : DFFPOSX1 port map( D => n1821, CLK => CLK, Q 
                           => currentPlainKey_35_port);
   currentPlainKey_reg_34_inst : DFFPOSX1 port map( D => n1820, CLK => CLK, Q 
                           => currentPlainKey_34_port);
   currentPlainKey_reg_33_inst : DFFPOSX1 port map( D => n1819, CLK => CLK, Q 
                           => currentPlainKey_33_port);
   currentPlainKey_reg_32_inst : DFFPOSX1 port map( D => n1818, CLK => CLK, Q 
                           => currentPlainKey_32_port);
   currentPlainKey_reg_31_inst : DFFPOSX1 port map( D => n1817, CLK => CLK, Q 
                           => currentPlainKey_31_port);
   currentPlainKey_reg_30_inst : DFFPOSX1 port map( D => n1816, CLK => CLK, Q 
                           => currentPlainKey_30_port);
   currentPlainKey_reg_29_inst : DFFPOSX1 port map( D => n1815, CLK => CLK, Q 
                           => currentPlainKey_29_port);
   currentPlainKey_reg_28_inst : DFFPOSX1 port map( D => n1814, CLK => CLK, Q 
                           => currentPlainKey_28_port);
   currentPlainKey_reg_27_inst : DFFPOSX1 port map( D => n1813, CLK => CLK, Q 
                           => currentPlainKey_27_port);
   currentPlainKey_reg_26_inst : DFFPOSX1 port map( D => n1812, CLK => CLK, Q 
                           => currentPlainKey_26_port);
   currentPlainKey_reg_25_inst : DFFPOSX1 port map( D => n1811, CLK => CLK, Q 
                           => currentPlainKey_25_port);
   currentPlainKey_reg_24_inst : DFFPOSX1 port map( D => n1810, CLK => CLK, Q 
                           => currentPlainKey_24_port);
   currentPlainKey_reg_23_inst : DFFPOSX1 port map( D => n1809, CLK => CLK, Q 
                           => currentPlainKey_23_port);
   currentPlainKey_reg_22_inst : DFFPOSX1 port map( D => n1808, CLK => CLK, Q 
                           => currentPlainKey_22_port);
   currentPlainKey_reg_21_inst : DFFPOSX1 port map( D => n1807, CLK => CLK, Q 
                           => currentPlainKey_21_port);
   currentPlainKey_reg_20_inst : DFFPOSX1 port map( D => n1806, CLK => CLK, Q 
                           => currentPlainKey_20_port);
   currentPlainKey_reg_19_inst : DFFPOSX1 port map( D => n1805, CLK => CLK, Q 
                           => currentPlainKey_19_port);
   currentPlainKey_reg_18_inst : DFFPOSX1 port map( D => n1804, CLK => CLK, Q 
                           => currentPlainKey_18_port);
   currentPlainKey_reg_17_inst : DFFPOSX1 port map( D => n1803, CLK => CLK, Q 
                           => currentPlainKey_17_port);
   currentPlainKey_reg_16_inst : DFFPOSX1 port map( D => n1802, CLK => CLK, Q 
                           => currentPlainKey_16_port);
   currentPlainKey_reg_15_inst : DFFPOSX1 port map( D => n1801, CLK => CLK, Q 
                           => currentPlainKey_15_port);
   currentPlainKey_reg_14_inst : DFFPOSX1 port map( D => n1800, CLK => CLK, Q 
                           => currentPlainKey_14_port);
   currentPlainKey_reg_13_inst : DFFPOSX1 port map( D => n1799_port, CLK => CLK
                           , Q => currentPlainKey_13_port);
   currentPlainKey_reg_12_inst : DFFPOSX1 port map( D => n1798_port, CLK => CLK
                           , Q => currentPlainKey_12_port);
   currentPlainKey_reg_11_inst : DFFPOSX1 port map( D => n1797_port, CLK => CLK
                           , Q => currentPlainKey_11_port);
   currentPlainKey_reg_10_inst : DFFPOSX1 port map( D => n1796_port, CLK => CLK
                           , Q => currentPlainKey_10_port);
   currentPlainKey_reg_9_inst : DFFPOSX1 port map( D => n1795_port, CLK => CLK,
                           Q => currentPlainKey_9_port);
   currentPlainKey_reg_8_inst : DFFPOSX1 port map( D => n1794_port, CLK => CLK,
                           Q => currentPlainKey_8_port);
   currentPlainKey_reg_7_inst : DFFPOSX1 port map( D => n1793_port, CLK => CLK,
                           Q => currentPlainKey_7_port);
   currentPlainKey_reg_6_inst : DFFPOSX1 port map( D => n1792_port, CLK => CLK,
                           Q => currentPlainKey_6_port);
   currentPlainKey_reg_5_inst : DFFPOSX1 port map( D => n1791, CLK => CLK, Q =>
                           currentPlainKey_5_port);
   currentPlainKey_reg_4_inst : DFFPOSX1 port map( D => n1790, CLK => CLK, Q =>
                           currentPlainKey_4_port);
   currentPlainKey_reg_3_inst : DFFPOSX1 port map( D => n1789, CLK => CLK, Q =>
                           currentPlainKey_3_port);
   currentPlainKey_reg_2_inst : DFFPOSX1 port map( D => n1788, CLK => CLK, Q =>
                           currentPlainKey_2_port);
   currentPlainKey_reg_1_inst : DFFPOSX1 port map( D => n1787, CLK => CLK, Q =>
                           currentPlainKey_1_port);
   currentPlainKey_reg_0_inst : DFFPOSX1 port map( D => n1786, CLK => CLK, Q =>
                           currentPlainKey_0_port);
   PLAINKEY_reg_63_inst : DFFPOSX1 port map( D => n1856, CLK => CLK, Q => 
                           PLAINKEY_63_port);
   PLAINKEY_reg_62_inst : DFFPOSX1 port map( D => n1857, CLK => CLK, Q => 
                           PLAINKEY_62_port);
   PLAINKEY_reg_61_inst : DFFPOSX1 port map( D => n1858, CLK => CLK, Q => 
                           PLAINKEY_61_port);
   PLAINKEY_reg_60_inst : DFFPOSX1 port map( D => n1859, CLK => CLK, Q => 
                           PLAINKEY_60_port);
   PLAINKEY_reg_59_inst : DFFPOSX1 port map( D => n1860, CLK => CLK, Q => 
                           PLAINKEY_59_port);
   PLAINKEY_reg_58_inst : DFFPOSX1 port map( D => n1861, CLK => CLK, Q => 
                           PLAINKEY_58_port);
   PLAINKEY_reg_57_inst : DFFPOSX1 port map( D => n1862, CLK => CLK, Q => 
                           PLAINKEY_57_port);
   PLAINKEY_reg_56_inst : DFFPOSX1 port map( D => n1863, CLK => CLK, Q => 
                           PLAINKEY_56_port);
   PLAINKEY_reg_55_inst : DFFPOSX1 port map( D => n1864, CLK => CLK, Q => 
                           PLAINKEY_55_port);
   PLAINKEY_reg_54_inst : DFFPOSX1 port map( D => n1865, CLK => CLK, Q => 
                           PLAINKEY_54_port);
   PLAINKEY_reg_53_inst : DFFPOSX1 port map( D => n1866, CLK => CLK, Q => 
                           PLAINKEY_53_port);
   PLAINKEY_reg_52_inst : DFFPOSX1 port map( D => n1867, CLK => CLK, Q => 
                           PLAINKEY_52_port);
   PLAINKEY_reg_51_inst : DFFPOSX1 port map( D => n1868, CLK => CLK, Q => 
                           PLAINKEY_51_port);
   PLAINKEY_reg_50_inst : DFFPOSX1 port map( D => n1869, CLK => CLK, Q => 
                           PLAINKEY_50_port);
   PLAINKEY_reg_49_inst : DFFPOSX1 port map( D => n1870, CLK => CLK, Q => 
                           PLAINKEY_49_port);
   PLAINKEY_reg_48_inst : DFFPOSX1 port map( D => n1871, CLK => CLK, Q => 
                           PLAINKEY_48_port);
   PLAINKEY_reg_47_inst : DFFPOSX1 port map( D => n1872, CLK => CLK, Q => 
                           PLAINKEY_47_port);
   PLAINKEY_reg_46_inst : DFFPOSX1 port map( D => n1873, CLK => CLK, Q => 
                           PLAINKEY_46_port);
   PLAINKEY_reg_45_inst : DFFPOSX1 port map( D => n1874, CLK => CLK, Q => 
                           PLAINKEY_45_port);
   PLAINKEY_reg_44_inst : DFFPOSX1 port map( D => n1875, CLK => CLK, Q => 
                           PLAINKEY_44_port);
   PLAINKEY_reg_43_inst : DFFPOSX1 port map( D => n1876, CLK => CLK, Q => 
                           PLAINKEY_43_port);
   PLAINKEY_reg_42_inst : DFFPOSX1 port map( D => n1877, CLK => CLK, Q => 
                           PLAINKEY_42_port);
   PLAINKEY_reg_41_inst : DFFPOSX1 port map( D => n1878, CLK => CLK, Q => 
                           PLAINKEY_41_port);
   PLAINKEY_reg_40_inst : DFFPOSX1 port map( D => n1879, CLK => CLK, Q => 
                           PLAINKEY_40_port);
   PLAINKEY_reg_39_inst : DFFPOSX1 port map( D => n1880, CLK => CLK, Q => 
                           PLAINKEY_39_port);
   PLAINKEY_reg_38_inst : DFFPOSX1 port map( D => n1881, CLK => CLK, Q => 
                           PLAINKEY_38_port);
   PLAINKEY_reg_37_inst : DFFPOSX1 port map( D => n1882, CLK => CLK, Q => 
                           PLAINKEY_37_port);
   PLAINKEY_reg_36_inst : DFFPOSX1 port map( D => n1883, CLK => CLK, Q => 
                           PLAINKEY_36_port);
   PLAINKEY_reg_35_inst : DFFPOSX1 port map( D => n1884, CLK => CLK, Q => 
                           PLAINKEY_35_port);
   PLAINKEY_reg_34_inst : DFFPOSX1 port map( D => n1885, CLK => CLK, Q => 
                           PLAINKEY_34_port);
   PLAINKEY_reg_33_inst : DFFPOSX1 port map( D => n1886, CLK => CLK, Q => 
                           PLAINKEY_33_port);
   PLAINKEY_reg_32_inst : DFFPOSX1 port map( D => n1887, CLK => CLK, Q => 
                           PLAINKEY_32_port);
   PLAINKEY_reg_31_inst : DFFPOSX1 port map( D => n1888, CLK => CLK, Q => 
                           PLAINKEY_31_port);
   PLAINKEY_reg_30_inst : DFFPOSX1 port map( D => n1889, CLK => CLK, Q => 
                           PLAINKEY_30_port);
   PLAINKEY_reg_29_inst : DFFPOSX1 port map( D => n1890, CLK => CLK, Q => 
                           PLAINKEY_29_port);
   PLAINKEY_reg_28_inst : DFFPOSX1 port map( D => n1891, CLK => CLK, Q => 
                           PLAINKEY_28_port);
   PLAINKEY_reg_27_inst : DFFPOSX1 port map( D => n1892, CLK => CLK, Q => 
                           PLAINKEY_27_port);
   PLAINKEY_reg_26_inst : DFFPOSX1 port map( D => n1893, CLK => CLK, Q => 
                           PLAINKEY_26_port);
   PLAINKEY_reg_25_inst : DFFPOSX1 port map( D => n1894, CLK => CLK, Q => 
                           PLAINKEY_25_port);
   PLAINKEY_reg_24_inst : DFFPOSX1 port map( D => n1895, CLK => CLK, Q => 
                           PLAINKEY_24_port);
   PLAINKEY_reg_23_inst : DFFPOSX1 port map( D => n1896, CLK => CLK, Q => 
                           PLAINKEY_23_port);
   PLAINKEY_reg_22_inst : DFFPOSX1 port map( D => n1897, CLK => CLK, Q => 
                           PLAINKEY_22_port);
   PLAINKEY_reg_21_inst : DFFPOSX1 port map( D => n1898, CLK => CLK, Q => 
                           PLAINKEY_21_port);
   PLAINKEY_reg_20_inst : DFFPOSX1 port map( D => n1899, CLK => CLK, Q => 
                           PLAINKEY_20_port);
   PLAINKEY_reg_19_inst : DFFPOSX1 port map( D => n1900, CLK => CLK, Q => 
                           PLAINKEY_19_port);
   PLAINKEY_reg_18_inst : DFFPOSX1 port map( D => n1901, CLK => CLK, Q => 
                           PLAINKEY_18_port);
   PLAINKEY_reg_17_inst : DFFPOSX1 port map( D => n1902, CLK => CLK, Q => 
                           PLAINKEY_17_port);
   PLAINKEY_reg_16_inst : DFFPOSX1 port map( D => n1903, CLK => CLK, Q => 
                           PLAINKEY_16_port);
   PLAINKEY_reg_15_inst : DFFPOSX1 port map( D => n1904, CLK => CLK, Q => 
                           PLAINKEY_15_port);
   PLAINKEY_reg_14_inst : DFFPOSX1 port map( D => n1905, CLK => CLK, Q => 
                           PLAINKEY_14_port);
   PLAINKEY_reg_13_inst : DFFPOSX1 port map( D => n1906, CLK => CLK, Q => 
                           PLAINKEY_13_port);
   PLAINKEY_reg_12_inst : DFFPOSX1 port map( D => n1907, CLK => CLK, Q => 
                           PLAINKEY_12_port);
   PLAINKEY_reg_11_inst : DFFPOSX1 port map( D => n1908, CLK => CLK, Q => 
                           PLAINKEY_11_port);
   PLAINKEY_reg_10_inst : DFFPOSX1 port map( D => n1909, CLK => CLK, Q => 
                           PLAINKEY_10_port);
   PLAINKEY_reg_9_inst : DFFPOSX1 port map( D => n1910, CLK => CLK, Q => 
                           PLAINKEY_9_port);
   PLAINKEY_reg_8_inst : DFFPOSX1 port map( D => n1911, CLK => CLK, Q => 
                           PLAINKEY_8_port);
   PLAINKEY_reg_7_inst : DFFPOSX1 port map( D => n1912, CLK => CLK, Q => 
                           PLAINKEY_7_port);
   PLAINKEY_reg_6_inst : DFFPOSX1 port map( D => n1913, CLK => CLK, Q => 
                           PLAINKEY_6_port);
   PLAINKEY_reg_5_inst : DFFPOSX1 port map( D => n1914, CLK => CLK, Q => 
                           PLAINKEY_5_port);
   PLAINKEY_reg_4_inst : DFFPOSX1 port map( D => n1915, CLK => CLK, Q => 
                           PLAINKEY_4_port);
   PLAINKEY_reg_3_inst : DFFPOSX1 port map( D => n1916, CLK => CLK, Q => 
                           PLAINKEY_3_port);
   PLAINKEY_reg_2_inst : DFFPOSX1 port map( D => n1917, CLK => CLK, Q => 
                           PLAINKEY_2_port);
   PLAINKEY_reg_1_inst : DFFPOSX1 port map( D => n1918, CLK => CLK, Q => 
                           PLAINKEY_1_port);
   PLAINKEY_reg_0_inst : DFFPOSX1 port map( D => n1919, CLK => CLK, Q => 
                           PLAINKEY_0_port);
   U9 : NAND3X1 port map( A => parityAccumulator_7_port, B => 
                           parityAccumulator_6_port, C => n1986, Y => n1987);
   U10 : NOR2X1 port map( A => n1692, B => n1693, Y => n1986);
   U11 : NAND3X1 port map( A => parityAccumulator_3_port, B => 
                           parityAccumulator_2_port, C => n1985, Y => n1988);
   U12 : NOR2X1 port map( A => n1688, B => n1689, Y => n1985);
   U13 : OAI21X1 port map( A => RST, B => n1759, C => n1984, Y => n1919);
   U14 : NAND2X1 port map( A => PLAINKEY_0_port, B => n286, Y => n1984);
   U15 : OAI21X1 port map( A => n284, B => n1758, C => n1983, Y => n1918);
   U16 : NAND2X1 port map( A => PLAINKEY_1_port, B => n288, Y => n1983);
   U17 : OAI21X1 port map( A => n285, B => n1757, C => n1982, Y => n1917);
   U18 : NAND2X1 port map( A => PLAINKEY_2_port, B => n288, Y => n1982);
   U19 : OAI21X1 port map( A => n287, B => n1756, C => n1981, Y => n1916);
   U20 : NAND2X1 port map( A => PLAINKEY_3_port, B => n288, Y => n1981);
   U21 : OAI21X1 port map( A => RST, B => n1755, C => n1980, Y => n1915);
   U22 : NAND2X1 port map( A => PLAINKEY_4_port, B => n288, Y => n1980);
   U24 : OAI21X1 port map( A => n286, B => n1754, C => n1979, Y => n1914);
   U25 : NAND2X1 port map( A => PLAINKEY_5_port, B => n288, Y => n1979);
   U27 : OAI21X1 port map( A => n284, B => n1753, C => n1978, Y => n1913);
   U28 : NAND2X1 port map( A => PLAINKEY_6_port, B => n288, Y => n1978);
   U30 : OAI21X1 port map( A => RST, B => n1752, C => n1977, Y => n1912);
   U31 : NAND2X1 port map( A => PLAINKEY_7_port, B => n288, Y => n1977);
   U33 : OAI21X1 port map( A => n288, B => n1751, C => n1976, Y => n1911);
   U34 : NAND2X1 port map( A => PLAINKEY_8_port, B => n288, Y => n1976);
   U36 : OAI21X1 port map( A => n284, B => n1750, C => n1975, Y => n1910);
   U37 : NAND2X1 port map( A => PLAINKEY_9_port, B => n288, Y => n1975);
   U39 : OAI21X1 port map( A => n284, B => n1749, C => n1974, Y => n1909);
   U40 : NAND2X1 port map( A => PLAINKEY_10_port, B => n288, Y => n1974);
   U42 : OAI21X1 port map( A => n284, B => n1748, C => n1973, Y => n1908);
   U43 : NAND2X1 port map( A => PLAINKEY_11_port, B => n288, Y => n1973);
   U45 : OAI21X1 port map( A => n284, B => n1747, C => n1972, Y => n1907);
   U46 : NAND2X1 port map( A => PLAINKEY_12_port, B => n288, Y => n1972);
   U48 : OAI21X1 port map( A => n284, B => n1746, C => n1971, Y => n1906);
   U49 : NAND2X1 port map( A => PLAINKEY_13_port, B => n288, Y => n1971);
   U51 : OAI21X1 port map( A => n284, B => n1745, C => n1970, Y => n1905);
   U52 : NAND2X1 port map( A => PLAINKEY_14_port, B => n288, Y => n1970);
   U54 : OAI21X1 port map( A => n284, B => n1744, C => n1969, Y => n1904);
   U55 : NAND2X1 port map( A => PLAINKEY_15_port, B => n288, Y => n1969);
   U57 : OAI21X1 port map( A => n285, B => n1743, C => n1968, Y => n1903);
   U58 : NAND2X1 port map( A => PLAINKEY_16_port, B => n288, Y => n1968);
   U60 : OAI21X1 port map( A => n285, B => n1742, C => n1967, Y => n1902);
   U61 : NAND2X1 port map( A => PLAINKEY_17_port, B => n288, Y => n1967);
   U63 : OAI21X1 port map( A => n285, B => n1741, C => n1966, Y => n1901);
   U64 : NAND2X1 port map( A => PLAINKEY_18_port, B => n288, Y => n1966);
   U66 : OAI21X1 port map( A => n285, B => n1740, C => n1965, Y => n1900);
   U67 : NAND2X1 port map( A => PLAINKEY_19_port, B => n288, Y => n1965);
   U69 : OAI21X1 port map( A => n285, B => n1739, C => n1964, Y => n1899);
   U70 : NAND2X1 port map( A => PLAINKEY_20_port, B => n288, Y => n1964);
   U72 : OAI21X1 port map( A => n285, B => n1738, C => n1963, Y => n1898);
   U73 : NAND2X1 port map( A => PLAINKEY_21_port, B => n288, Y => n1963);
   U75 : OAI21X1 port map( A => n285, B => n1737, C => n1962, Y => n1897);
   U76 : NAND2X1 port map( A => PLAINKEY_22_port, B => n288, Y => n1962);
   U78 : OAI21X1 port map( A => n286, B => n1736, C => n1961, Y => n1896);
   U79 : NAND2X1 port map( A => PLAINKEY_23_port, B => n287, Y => n1961);
   U81 : OAI21X1 port map( A => n285, B => n1735, C => n1960, Y => n1895);
   U82 : NAND2X1 port map( A => PLAINKEY_24_port, B => n285, Y => n1960);
   U84 : OAI21X1 port map( A => n284, B => n1734, C => n1959, Y => n1894);
   U85 : NAND2X1 port map( A => PLAINKEY_25_port, B => n287, Y => n1959);
   U87 : OAI21X1 port map( A => n286, B => n1733, C => n1958, Y => n1893);
   U88 : NAND2X1 port map( A => PLAINKEY_26_port, B => n286, Y => n1958);
   U90 : OAI21X1 port map( A => n286, B => n1732, C => n1957, Y => n1892);
   U91 : NAND2X1 port map( A => PLAINKEY_27_port, B => n285, Y => n1957);
   U93 : OAI21X1 port map( A => n285, B => n1731, C => n1956, Y => n1891);
   U94 : NAND2X1 port map( A => PLAINKEY_28_port, B => n284, Y => n1956);
   U96 : OAI21X1 port map( A => n286, B => n1730, C => n1955, Y => n1890);
   U97 : NAND2X1 port map( A => PLAINKEY_29_port, B => n284, Y => n1955);
   U99 : OAI21X1 port map( A => n286, B => n1729, C => n1954, Y => n1889);
   U100 : NAND2X1 port map( A => PLAINKEY_30_port, B => RST, Y => n1954);
   U102 : OAI21X1 port map( A => n287, B => n1728, C => n1953, Y => n1888);
   U103 : NAND2X1 port map( A => PLAINKEY_31_port, B => n288, Y => n1953);
   U105 : OAI21X1 port map( A => n287, B => n1727, C => n1952, Y => n1887);
   U106 : NAND2X1 port map( A => PLAINKEY_32_port, B => n286, Y => n1952);
   U108 : OAI21X1 port map( A => n286, B => n1726, C => n1951, Y => n1886);
   U109 : NAND2X1 port map( A => PLAINKEY_33_port, B => n287, Y => n1951);
   U111 : OAI21X1 port map( A => n287, B => n1725, C => n1950, Y => n1885);
   U112 : NAND2X1 port map( A => PLAINKEY_34_port, B => n285, Y => n1950);
   U114 : OAI21X1 port map( A => n286, B => n1724, C => n1949, Y => n1884);
   U115 : NAND2X1 port map( A => PLAINKEY_35_port, B => n284, Y => n1949);
   U117 : OAI21X1 port map( A => n286, B => n1723, C => n1948, Y => n1883);
   U118 : NAND2X1 port map( A => PLAINKEY_36_port, B => RST, Y => n1948);
   U120 : OAI21X1 port map( A => n287, B => n1722, C => n1947, Y => n1882);
   U121 : NAND2X1 port map( A => PLAINKEY_37_port, B => n286, Y => n1947);
   U123 : OAI21X1 port map( A => n287, B => n1721, C => n1946, Y => n1881);
   U124 : NAND2X1 port map( A => PLAINKEY_38_port, B => RST, Y => n1946);
   U126 : OAI21X1 port map( A => n287, B => n1720, C => n1945, Y => n1880);
   U127 : NAND2X1 port map( A => PLAINKEY_39_port, B => n288, Y => n1945);
   U129 : OAI21X1 port map( A => n287, B => n1719, C => n1944, Y => n1879);
   U130 : NAND2X1 port map( A => PLAINKEY_40_port, B => RST, Y => n1944);
   U132 : OAI21X1 port map( A => n287, B => n1718, C => n1943, Y => n1878);
   U133 : NAND2X1 port map( A => PLAINKEY_41_port, B => n287, Y => n1943);
   U135 : OAI21X1 port map( A => n286, B => n1717, C => n1942, Y => n1877);
   U136 : NAND2X1 port map( A => PLAINKEY_42_port, B => n285, Y => n1942);
   U138 : OAI21X1 port map( A => n287, B => n1716, C => n1941, Y => n1876);
   U139 : NAND2X1 port map( A => PLAINKEY_43_port, B => n286, Y => n1941);
   U141 : OAI21X1 port map( A => n287, B => n1715, C => n1940, Y => n1875);
   U142 : NAND2X1 port map( A => PLAINKEY_44_port, B => n287, Y => n1940);
   U144 : OAI21X1 port map( A => n287, B => n1714, C => n1939, Y => n1874);
   U145 : NAND2X1 port map( A => PLAINKEY_45_port, B => n284, Y => n1939);
   U147 : OAI21X1 port map( A => n287, B => n1713, C => n1938, Y => n1873);
   U148 : NAND2X1 port map( A => PLAINKEY_46_port, B => RST, Y => n1938);
   U150 : OAI21X1 port map( A => n284, B => n1712, C => n1937, Y => n1872);
   U151 : NAND2X1 port map( A => PLAINKEY_47_port, B => n287, Y => n1937);
   U153 : OAI21X1 port map( A => n286, B => n1711, C => n1936, Y => n1871);
   U154 : NAND2X1 port map( A => PLAINKEY_48_port, B => n285, Y => n1936);
   U156 : OAI21X1 port map( A => n286, B => n1710, C => n1935, Y => n1870);
   U157 : NAND2X1 port map( A => PLAINKEY_49_port, B => n287, Y => n1935);
   U159 : OAI21X1 port map( A => n286, B => n1709, C => n1934, Y => n1869);
   U160 : NAND2X1 port map( A => PLAINKEY_50_port, B => n284, Y => n1934);
   U162 : OAI21X1 port map( A => n285, B => n1708, C => n1933, Y => n1868);
   U163 : NAND2X1 port map( A => PLAINKEY_51_port, B => n286, Y => n1933);
   U165 : OAI21X1 port map( A => n286, B => n1707, C => n1932, Y => n1867);
   U166 : NAND2X1 port map( A => PLAINKEY_52_port, B => RST, Y => n1932);
   U168 : OAI21X1 port map( A => n285, B => n1706, C => n1931, Y => n1866);
   U169 : NAND2X1 port map( A => PLAINKEY_53_port, B => n285, Y => n1931);
   U171 : OAI21X1 port map( A => n285, B => n1705, C => n1930, Y => n1865);
   U172 : NAND2X1 port map( A => PLAINKEY_54_port, B => n286, Y => n1930);
   U174 : OAI21X1 port map( A => n284, B => n1704, C => n1929, Y => n1864);
   U175 : NAND2X1 port map( A => PLAINKEY_55_port, B => n287, Y => n1929);
   U177 : OAI21X1 port map( A => n285, B => n1703, C => n1928, Y => n1863);
   U178 : NAND2X1 port map( A => PLAINKEY_56_port, B => RST, Y => n1928);
   U180 : OAI21X1 port map( A => n284, B => n1702, C => n1927, Y => n1862);
   U181 : NAND2X1 port map( A => PLAINKEY_57_port, B => n288, Y => n1927);
   U183 : OAI21X1 port map( A => n284, B => n1701, C => n1926, Y => n1861);
   U184 : NAND2X1 port map( A => PLAINKEY_58_port, B => n285, Y => n1926);
   U186 : OAI21X1 port map( A => n284, B => n1700, C => n1925, Y => n1860);
   U187 : NAND2X1 port map( A => PLAINKEY_59_port, B => n287, Y => n1925);
   U188 : OAI21X1 port map( A => RST, B => n1699, C => n1924, Y => n1859);
   U189 : NAND2X1 port map( A => PLAINKEY_60_port, B => n285, Y => n1924);
   U191 : OAI21X1 port map( A => RST, B => n1698, C => n1923, Y => n1858);
   U192 : NAND2X1 port map( A => PLAINKEY_61_port, B => n288, Y => n1923);
   U194 : OAI21X1 port map( A => n288, B => n1685, C => n1922, Y => n1857);
   U195 : NAND2X1 port map( A => PLAINKEY_62_port, B => n284, Y => n1922);
   U196 : OAI21X1 port map( A => n286, B => n1697, C => n1921, Y => n1856);
   U197 : NAND2X1 port map( A => PLAINKEY_63_port, B => n284, Y => n1921);
   U1305 : NAND2X1 port map( A => n1648, B => n1760, Y => n1920);
   n1855 <= '1';
   n1854 <= '1';
   n1853 <= '1';
   n1852 <= '1';
   n1851 <= '1';
   n1850 <= '1';
   r577 : keyreg_0_DW01_add_1 port map( A(7) => parityAccumulator_7_port, A(6) 
                           => parityAccumulator_6_port, A(5) => 
                           parityAccumulator_5_port, A(4) => 
                           parityAccumulator_4_port, A(3) => 
                           parityAccumulator_3_port, A(2) => 
                           parityAccumulator_2_port, A(1) => 
                           parityAccumulator_1_port, A(0) => 
                           parityAccumulator_0_port, B(7) => RCV_DATA(7), B(6) 
                           => RCV_DATA(6), B(5) => RCV_DATA(5), B(4) => 
                           RCV_DATA(4), B(3) => RCV_DATA(3), B(2) => n281, B(1)
                           => RCV_DATA(1), B(0) => n220, CI => n1989, SUM(7) =>
                           N1799, SUM(6) => N1798, SUM(5) => N1797, SUM(4) => 
                           N1796, SUM(3) => N1795, SUM(2) => N1794, SUM(1) => 
                           N1793, SUM(0) => N1792, CO => n_1020);
   U3 : INVX2 port map( A => n747, Y => n678);
   U4 : INVX1 port map( A => n135, Y => n1163);
   U5 : INVX1 port map( A => n137, Y => n849);
   U7 : INVX2 port map( A => n849, Y => n785);
   U8 : INVX2 port map( A => n164, Y => n303);
   U23 : INVX4 port map( A => n67, Y => n177);
   U26 : INVX2 port map( A => n1372, Y => n1520);
   U29 : BUFX2 port map( A => n550, Y => n53);
   U32 : INVX1 port map( A => n691, Y => n103);
   U35 : INVX1 port map( A => n968, Y => n152);
   U38 : INVX1 port map( A => n1039, Y => n107);
   U41 : BUFX2 port map( A => n190, Y => n277);
   U44 : INVX4 port map( A => n163, Y => n164);
   U47 : INVX2 port map( A => n1021, Y => n1051);
   U50 : INVX2 port map( A => n1480, Y => n1437);
   U53 : INVX2 port map( A => n744, Y => n774);
   U56 : INVX1 port map( A => n205, Y => n206);
   U59 : INVX2 port map( A => n1542, Y => n205);
   U62 : AND2X1 port map( A => n188, B => n221, Y => n1);
   U65 : INVX2 port map( A => n847, Y => n824);
   U68 : AND2X2 port map( A => n312, B => n727, Y => n2);
   U71 : INVX2 port map( A => n637, Y => n614);
   U74 : INVX2 port map( A => n604, Y => n585);
   U77 : INVX2 port map( A => n1481, Y => n1444);
   U80 : INVX2 port map( A => n201, Y => n202);
   U83 : INVX2 port map( A => n1506, Y => n201);
   U86 : INVX2 port map( A => n1122, Y => n1105);
   U89 : INVX1 port map( A => n283, Y => n282);
   U92 : INVX1 port map( A => n1372, Y => n69);
   U95 : INVX4 port map( A => n117, Y => n275);
   U98 : INVX2 port map( A => n916, Y => n892);
   U101 : AND2X1 port map( A => n1462, B => n1464, Y => n4);
   U104 : INVX1 port map( A => n1515, Y => n5);
   U107 : INVX1 port map( A => n946, Y => n6);
   U110 : BUFX2 port map( A => n1504, Y => n7);
   U113 : BUFX2 port map( A => n413, Y => n8);
   U116 : INVX1 port map( A => n1155, Y => n9);
   U119 : INVX2 port map( A => n1121, Y => n1155);
   U122 : INVX1 port map( A => n1190, Y => n10);
   U125 : INVX1 port map( A => n910, Y => n11);
   U128 : NAND2X1 port map( A => n1660, B => n319, Y => n14);
   U131 : INVX4 port map( A => n197, Y => n1660);
   U134 : BUFX4 port map( A => n1482, Y => n251);
   U137 : BUFX4 port map( A => n1466, Y => n16);
   U140 : OR2X2 port map( A => n1529, B => n111, Y => n17);
   U143 : INVX1 port map( A => n17, Y => n115);
   U146 : INVX1 port map( A => n632, Y => n19);
   U149 : INVX2 port map( A => n1364, Y => n20);
   U152 : INVX1 port map( A => n1460, Y => n21);
   U155 : INVX2 port map( A => n1651, Y => n23);
   U158 : INVX2 port map( A => n648, Y => n25);
   U161 : INVX2 port map( A => n1444, Y => n27);
   U164 : INVX4 port map( A => n739, Y => n29);
   U167 : INVX2 port map( A => n708, Y => n739);
   U170 : INVX4 port map( A => n841, Y => n31);
   U173 : INVX2 port map( A => n814, Y => n841);
   U176 : INVX4 port map( A => n1016, Y => n33);
   U179 : INVX2 port map( A => n985, Y => n1016);
   U182 : BUFX2 port map( A => n1602, Y => n35);
   U185 : INVX4 port map( A => n809, Y => n37);
   U190 : INVX2 port map( A => n779, Y => n809);
   U193 : INVX4 port map( A => n1084, Y => n39);
   U198 : INVX2 port map( A => n1056, Y => n1084);
   U199 : INVX1 port map( A => n980, Y => n41);
   U200 : INVX2 port map( A => n1407, Y => n43);
   U201 : INVX2 port map( A => n926, Y => n45);
   U202 : INVX1 port map( A => n952, Y => n926);
   U203 : AND2X2 port map( A => n49, B => n327, Y => n47);
   U204 : INVX1 port map( A => n47, Y => n1142);
   U205 : NOR2X1 port map( A => address_1_port, B => address_0_port, Y => n49);
   U206 : INVX1 port map( A => n1419, Y => n51);
   U207 : INVX1 port map( A => n703, Y => n55);
   U208 : BUFX2 port map( A => n567, Y => n57);
   U209 : INVX1 port map( A => n1384, Y => n59);
   U210 : INVX2 port map( A => n1195, Y => n1384);
   U211 : INVX2 port map( A => n1557, Y => n61);
   U212 : INVX4 port map( A => n1578, Y => n1557);
   U213 : INVX4 port map( A => n1571, Y => n63);
   U214 : INVX4 port map( A => n1503, Y => n1571);
   U215 : INVX2 port map( A => n1437, Y => n65);
   U216 : INVX1 port map( A => address_0_port, Y => n324);
   U217 : OR2X2 port map( A => n335, B => n222, Y => n67);
   U218 : INVX2 port map( A => n335, Y => n586);
   U219 : INVX2 port map( A => n1424, Y => n1460);
   U220 : INVX1 port map( A => n69, Y => n71);
   U221 : INVX2 port map( A => n603, Y => n632);
   U222 : AND2X2 port map( A => n604, B => n603, Y => n123);
   U223 : INVX2 port map( A => n1176, Y => n73);
   U224 : INVX1 port map( A => n73, Y => n75);
   U225 : INVX2 port map( A => n189, Y => n77);
   U226 : INVX4 port map( A => n77, Y => n79);
   U227 : BUFX2 port map( A => n131, Y => n81);
   U228 : INVX4 port map( A => n562, Y => n83);
   U229 : INVX4 port map( A => n545, Y => n562);
   U230 : MUX2X1 port map( B => n271, A => n1489, S => n1524, Y => n1490);
   U231 : INVX1 port map( A => n1524, Y => n1596);
   U232 : BUFX2 port map( A => n125, Y => n85);
   U233 : INVX4 port map( A => n497, Y => n87);
   U234 : INVX4 port map( A => n478, Y => n497);
   U235 : INVX1 port map( A => n1175, Y => n89);
   U236 : NAND2X1 port map( A => n1463, B => n4, Y => n1842);
   U237 : AND2X2 port map( A => n916, B => n915, Y => n149);
   U238 : MUX2X1 port map( B => n283, A => n1491, S => n1529, Y => n1492);
   U239 : INVX1 port map( A => n1529, Y => n1598);
   U240 : BUFX2 port map( A => n174, Y => n91);
   U241 : INVX1 port map( A => n863, Y => n93);
   U242 : INVX1 port map( A => n125, Y => n457);
   U243 : INVX2 port map( A => n1160, Y => n1190);
   U244 : AND2X2 port map( A => n1090, B => n1089, Y => n95);
   U245 : INVX1 port map( A => n95, Y => n1092);
   U246 : INVX2 port map( A => n1092, Y => n1102);
   U247 : BUFX2 port map( A => n73, Y => n159);
   U248 : INVX2 port map( A => n881, Y => n910);
   U249 : AND2X1 port map( A => n745, B => n744, Y => n97);
   U250 : INVX1 port map( A => n97, Y => n747);
   U251 : AND2X1 port map( A => n1022, B => n1021, Y => n99);
   U252 : INVX1 port map( A => n99, Y => n1024);
   U253 : INVX2 port map( A => n1024, Y => n1036);
   U254 : INVX2 port map( A => n585, Y => n101);
   U255 : MUX2X1 port map( B => n262, A => n665, S => n103, Y => n667);
   U256 : BUFX2 port map( A => address_2_port, Y => n105);
   U257 : AND2X2 port map( A => n1196, B => n1195, Y => n154);
   U258 : INVX1 port map( A => n37, Y => n756);
   U259 : MUX2X1 port map( B => n261, A => n1013, S => n107, Y => n1015);
   U260 : INVX1 port map( A => n29, Y => n684);
   U261 : NAND2X1 port map( A => n299, B => n109, Y => n1664);
   U262 : AND2X1 port map( A => n226, B => n164, Y => n109);
   U263 : OR2X2 port map( A => n1529, B => n271, Y => n113);
   U264 : INVX1 port map( A => n168, Y => n111);
   U265 : AND2X2 port map( A => RCV_DATA(6), B => n228, Y => n117);
   U266 : INVX2 port map( A => n672, Y => n703);
   U267 : AND2X2 port map( A => n479, B => n478, Y => n125);
   U268 : INVX2 port map( A => n888, Y => n1141);
   U269 : INVX2 port map( A => n951, Y => n980);
   U270 : AND2X2 port map( A => n1465, B => n1453, Y => n119);
   U271 : INVX1 port map( A => n119, Y => n1493);
   U272 : BUFX4 port map( A => n1577, Y => n266);
   U273 : BUFX2 port map( A => n450, Y => n121);
   U274 : INVX2 port map( A => n1389, Y => n1419);
   U275 : INVX2 port map( A => n782, Y => n753);
   U276 : INVX2 port map( A => n711, Y => n681);
   U277 : INVX1 port map( A => n123, Y => n606);
   U278 : AND2X2 port map( A => n673, B => n672, Y => n141);
   U279 : INVX2 port map( A => n673, Y => n656);
   U280 : INVX1 port map( A => n39, Y => n1032);
   U281 : INVX1 port map( A => n1059, Y => n993);
   U282 : BUFX2 port map( A => n14, Y => n230);
   U283 : INVX1 port map( A => n988, Y => n921);
   U284 : AND2X1 port map( A => n1122, B => n1121, Y => n127);
   U285 : INVX2 port map( A => n127, Y => n1124);
   U286 : INVX2 port map( A => n1124, Y => n1137);
   U287 : BUFX4 port map( A => n190, Y => n280);
   U288 : OR2X2 port map( A => n166, B => n1644, Y => n1613);
   U289 : INVX2 port map( A => n166, Y => n1609);
   U290 : INVX2 port map( A => state_0_port, Y => n163);
   U291 : OR2X2 port map( A => n230, B => n283, Y => n1466);
   U292 : AND2X2 port map( A => n1425, B => n1424, Y => n129);
   U293 : INVX2 port map( A => n129, Y => n1427);
   U294 : INVX2 port map( A => n1427, Y => n1441);
   U295 : AND2X2 port map( A => n546, B => n545, Y => n131);
   U296 : INVX1 port map( A => n131, Y => n524);
   U297 : INVX4 port map( A => n155, Y => n169);
   U298 : AND2X2 port map( A => n513, B => n512, Y => n133);
   U299 : INVX1 port map( A => n133, Y => n491);
   U300 : AND2X2 port map( A => n1161, B => n1160, Y => n135);
   U301 : AND2X1 port map( A => n847, B => n846, Y => n137);
   U302 : AND2X2 port map( A => n882, B => n881, Y => n139);
   U303 : INVX2 port map( A => n139, Y => n884);
   U304 : INVX2 port map( A => n884, Y => n896);
   U305 : BUFX4 port map( A => n184, Y => n242);
   U306 : BUFX4 port map( A => n1428, Y => n231);
   U307 : INVX2 port map( A => n141, Y => n675);
   U308 : INVX2 port map( A => n675, Y => n688);
   U309 : BUFX4 port map( A => n184, Y => n243);
   U310 : INVX8 port map( A => n243, Y => n240);
   U311 : INVX1 port map( A => n1551, Y => n143);
   U312 : INVX2 port map( A => n1519, Y => n1551);
   U313 : AND2X2 port map( A => n1390, B => n1389, Y => n145);
   U314 : INVX2 port map( A => n145, Y => n1392);
   U315 : INVX2 port map( A => n1392, Y => n1404);
   U316 : AND2X2 port map( A => n1481, B => n1480, Y => n147);
   U317 : INVX1 port map( A => n147, Y => n1454);
   U318 : BUFX4 port map( A => n1482, Y => n249);
   U319 : INVX4 port map( A => n181, Y => n264);
   U320 : INVX2 port map( A => n264, Y => n263);
   U321 : BUFX4 port map( A => n184, Y => n245);
   U322 : INVX2 port map( A => n149, Y => n918);
   U323 : INVX2 port map( A => n918, Y => n931);
   U324 : AND2X1 port map( A => n638, B => n637, Y => n150);
   U325 : INVX1 port map( A => n150, Y => n640);
   U326 : INVX2 port map( A => n640, Y => n653);
   U327 : INVX4 port map( A => n117, Y => n276);
   U328 : INVX4 port map( A => n256, Y => n253);
   U329 : INVX1 port map( A => n328, Y => n151);
   U330 : INVX8 port map( A => n249, Y => n248);
   U331 : MUX2X1 port map( B => n261, A => n943, S => n152, Y => n945);
   U332 : INVX1 port map( A => n568, Y => n550);
   U333 : AND2X1 port map( A => n952, B => n951, Y => n153);
   U334 : INVX1 port map( A => n153, Y => n954);
   U335 : INVX2 port map( A => n954, Y => n965);
   U336 : INVX1 port map( A => n673, Y => n648);
   U337 : INVX1 port map( A => n154, Y => n1268);
   U338 : INVX2 port map( A => n1268, Y => n1368);
   U339 : INVX4 port map( A => n161, Y => n182);
   U340 : INVX1 port map( A => n1390, Y => n1364);
   U341 : INVX8 port map( A => n244, Y => n239);
   U342 : INVX8 port map( A => n249, Y => n247);
   U343 : INVX4 port map( A => n256, Y => n254);
   U344 : BUFX4 port map( A => n1466, Y => n238);
   U345 : INVX1 port map( A => n224, Y => n306);
   U346 : OR2X2 port map( A => n1582, B => n222, Y => n155);
   U347 : INVX2 port map( A => n1582, Y => n1561);
   U348 : MUX2X1 port map( B => n247, A => n1052, S => n1021, Y => n1054);
   U349 : NAND2X1 port map( A => n1660, B => n319, Y => n156);
   U350 : INVX4 port map( A => n191, Y => n204);
   U351 : AND2X2 port map( A => address_1_port, B => address_2_port, Y => n194)
                           ;
   U352 : AND2X2 port map( A => n1520, B => n223, Y => n157);
   U353 : BUFX2 port map( A => n864, Y => n158);
   U354 : INVX2 port map( A => n610, Y => n864);
   U355 : INVX1 port map( A => address_6_port, Y => n1696);
   U356 : INVX1 port map( A => n1453, Y => n1534);
   U357 : INVX1 port map( A => n782, Y => n716);
   U358 : INVX1 port map( A => n31, Y => n791);
   U359 : INVX1 port map( A => n817, Y => n750);
   U360 : INVX8 port map( A => n250, Y => n246);
   U361 : INVX1 port map( A => n711, Y => n643);
   U362 : INVX4 port map( A => n258, Y => n256);
   U363 : INVX2 port map( A => n256, Y => n255);
   U364 : INVX1 port map( A => n55, Y => n649);
   U365 : BUFX2 port map( A => address_0_port, Y => n160);
   U366 : OR2X2 port map( A => n888, B => n222, Y => n161);
   U367 : BUFX2 port map( A => n1520, Y => n162);
   U368 : INVX2 port map( A => n1612, Y => n165);
   U369 : INVX4 port map( A => n165, Y => n166);
   U370 : INVX4 port map( A => n265, Y => n262);
   U371 : INVX4 port map( A => n265, Y => n261);
   U372 : BUFX4 port map( A => n1466, Y => n237);
   U373 : INVX1 port map( A => n21, Y => n1400);
   U374 : INVX1 port map( A => n41, Y => n927);
   U375 : INVX4 port map( A => n264, Y => n260);
   U376 : INVX1 port map( A => n1664, Y => n1651);
   U377 : INVX1 port map( A => n245, Y => n167);
   U378 : INVX2 port map( A => n264, Y => n259);
   U379 : INVX1 port map( A => n172, Y => n235);
   U380 : BUFX4 port map( A => n184, Y => n244);
   U381 : INVX4 port map( A => n257, Y => n252);
   U382 : INVX4 port map( A => n283, Y => n281);
   U383 : INVX2 port map( A => n1505, Y => n258);
   U384 : INVX2 port map( A => n1584, Y => n274);
   U385 : INVX2 port map( A => address_3_port, Y => n221);
   U386 : INVX2 port map( A => n290, Y => n286);
   U387 : INVX2 port map( A => n290, Y => n285);
   U388 : INVX2 port map( A => n289, Y => n284);
   U389 : INVX2 port map( A => n291, Y => n287);
   U390 : INVX2 port map( A => n291, Y => n288);
   U391 : AND2X2 port map( A => n1468, B => n228, Y => n168);
   U392 : BUFX2 port map( A => n293, Y => n291);
   U393 : BUFX2 port map( A => n293, Y => n290);
   U394 : BUFX2 port map( A => n293, Y => n289);
   U395 : BUFX2 port map( A => n289, Y => n292);
   U396 : BUFX2 port map( A => n1577, Y => n267);
   U397 : BUFX2 port map( A => n1577, Y => n269);
   U398 : INVX4 port map( A => n156, Y => n229);
   U399 : INVX4 port map( A => n232, Y => n227);
   U400 : INVX2 port map( A => n172, Y => n233);
   U401 : INVX2 port map( A => n172, Y => n234);
   U402 : AND2X2 port map( A => n176, B => n1561, Y => n170);
   U403 : BUFX2 port map( A => n1577, Y => n270);
   U404 : INVX2 port map( A => n242, Y => n241);
   U405 : INVX2 port map( A => RST, Y => n293);
   U406 : AND2X2 port map( A => n325, B => n176, Y => n171);
   U407 : AND2X2 port map( A => n403, B => n185, Y => n172);
   U408 : AND2X2 port map( A => n1520, B => n223, Y => n173);
   U409 : AND2X2 port map( A => n73, B => n223, Y => n174);
   U410 : AND2X2 port map( A => n201, B => n223, Y => n175);
   U411 : AND2X2 port map( A => n205, B => n223, Y => n176);
   U412 : INVX2 port map( A => n181, Y => n265);
   U413 : AND2X2 port map( A => n223, B => n47, Y => n178);
   U414 : AND2X2 port map( A => n191, B => n223, Y => n179);
   U415 : INVX2 port map( A => n207, Y => n208);
   U416 : INVX2 port map( A => n207, Y => n209);
   U417 : AND2X2 port map( A => n325, B => n91, Y => n180);
   U418 : INVX2 port map( A => n571, Y => n207);
   U419 : BUFX2 port map( A => n190, Y => n278);
   U420 : BUFX2 port map( A => n190, Y => n279);
   U421 : AND2X2 port map( A => n343, B => n185, Y => n181);
   U422 : INVX2 port map( A => n274, Y => n272);
   U423 : INVX2 port map( A => n274, Y => n271);
   U424 : INVX2 port map( A => n1, Y => n218);
   U425 : AND2X2 port map( A => n864, B => n221, Y => n183);
   U426 : AND2X2 port map( A => n339, B => n185, Y => n184);
   U427 : AND2X2 port map( A => n319, B => n309, Y => n185);
   U428 : INVX2 port map( A => n258, Y => n257);
   U429 : AND2X2 port map( A => n194, B => n324, Y => n186);
   U430 : AND2X2 port map( A => n226, B => n225, Y => n187);
   U431 : INVX2 port map( A => n221, Y => n223);
   U432 : INVX2 port map( A => n274, Y => n273);
   U433 : INVX2 port map( A => n221, Y => n222);
   U434 : INVX2 port map( A => RCV_DATA(2), Y => n283);
   U435 : BUFX4 port map( A => state_2_port, Y => n225);
   U436 : BUFX4 port map( A => state_1_port, Y => n226);
   U437 : INVX2 port map( A => n210, Y => n211);
   U438 : INVX2 port map( A => n712, Y => n210);
   U439 : INVX2 port map( A => n214, Y => n215);
   U440 : INVX2 port map( A => n989, Y => n214);
   U441 : INVX4 port map( A => n212, Y => n213);
   U442 : INVX2 port map( A => n850, Y => n212);
   U443 : INVX4 port map( A => n216, Y => n217);
   U444 : INVX2 port map( A => n1125, Y => n216);
   U445 : INVX4 port map( A => n219, Y => n220);
   U446 : INVX2 port map( A => RCV_DATA(0), Y => n219);
   U447 : AND2X2 port map( A => address_4_port, B => address_5_port, Y => n188)
                           ;
   U448 : NOR2X1 port map( A => address_6_port, B => address_7_port, Y => n189)
                           ;
   U449 : AND2X2 port map( A => RCV_DATA(6), B => n228, Y => n190);
   U450 : AND2X2 port map( A => n194, B => n160, Y => n191);
   U451 : INVX4 port map( A => n2, Y => n203);
   U452 : NOR2X1 port map( A => n224, B => n164, Y => n192);
   U453 : NOR2X1 port map( A => n226, B => n164, Y => n193);
   U454 : INVX2 port map( A => n1469, Y => n195);
   U455 : INVX1 port map( A => n195, Y => n196);
   U456 : BUFX4 port map( A => n1672, Y => n197);
   U457 : BUFX2 port map( A => n1672, Y => n198);
   U458 : INVX1 port map( A => n186, Y => n199);
   U459 : INVX1 port map( A => n186, Y => n200);
   U460 : BUFX4 port map( A => state_3_port, Y => n224);
   U461 : INVX1 port map( A => n166, Y => n1611);
   U462 : BUFX2 port map( A => n14, Y => n232);
   U463 : INVX8 port map( A => n231, Y => n228);
   U464 : BUFX4 port map( A => n1466, Y => n236);
   U465 : BUFX4 port map( A => n1482, Y => n250);
   U466 : BUFX4 port map( A => n1577, Y => n268);
   U467 : NOR2X1 port map( A => n224, B => n225, Y => n294);
   U468 : NAND3X1 port map( A => n226, B => n303, C => n294, Y => n1672);
   U469 : INVX2 port map( A => n226, Y => n297);
   U470 : NOR2X1 port map( A => n224, B => n297, Y => n295);
   U471 : NAND3X1 port map( A => n225, B => n164, C => n295, Y => n1642);
   U472 : NAND2X1 port map( A => n197, B => n1642, Y => CLR_RBUFF_port);
   U473 : NOR2X1 port map( A => n224, B => n164, Y => n296);
   U474 : NAND3X1 port map( A => n225, B => n297, C => n296, Y => n1620);
   U475 : INVX2 port map( A => n1620, Y => PROG_ERROR);
   U476 : NOR2X1 port map( A => n226, B => n225, Y => n298);
   U477 : NAND2X1 port map( A => n298, B => n303, Y => n1662);
   U478 : NOR2X1 port map( A => n224, B => n225, Y => n299);
   U479 : OAI21X1 port map( A => n224, B => n1662, C => n1664, Y => n301);
   U480 : NAND2X1 port map( A => n187, B => n192, Y => n1661);
   U481 : NAND2X1 port map( A => n1661, B => n1620, Y => n300);
   U482 : NOR3X1 port map( A => CLR_RBUFF_port, B => n301, C => n300, Y => 
                           n1602);
   U483 : NOR2X1 port map( A => n225, B => n306, Y => n302);
   U484 : NAND2X1 port map( A => n302, B => n193, Y => n1663);
   U485 : NOR2X1 port map( A => n224, B => n303, Y => n304);
   U486 : NAND3X1 port map( A => n225, B => n297, C => n304, Y => n1669);
   U487 : INVX2 port map( A => n1669, Y => n1647);
   U488 : NOR2X1 port map( A => n226, B => n225, Y => n305);
   U489 : NAND3X1 port map( A => n164, B => n306, C => n305, Y => n1657);
   U490 : INVX2 port map( A => n1657, Y => n1615);
   U491 : AOI21X1 port map( A => n1647, B => parityError, C => n1615, Y => n307
                           );
   U492 : NAND3X1 port map( A => n35, B => n1663, C => n307, Y => KEY_ERROR);
   U493 : INVX2 port map( A => currentPlainKey_63_port, Y => n1697);
   U494 : INVX2 port map( A => currentPlainKey_62_port, Y => n1685);
   U495 : INVX2 port map( A => currentPlainKey_3_port, Y => n1756);
   U496 : INVX2 port map( A => currentPlainKey_2_port, Y => n1757);
   U497 : INVX2 port map( A => currentPlainKey_1_port, Y => n1758);
   U498 : INVX2 port map( A => currentPlainKey_0_port, Y => n1759);
   U499 : INVX2 port map( A => parityAccumulator_4_port, Y => n1692);
   U500 : INVX2 port map( A => parityAccumulator_5_port, Y => n1693);
   U501 : AOI21X1 port map( A => n187, B => n192, C => n287, Y => n308);
   U502 : AND2X2 port map( A => n308, B => n1664, Y => n319);
   U503 : AND2X2 port map( A => n1657, B => n1620, Y => n309);
   U504 : NAND3X1 port map( A => n1663, B => n1642, C => n185, Y => n310);
   U505 : INVX2 port map( A => n310, Y => n1683);
   U506 : NAND2X1 port map( A => n1683, B => n1669, Y => n1577);
   U507 : NAND2X1 port map( A => n270, B => currentPlainKey_0_port, Y => n333);
   U508 : NAND3X1 port map( A => address_6_port, B => address_7_port, C => n188
                           , Y => n329);
   U509 : INVX2 port map( A => n329, Y => n325);
   U510 : INVX2 port map( A => address_1_port, Y => n328);
   U511 : NAND3X1 port map( A => address_2_port, B => n324, C => n328, Y => 
                           n1372);
   U512 : NAND2X1 port map( A => n325, B => n173, Y => n311);
   U513 : INVX2 port map( A => n311, Y => n380);
   U514 : INVX2 port map( A => RCV_DATA(4), Y => n342);
   U515 : NAND2X1 port map( A => n380, B => n342, Y => n323);
   U516 : NAND2X1 port map( A => n186, B => n223, Y => n1581);
   U517 : INVX2 port map( A => n1581, Y => n1130);
   U518 : NAND2X1 port map( A => n325, B => n1130, Y => n412);
   U519 : INVX2 port map( A => n412, Y => n384);
   U520 : INVX2 port map( A => address_2_port, Y => n327);
   U521 : NAND3X1 port map( A => address_1_port, B => address_0_port, C => n327
                           , Y => n1506);
   U522 : NAND2X1 port map( A => n325, B => n175, Y => n345);
   U523 : NAND2X1 port map( A => n345, B => n311, Y => n361);
   U524 : AOI21X1 port map( A => n384, B => n281, C => n361, Y => n318);
   U525 : NOR2X1 port map( A => address_4_port, B => n222, Y => n312);
   U526 : INVX2 port map( A => address_5_port, Y => n727);
   U527 : INVX2 port map( A => n203, Y => n368);
   U528 : NAND2X1 port map( A => n368, B => n47, Y => n313);
   U529 : NAND2X1 port map( A => n220, B => n47, Y => n1144);
   U530 : INVX2 port map( A => n1144, Y => n1445);
   U531 : AOI22X1 port map( A => n313, B => currentPlainKey_0_port, C => n368, 
                           D => n1445, Y => n315);
   U532 : NAND2X1 port map( A => n325, B => n179, Y => n413);
   U533 : NAND2X1 port map( A => n412, B => n413, Y => n391);
   U534 : INVX2 port map( A => n413, Y => n430);
   U535 : NAND2X1 port map( A => n430, B => RCV_DATA(1), Y => n314);
   U536 : OAI21X1 port map( A => n315, B => n391, C => n314, Y => n316);
   U537 : NAND3X1 port map( A => address_2_port, B => address_0_port, C => n328
                           , Y => n1542);
   U538 : MUX2X1 port map( B => n316, A => RCV_DATA(3), S => n171, Y => n317);
   U539 : NAND2X1 port map( A => n318, B => n317, Y => n322);
   U540 : NAND2X1 port map( A => n1660, B => n319, Y => n1428);
   U541 : NAND2X1 port map( A => n229, B => n345, Y => n320);
   U542 : NAND3X1 port map( A => n185, B => RCV_DATA(5), C => n1660, Y => n1505
                           );
   U543 : NAND2X1 port map( A => n320, B => n257, Y => n321);
   U544 : NAND3X1 port map( A => n323, B => n322, C => n321, Y => n326);
   U545 : NAND3X1 port map( A => address_1_port, B => n324, C => n327, Y => 
                           n1176);
   U546 : MUX2X1 port map( B => n326, A => n276, S => n180, Y => n331);
   U547 : NAND2X1 port map( A => RCV_DATA(7), B => n228, Y => n1482);
   U548 : NAND3X1 port map( A => n328, B => address_0_port, C => n327, Y => 
                           n1469);
   U549 : NAND2X1 port map( A => n195, B => n223, Y => n484);
   U550 : NOR2X1 port map( A => n484, B => n329, Y => n330);
   U551 : MUX2X1 port map( B => n331, A => n248, S => n330, Y => n332);
   U552 : NAND2X1 port map( A => n333, B => n332, Y => n1786);
   U553 : NAND2X1 port map( A => n270, B => currentPlainKey_1_port, Y => n350);
   U554 : INVX2 port map( A => n391, Y => n411);
   U555 : NAND2X1 port map( A => n368, B => n195, Y => n334);
   U556 : NAND2X1 port map( A => n220, B => n195, Y => n469);
   U557 : INVX2 port map( A => n469, Y => n1470);
   U558 : AOI22X1 port map( A => n334, B => currentPlainKey_1_port, C => n368, 
                           D => n1470, Y => n336);
   U559 : INVX2 port map( A => RCV_DATA(1), Y => n1584);
   U560 : INVX2 port map( A => address_4_port, Y => n1004);
   U561 : NAND3X1 port map( A => n79, B => n1004, C => n727, Y => n335);
   U562 : NAND2X1 port map( A => n177, B => n47, Y => n446);
   U563 : INVX2 port map( A => n446, Y => n417);
   U564 : MUX2X1 port map( B => n336, A => n271, S => n417, Y => n338);
   U565 : NOR2X1 port map( A => n283, B => n413, Y => n337);
   U566 : AOI21X1 port map( A => n411, B => n338, C => n337, Y => n341);
   U567 : INVX2 port map( A => RCV_DATA(3), Y => n1589);
   U568 : NOR2X1 port map( A => n1589, B => n198, Y => n339);
   U569 : NAND2X1 port map( A => n384, B => n245, Y => n340);
   U570 : OAI21X1 port map( A => n341, B => n230, C => n340, Y => n344);
   U571 : NOR2X1 port map( A => n342, B => n198, Y => n343);
   U572 : MUX2X1 port map( B => n344, A => n261, S => n171, Y => n347);
   U573 : INVX2 port map( A => n345, Y => n351);
   U574 : AOI22X1 port map( A => n380, B => n253, C => n351, D => n280, Y => 
                           n346);
   U575 : OAI21X1 port map( A => n347, B => n361, C => n346, Y => n348);
   U576 : MUX2X1 port map( B => n348, A => n247, S => n180, Y => n349);
   U577 : NAND2X1 port map( A => n350, B => n349, Y => n1787);
   U578 : AOI22X1 port map( A => n267, B => currentPlainKey_2_port, C => n351, 
                           D => n246, Y => n367);
   U579 : NOR2X1 port map( A => n265, B => n412, Y => n364);
   U580 : NOR2X1 port map( A => n241, B => n8, Y => n359);
   U581 : NAND2X1 port map( A => n417, B => n281, Y => n357);
   U582 : OAI21X1 port map( A => n75, B => n203, C => currentPlainKey_2_port, Y
                           => n353);
   U583 : NAND2X1 port map( A => n73, B => n220, Y => n1179);
   U584 : INVX2 port map( A => n1179, Y => n1486);
   U585 : NAND2X1 port map( A => n368, B => n1486, Y => n352);
   U586 : NAND2X1 port map( A => n177, B => n195, Y => n445);
   U587 : NAND2X1 port map( A => n446, B => n445, Y => n424);
   U588 : AOI21X1 port map( A => n353, B => n352, C => n424, Y => n355);
   U589 : INVX2 port map( A => n445, Y => n463);
   U590 : AND2X2 port map( A => n463, B => RCV_DATA(1), Y => n354);
   U591 : OAI21X1 port map( A => n355, B => n354, C => n8, Y => n356);
   U592 : AOI21X1 port map( A => n357, B => n356, C => n230, Y => n358);
   U593 : OAI21X1 port map( A => n359, B => n358, C => n412, Y => n360);
   U594 : MUX2X1 port map( B => n360, A => n257, S => n171, Y => n363);
   U595 : INVX2 port map( A => n361, Y => n362);
   U596 : OAI21X1 port map( A => n364, B => n363, C => n362, Y => n366);
   U597 : NAND2X1 port map( A => n380, B => n278, Y => n365);
   U598 : NAND3X1 port map( A => n367, B => n366, C => n365, Y => n1788);
   U599 : NAND2X1 port map( A => n269, B => currentPlainKey_3_port, Y => n383);
   U600 : NOR2X1 port map( A => n257, B => n412, Y => n378);
   U601 : OAI21X1 port map( A => n202, B => n203, C => currentPlainKey_3_port, 
                           Y => n370);
   U602 : NAND2X1 port map( A => n220, B => n201, Y => n503);
   U603 : INVX2 port map( A => n503, Y => n1357);
   U604 : NAND2X1 port map( A => n368, B => n1357, Y => n369);
   U605 : NAND2X1 port map( A => n370, B => n369, Y => n371);
   U606 : NAND2X1 port map( A => n177, B => n159, Y => n479);
   U607 : INVX2 port map( A => n479, Y => n450);
   U608 : MUX2X1 port map( B => n371, A => RCV_DATA(1), S => n450, Y => n373);
   U609 : NAND2X1 port map( A => n463, B => n282, Y => n372);
   U610 : OAI21X1 port map( A => n373, B => n424, C => n372, Y => n374);
   U611 : AOI22X1 port map( A => n417, B => n242, C => n374, D => n227, Y => 
                           n376);
   U612 : NAND2X1 port map( A => n430, B => n263, Y => n375);
   U613 : OAI21X1 port map( A => n376, B => n391, C => n375, Y => n377);
   U614 : NOR2X1 port map( A => n378, B => n377, Y => n379);
   U615 : MUX2X1 port map( B => n379, A => n276, S => n171, Y => n381);
   U616 : MUX2X1 port map( B => n381, A => n247, S => n380, Y => n382);
   U617 : NAND2X1 port map( A => n383, B => n382, Y => n1789);
   U618 : NAND2X1 port map( A => n384, B => n278, Y => n400);
   U619 : NAND2X1 port map( A => n177, B => n201, Y => n478);
   U620 : NAND2X1 port map( A => n220, B => n1520, Y => n1521);
   U621 : OAI21X1 port map( A => n71, B => n203, C => currentPlainKey_4_port, Y
                           => n385);
   U622 : OAI21X1 port map( A => n1521, B => n203, C => n385, Y => n387);
   U623 : NOR2X1 port map( A => n271, B => n87, Y => n386);
   U624 : AOI21X1 port map( A => n125, B => n387, C => n386, Y => n389);
   U625 : NAND2X1 port map( A => n450, B => n282, Y => n388);
   U626 : OAI21X1 port map( A => n463, B => n389, C => n388, Y => n390);
   U627 : NAND2X1 port map( A => n229, B => n390, Y => n393);
   U628 : NAND2X1 port map( A => n463, B => n245, Y => n392);
   U629 : AOI21X1 port map( A => n393, B => n392, C => n391, Y => n394);
   U630 : MUX2X1 port map( B => n394, A => n262, S => n417, Y => n396);
   U631 : NAND2X1 port map( A => n430, B => n254, Y => n395);
   U632 : NAND2X1 port map( A => n396, B => n395, Y => n397);
   U633 : MUX2X1 port map( B => n397, A => n247, S => n171, Y => n399);
   U634 : NAND2X1 port map( A => currentPlainKey_4_port, B => n266, Y => n398);
   U635 : NAND3X1 port map( A => n400, B => n399, C => n398, Y => n1790);
   U636 : NAND2X1 port map( A => n463, B => n263, Y => n409);
   U637 : NAND2X1 port map( A => n220, B => n205, Y => n1544);
   U638 : OAI21X1 port map( A => n206, B => n203, C => currentPlainKey_5_port, 
                           Y => n401);
   U639 : OAI21X1 port map( A => n1544, B => n203, C => n401, Y => n402);
   U640 : NAND3X1 port map( A => n125, B => n228, C => n402, Y => n404);
   U641 : NOR2X1 port map( A => n273, B => n198, Y => n403);
   U642 : NAND2X1 port map( A => n177, B => n162, Y => n513);
   U643 : INVX2 port map( A => n513, Y => n483);
   U644 : MUX2X1 port map( B => n404, A => n233, S => n483, Y => n406);
   U645 : OAI22X1 port map( A => n241, B => n479, C => n236, D => n87, Y => 
                           n405);
   U646 : INVX2 port map( A => n424, Y => n444);
   U647 : OAI21X1 port map( A => n406, B => n405, C => n444, Y => n408);
   U648 : NAND2X1 port map( A => n417, B => n254, Y => n407);
   U649 : NAND3X1 port map( A => n409, B => n408, C => n407, Y => n410);
   U650 : NAND2X1 port map( A => n411, B => n410, Y => n416);
   U651 : OAI22X1 port map( A => n276, B => n8, C => n251, D => n412, Y => n414
                           );
   U652 : AOI21X1 port map( A => currentPlainKey_5_port, B => n269, C => n414, 
                           Y => n415);
   U653 : NAND2X1 port map( A => n416, B => n415, Y => n1791);
   U654 : NAND2X1 port map( A => n417, B => n280, Y => n434);
   U655 : NAND2X1 port map( A => n177, B => n205, Y => n512);
   U656 : NAND2X1 port map( A => n220, B => n186, Y => n1556);
   U657 : OAI21X1 port map( A => n200, B => n203, C => currentPlainKey_6_port, 
                           Y => n418);
   U658 : OAI21X1 port map( A => n1556, B => n203, C => n418, Y => n420);
   U659 : NOR2X1 port map( A => n273, B => n512, Y => n419);
   U660 : AOI21X1 port map( A => n133, B => n420, C => n419, Y => n422);
   U661 : NAND2X1 port map( A => n483, B => n282, Y => n421);
   U662 : OAI21X1 port map( A => n497, B => n422, C => n421, Y => n423);
   U663 : NAND2X1 port map( A => n229, B => n423, Y => n426);
   U664 : NAND2X1 port map( A => n497, B => n245, Y => n425);
   U665 : AOI21X1 port map( A => n426, B => n425, C => n424, Y => n427);
   U666 : MUX2X1 port map( B => n427, A => n262, S => n121, Y => n429);
   U667 : NAND2X1 port map( A => n463, B => n254, Y => n428);
   U668 : NAND2X1 port map( A => n429, B => n428, Y => n431);
   U669 : MUX2X1 port map( B => n431, A => n246, S => n430, Y => n433);
   U670 : NAND2X1 port map( A => currentPlainKey_6_port, B => n268, Y => n432);
   U671 : NAND3X1 port map( A => n434, B => n433, C => n432, Y => n1792_port);
   U672 : NAND2X1 port map( A => n497, B => n263, Y => n442);
   U673 : NAND2X1 port map( A => n220, B => n191, Y => n572);
   U674 : OAI21X1 port map( A => n204, B => n203, C => currentPlainKey_7_port, 
                           Y => n435);
   U675 : OAI21X1 port map( A => n572, B => n203, C => n435, Y => n436);
   U676 : NAND3X1 port map( A => n133, B => n228, C => n436, Y => n437);
   U677 : NAND2X1 port map( A => n177, B => n186, Y => n546);
   U678 : INVX2 port map( A => n546, Y => n517);
   U679 : MUX2X1 port map( B => n437, A => n233, S => n517, Y => n439);
   U680 : OAI22X1 port map( A => n240, B => n513, C => n236, D => n512, Y => 
                           n438);
   U681 : OAI21X1 port map( A => n439, B => n438, C => n85, Y => n441);
   U682 : NAND2X1 port map( A => n121, B => n254, Y => n440);
   U683 : NAND3X1 port map( A => n442, B => n441, C => n440, Y => n443);
   U684 : NAND2X1 port map( A => n444, B => n443, Y => n449);
   U685 : OAI22X1 port map( A => n250, B => n446, C => n276, D => n445, Y => 
                           n447);
   U686 : AOI21X1 port map( A => currentPlainKey_7_port, B => n269, C => n447, 
                           Y => n448);
   U687 : NAND2X1 port map( A => n449, B => n448, Y => n1793_port);
   U688 : NAND2X1 port map( A => n121, B => n279, Y => n467);
   U689 : INVX2 port map( A => n512, Y => n530);
   U690 : NAND2X1 port map( A => n177, B => n191, Y => n545);
   U691 : NAND3X1 port map( A => n222, B => n1004, C => n727, Y => n571);
   U692 : OAI21X1 port map( A => n1142, B => n209, C => currentPlainKey_8_port,
                           Y => n451);
   U693 : OAI21X1 port map( A => n1144, B => n208, C => n451, Y => n453);
   U694 : NOR2X1 port map( A => n273, B => n83, Y => n452);
   U695 : AOI21X1 port map( A => n131, B => n453, C => n452, Y => n455);
   U696 : NAND2X1 port map( A => n517, B => n282, Y => n454);
   U697 : OAI21X1 port map( A => n530, B => n455, C => n454, Y => n456);
   U698 : NAND2X1 port map( A => n229, B => n456, Y => n459);
   U699 : NAND2X1 port map( A => n530, B => n245, Y => n458);
   U700 : AOI21X1 port map( A => n459, B => n458, C => n457, Y => n460);
   U701 : MUX2X1 port map( B => n460, A => n262, S => n483, Y => n462);
   U702 : NAND2X1 port map( A => n497, B => n255, Y => n461);
   U703 : NAND2X1 port map( A => n462, B => n461, Y => n464);
   U704 : MUX2X1 port map( B => n464, A => n246, S => n463, Y => n466);
   U705 : NAND2X1 port map( A => currentPlainKey_8_port, B => n266, Y => n465);
   U706 : NAND3X1 port map( A => n467, B => n466, C => n465, Y => n1794_port);
   U707 : NAND2X1 port map( A => n530, B => n263, Y => n476);
   U708 : OAI21X1 port map( A => n196, B => n209, C => currentPlainKey_9_port, 
                           Y => n468);
   U709 : OAI21X1 port map( A => n469, B => n208, C => n468, Y => n470);
   U710 : NAND3X1 port map( A => n131, B => n228, C => n470, Y => n471);
   U711 : NAND2X1 port map( A => n586, B => n178, Y => n568);
   U712 : MUX2X1 port map( B => n471, A => n233, S => n53, Y => n473);
   U713 : OAI22X1 port map( A => n240, B => n546, C => n238, D => n83, Y => 
                           n472);
   U714 : OAI21X1 port map( A => n473, B => n472, C => n133, Y => n475);
   U715 : NAND2X1 port map( A => n483, B => n255, Y => n474);
   U716 : NAND3X1 port map( A => n476, B => n475, C => n474, Y => n477);
   U717 : NAND2X1 port map( A => n85, B => n477, Y => n482);
   U718 : OAI22X1 port map( A => n251, B => n479, C => n275, D => n87, Y => 
                           n480);
   U719 : AOI21X1 port map( A => currentPlainKey_9_port, B => n266, C => n480, 
                           Y => n481);
   U720 : NAND2X1 port map( A => n481, B => n482, Y => n1795_port);
   U721 : NAND2X1 port map( A => n483, B => n277, Y => n501);
   U722 : INVX2 port map( A => n484, Y => n1488);
   U723 : NAND2X1 port map( A => n586, B => n1488, Y => n567);
   U724 : NAND2X1 port map( A => n568, B => n567, Y => n570);
   U725 : INVX2 port map( A => n570, Y => n538);
   U726 : OAI21X1 port map( A => n75, B => n209, C => currentPlainKey_10_port, 
                           Y => n485);
   U727 : OAI21X1 port map( A => n1179, B => n208, C => n485, Y => n487);
   U728 : NOR2X1 port map( A => n273, B => n567, Y => n486);
   U729 : AOI21X1 port map( A => n538, B => n487, C => n486, Y => n489);
   U730 : NAND2X1 port map( A => n550, B => n282, Y => n488);
   U731 : OAI21X1 port map( A => n562, B => n489, C => n488, Y => n490);
   U732 : NAND2X1 port map( A => n229, B => n490, Y => n493);
   U733 : NAND2X1 port map( A => n562, B => n245, Y => n492);
   U734 : AOI21X1 port map( A => n493, B => n492, C => n491, Y => n494);
   U735 : MUX2X1 port map( B => n494, A => n262, S => n517, Y => n496);
   U736 : NAND2X1 port map( A => n530, B => n255, Y => n495);
   U737 : NAND2X1 port map( A => n496, B => n495, Y => n498);
   U738 : MUX2X1 port map( B => n498, A => n246, S => n497, Y => n500);
   U739 : NAND2X1 port map( A => currentPlainKey_10_port, B => n266, Y => n499)
                           ;
   U740 : NAND3X1 port map( A => n501, B => n500, C => n499, Y => n1796_port);
   U741 : NAND2X1 port map( A => n562, B => n262, Y => n510);
   U742 : OAI21X1 port map( A => n202, B => n209, C => currentPlainKey_11_port,
                           Y => n502);
   U743 : OAI21X1 port map( A => n503, B => n208, C => n502, Y => n504);
   U744 : NAND3X1 port map( A => n538, B => n228, C => n504, Y => n505);
   U745 : NAND2X1 port map( A => n586, B => n174, Y => n604);
   U746 : MUX2X1 port map( B => n505, A => n233, S => n585, Y => n507);
   U747 : OAI22X1 port map( A => n240, B => n568, C => n236, D => n57, Y => 
                           n506);
   U748 : OAI21X1 port map( A => n507, B => n506, C => n81, Y => n509);
   U749 : NAND2X1 port map( A => n517, B => n253, Y => n508);
   U750 : NAND3X1 port map( A => n510, B => n509, C => n508, Y => n511);
   U751 : NAND2X1 port map( A => n133, B => n511, Y => n516);
   U752 : OAI22X1 port map( A => n249, B => n513, C => n276, D => n512, Y => 
                           n514);
   U753 : AOI21X1 port map( A => currentPlainKey_11_port, B => n268, C => n514,
                           Y => n515);
   U754 : NAND2X1 port map( A => n516, B => n515, Y => n1797_port);
   U755 : NAND2X1 port map( A => n517, B => n278, Y => n534);
   U756 : INVX2 port map( A => n567, Y => n598);
   U757 : NAND2X1 port map( A => n586, B => n175, Y => n603);
   U758 : OAI21X1 port map( A => n71, B => n209, C => currentPlainKey_12_port, 
                           Y => n518);
   U759 : OAI21X1 port map( A => n1521, B => n208, C => n518, Y => n520);
   U760 : NOR2X1 port map( A => n273, B => n603, Y => n519);
   U761 : AOI21X1 port map( A => n123, B => n520, C => n519, Y => n522);
   U762 : NAND2X1 port map( A => n585, B => n282, Y => n521);
   U763 : OAI21X1 port map( A => n522, B => n598, C => n521, Y => n523);
   U764 : NAND2X1 port map( A => n229, B => n523, Y => n526);
   U765 : NAND2X1 port map( A => n598, B => n245, Y => n525);
   U766 : AOI21X1 port map( A => n526, B => n525, C => n524, Y => n527);
   U767 : MUX2X1 port map( B => n527, A => n262, S => n53, Y => n529);
   U768 : NAND2X1 port map( A => n562, B => n255, Y => n528);
   U769 : NAND2X1 port map( A => n529, B => n528, Y => n531);
   U770 : MUX2X1 port map( B => n531, A => n246, S => n530, Y => n533);
   U771 : NAND2X1 port map( A => currentPlainKey_12_port, B => n270, Y => n532)
                           ;
   U772 : NAND3X1 port map( A => n534, B => n533, C => n532, Y => n1798_port);
   U773 : NAND2X1 port map( A => n598, B => n263, Y => n543);
   U774 : OAI21X1 port map( A => n206, B => n209, C => currentPlainKey_13_port,
                           Y => n535);
   U775 : OAI21X1 port map( A => n1544, B => n208, C => n535, Y => n536);
   U776 : NAND3X1 port map( A => n123, B => n228, C => n536, Y => n537);
   U777 : NAND2X1 port map( A => n586, B => n157, Y => n638);
   U778 : INVX2 port map( A => n638, Y => n620);
   U779 : MUX2X1 port map( B => n537, A => n233, S => n620, Y => n540);
   U780 : OAI22X1 port map( A => n240, B => n101, C => n16, D => n19, Y => n539
                           );
   U781 : OAI21X1 port map( A => n540, B => n539, C => n538, Y => n542);
   U782 : NAND2X1 port map( A => n53, B => n255, Y => n541);
   U783 : NAND3X1 port map( A => n543, B => n542, C => n541, Y => n544);
   U784 : NAND2X1 port map( A => n81, B => n544, Y => n549);
   U785 : OAI22X1 port map( A => n249, B => n546, C => n276, D => n83, Y => 
                           n547);
   U786 : AOI21X1 port map( A => currentPlainKey_13_port, B => n268, C => n547,
                           Y => n548);
   U787 : NAND2X1 port map( A => n548, B => n549, Y => n1799_port);
   U788 : NAND2X1 port map( A => n53, B => n279, Y => n566);
   U789 : NAND2X1 port map( A => n586, B => n176, Y => n637);
   U790 : OAI21X1 port map( A => n199, B => n209, C => currentPlainKey_14_port,
                           Y => n551);
   U791 : OAI21X1 port map( A => n1556, B => n208, C => n551, Y => n553);
   U792 : NOR2X1 port map( A => n272, B => n637, Y => n552);
   U793 : AOI21X1 port map( A => n150, B => n553, C => n552, Y => n555);
   U794 : NAND2X1 port map( A => n620, B => n282, Y => n554);
   U795 : OAI21X1 port map( A => n632, B => n555, C => n554, Y => n556);
   U796 : NAND2X1 port map( A => n229, B => n556, Y => n558);
   U797 : NAND2X1 port map( A => n632, B => n245, Y => n557);
   U798 : AOI21X1 port map( A => n558, B => n557, C => n570, Y => n559);
   U799 : MUX2X1 port map( B => n559, A => n262, S => n585, Y => n561);
   U800 : NAND2X1 port map( A => n598, B => n255, Y => n560);
   U801 : NAND2X1 port map( A => n561, B => n560, Y => n563);
   U802 : MUX2X1 port map( B => n563, A => n246, S => n562, Y => n565);
   U803 : NAND2X1 port map( A => currentPlainKey_14_port, B => n266, Y => n564)
                           ;
   U804 : NAND3X1 port map( A => n566, B => n565, C => n564, Y => n1800);
   U805 : OAI22X1 port map( A => n249, B => n568, C => n276, D => n57, Y => 
                           n569);
   U806 : AOI21X1 port map( A => currentPlainKey_15_port, B => n266, C => n569,
                           Y => n584);
   U807 : OAI21X1 port map( A => n204, B => n209, C => currentPlainKey_15_port,
                           Y => n575);
   U808 : INVX2 port map( A => n208, Y => n573);
   U809 : INVX2 port map( A => n572, Y => n1430);
   U810 : NAND2X1 port map( A => n573, B => n1430, Y => n574);
   U811 : NAND2X1 port map( A => n575, B => n574, Y => n576);
   U812 : NAND3X1 port map( A => n228, B => n576, C => n653, Y => n577);
   U813 : NAND2X1 port map( A => n586, B => n1130, Y => n673);
   U814 : MUX2X1 port map( B => n577, A => n233, S => n656, Y => n579);
   U815 : OAI22X1 port map( A => n240, B => n638, C => n16, D => n637, Y => 
                           n578);
   U816 : OAI21X1 port map( A => n579, B => n578, C => n123, Y => n581);
   U817 : AOI22X1 port map( A => n632, B => n260, C => n585, D => n253, Y => 
                           n580);
   U818 : NAND2X1 port map( A => n581, B => n580, Y => n582);
   U819 : NAND2X1 port map( A => n538, B => n582, Y => n583);
   U820 : NAND2X1 port map( A => n584, B => n583, Y => n1801);
   U821 : NAND2X1 port map( A => n585, B => n277, Y => n602);
   U822 : NAND2X1 port map( A => n586, B => n179, Y => n672);
   U823 : NAND3X1 port map( A => address_4_port, B => n221, C => n727, Y => 
                           n712);
   U824 : OAI21X1 port map( A => n1142, B => n211, C => currentPlainKey_16_port
                           , Y => n587);
   U825 : OAI21X1 port map( A => n1144, B => n211, C => n587, Y => n589);
   U826 : NOR2X1 port map( A => n272, B => n672, Y => n588);
   U827 : AOI21X1 port map( A => n141, B => n589, C => n588, Y => n591);
   U828 : NAND2X1 port map( A => n656, B => n282, Y => n590);
   U829 : OAI21X1 port map( A => n614, B => n591, C => n590, Y => n592);
   U830 : NAND2X1 port map( A => n229, B => n592, Y => n594);
   U831 : NAND2X1 port map( A => n614, B => n245, Y => n593);
   U832 : AOI21X1 port map( A => n594, B => n593, C => n606, Y => n595);
   U833 : MUX2X1 port map( B => n595, A => n262, S => n620, Y => n597);
   U834 : NAND2X1 port map( A => n632, B => n255, Y => n596);
   U835 : NAND2X1 port map( A => n597, B => n596, Y => n599);
   U836 : MUX2X1 port map( B => n599, A => n246, S => n598, Y => n601);
   U837 : NAND2X1 port map( A => currentPlainKey_16_port, B => n268, Y => n600)
                           ;
   U838 : NAND3X1 port map( A => n602, B => n601, C => n600, Y => n1802);
   U839 : OAI22X1 port map( A => n250, B => n101, C => n276, D => n19, Y => 
                           n605);
   U840 : AOI21X1 port map( A => currentPlainKey_17_port, B => n266, C => n605,
                           Y => n619);
   U841 : OAI21X1 port map( A => n196, B => n211, C => currentPlainKey_17_port,
                           Y => n608);
   U842 : INVX2 port map( A => n211, Y => n713);
   U843 : NAND2X1 port map( A => n713, B => n1470, Y => n607);
   U844 : NAND2X1 port map( A => n608, B => n607, Y => n609);
   U845 : NAND3X1 port map( A => n227, B => n609, C => n688, Y => n611);
   U846 : NAND3X1 port map( A => n79, B => address_4_port, C => n727, Y => n610
                           );
   U847 : NAND2X1 port map( A => n183, B => n47, Y => n709);
   U848 : INVX2 port map( A => n709, Y => n691);
   U849 : MUX2X1 port map( B => n611, A => n233, S => n691, Y => n613);
   U850 : OAI22X1 port map( A => n240, B => n25, C => n238, D => n55, Y => n612
                           );
   U851 : OAI21X1 port map( A => n613, B => n612, C => n653, Y => n616);
   U852 : AOI22X1 port map( A => n614, B => n260, C => n620, D => n253, Y => 
                           n615);
   U853 : NAND2X1 port map( A => n616, B => n615, Y => n617);
   U854 : NAND2X1 port map( A => n123, B => n617, Y => n618);
   U855 : NAND2X1 port map( A => n619, B => n618, Y => n1803);
   U856 : NAND2X1 port map( A => n620, B => n279, Y => n636);
   U857 : NAND2X1 port map( A => n183, B => n195, Y => n708);
   U858 : NAND2X1 port map( A => n709, B => n708, Y => n711);
   U859 : OAI21X1 port map( A => n75, B => n211, C => currentPlainKey_18_port, 
                           Y => n621);
   U860 : OAI21X1 port map( A => n1179, B => n211, C => n621, Y => n623);
   U861 : NOR2X1 port map( A => n272, B => n29, Y => n622);
   U862 : AOI21X1 port map( A => n681, B => n623, C => n622, Y => n625);
   U863 : NAND2X1 port map( A => n691, B => n282, Y => n624);
   U864 : OAI21X1 port map( A => n703, B => n625, C => n624, Y => n626);
   U865 : NAND2X1 port map( A => n229, B => n626, Y => n628);
   U866 : NAND2X1 port map( A => n703, B => n245, Y => n627);
   U867 : AOI21X1 port map( A => n628, B => n627, C => n640, Y => n629);
   U868 : MUX2X1 port map( B => n629, A => n262, S => n656, Y => n631);
   U869 : NAND2X1 port map( A => n614, B => n255, Y => n630);
   U870 : NAND2X1 port map( A => n631, B => n630, Y => n633);
   U871 : MUX2X1 port map( B => n633, A => n246, S => n632, Y => n635);
   U872 : NAND2X1 port map( A => currentPlainKey_18_port, B => n268, Y => n634)
                           ;
   U873 : NAND3X1 port map( A => n636, B => n635, C => n634, Y => n1804);
   U874 : OAI22X1 port map( A => n250, B => n638, C => n276, D => n637, Y => 
                           n639);
   U875 : AOI21X1 port map( A => currentPlainKey_19_port, B => n266, C => n639,
                           Y => n655);
   U876 : OAI21X1 port map( A => n202, B => n211, C => currentPlainKey_19_port,
                           Y => n642);
   U877 : NAND2X1 port map( A => n713, B => n1357, Y => n641);
   U878 : NAND2X1 port map( A => n642, B => n641, Y => n644);
   U879 : NAND3X1 port map( A => n228, B => n644, C => n643, Y => n645);
   U880 : NAND2X1 port map( A => n183, B => n159, Y => n745);
   U881 : INVX2 port map( A => n745, Y => n726);
   U882 : MUX2X1 port map( B => n645, A => n233, S => n726, Y => n647);
   U883 : OAI22X1 port map( A => n240, B => n709, C => n238, D => n29, Y => 
                           n646);
   U884 : OAI21X1 port map( A => n647, B => n646, C => n688, Y => n651);
   U885 : AOI22X1 port map( A => n649, B => n260, C => n648, D => n253, Y => 
                           n650);
   U886 : NAND2X1 port map( A => n651, B => n650, Y => n652);
   U887 : NAND2X1 port map( A => n653, B => n652, Y => n654);
   U888 : NAND2X1 port map( A => n655, B => n654, Y => n1805);
   U889 : NAND2X1 port map( A => n656, B => n277, Y => n671);
   U890 : NAND2X1 port map( A => n183, B => n201, Y => n744);
   U891 : OAI21X1 port map( A => n71, B => n211, C => currentPlainKey_20_port, 
                           Y => n657);
   U892 : OAI21X1 port map( A => n1521, B => n211, C => n657, Y => n659);
   U893 : NOR2X1 port map( A => n272, B => n744, Y => n658);
   U894 : AOI21X1 port map( A => n97, B => n659, C => n658, Y => n661);
   U895 : NAND2X1 port map( A => n726, B => n281, Y => n660);
   U896 : OAI21X1 port map( A => n661, B => n739, C => n660, Y => n662);
   U897 : NAND2X1 port map( A => n229, B => n662, Y => n664);
   U898 : NAND2X1 port map( A => n739, B => n245, Y => n663);
   U899 : AOI21X1 port map( A => n664, B => n663, C => n675, Y => n665);
   U900 : NAND2X1 port map( A => n703, B => n255, Y => n666);
   U901 : NAND2X1 port map( A => n667, B => n666, Y => n668);
   U902 : MUX2X1 port map( B => n668, A => n246, S => n614, Y => n670);
   U903 : NAND2X1 port map( A => currentPlainKey_20_port, B => n269, Y => n669)
                           ;
   U904 : NAND3X1 port map( A => n671, B => n670, C => n669, Y => n1806);
   U905 : OAI22X1 port map( A => n250, B => n25, C => n275, D => n55, Y => n674
                           );
   U906 : AOI21X1 port map( A => currentPlainKey_21_port, B => n268, C => n674,
                           Y => n690);
   U907 : OAI21X1 port map( A => n206, B => n211, C => currentPlainKey_21_port,
                           Y => n677);
   U908 : INVX2 port map( A => n1544, Y => n1393);
   U909 : NAND2X1 port map( A => n713, B => n1393, Y => n676);
   U910 : NAND2X1 port map( A => n677, B => n676, Y => n679);
   U911 : NAND3X1 port map( A => n228, B => n679, C => n678, Y => n680);
   U912 : NAND2X1 port map( A => n183, B => n1520, Y => n780);
   U913 : INVX2 port map( A => n780, Y => n762);
   U914 : MUX2X1 port map( B => n680, A => n233, S => n762, Y => n683);
   U915 : OAI22X1 port map( A => n240, B => n745, C => n16, D => n744, Y => 
                           n682);
   U916 : OAI21X1 port map( A => n683, B => n682, C => n681, Y => n686);
   U917 : AOI22X1 port map( A => n684, B => n260, C => n691, D => n253, Y => 
                           n685);
   U918 : NAND2X1 port map( A => n686, B => n685, Y => n687);
   U919 : NAND2X1 port map( A => n688, B => n687, Y => n689);
   U920 : NAND2X1 port map( A => n690, B => n689, Y => n1807);
   U921 : NAND2X1 port map( A => n691, B => n280, Y => n707);
   U922 : NAND2X1 port map( A => n183, B => n205, Y => n779);
   U923 : NAND2X1 port map( A => n780, B => n779, Y => n782);
   U924 : OAI21X1 port map( A => n200, B => n211, C => currentPlainKey_22_port,
                           Y => n692);
   U925 : OAI21X1 port map( A => n1556, B => n211, C => n692, Y => n694);
   U926 : NOR2X1 port map( A => n272, B => n37, Y => n693);
   U927 : AOI21X1 port map( A => n753, B => n694, C => n693, Y => n696);
   U928 : NAND2X1 port map( A => n762, B => n281, Y => n695);
   U929 : OAI21X1 port map( A => n774, B => n696, C => n695, Y => n697);
   U930 : NAND2X1 port map( A => n229, B => n697, Y => n699);
   U931 : NAND2X1 port map( A => n774, B => n243, Y => n698);
   U932 : AOI21X1 port map( A => n699, B => n698, C => n711, Y => n700);
   U933 : MUX2X1 port map( B => n700, A => n262, S => n726, Y => n702);
   U934 : NAND2X1 port map( A => n739, B => n255, Y => n701);
   U935 : NAND2X1 port map( A => n702, B => n701, Y => n704);
   U936 : MUX2X1 port map( B => n704, A => n248, S => n703, Y => n706);
   U937 : NAND2X1 port map( A => currentPlainKey_22_port, B => n266, Y => n705)
                           ;
   U938 : NAND3X1 port map( A => n707, B => n706, C => n705, Y => n1808);
   U939 : OAI22X1 port map( A => n251, B => n709, C => n276, D => n29, Y => 
                           n710);
   U940 : AOI21X1 port map( A => currentPlainKey_23_port, B => n270, C => n710,
                           Y => n725);
   U941 : OAI21X1 port map( A => n204, B => n211, C => currentPlainKey_23_port,
                           Y => n715);
   U942 : NAND2X1 port map( A => n713, B => n1430, Y => n714);
   U943 : NAND2X1 port map( A => n715, B => n714, Y => n717);
   U944 : NAND3X1 port map( A => n228, B => n717, C => n716, Y => n718);
   U945 : NAND2X1 port map( A => n183, B => n186, Y => n815);
   U946 : INVX2 port map( A => n815, Y => n797);
   U947 : MUX2X1 port map( B => n718, A => n233, S => n797, Y => n720);
   U948 : OAI22X1 port map( A => n240, B => n780, C => n238, D => n37, Y => 
                           n719);
   U949 : OAI21X1 port map( A => n720, B => n719, C => n678, Y => n722);
   U950 : AOI22X1 port map( A => n774, B => n260, C => n726, D => n253, Y => 
                           n721);
   U951 : NAND2X1 port map( A => n722, B => n721, Y => n723);
   U952 : NAND2X1 port map( A => n643, B => n723, Y => n724);
   U953 : NAND2X1 port map( A => n725, B => n724, Y => n1809);
   U954 : NAND2X1 port map( A => n726, B => n278, Y => n743);
   U955 : NAND2X1 port map( A => n183, B => n191, Y => n814);
   U956 : NAND2X1 port map( A => n815, B => n814, Y => n817);
   U957 : INVX2 port map( A => n817, Y => n788);
   U958 : NAND3X1 port map( A => n222, B => address_4_port, C => n727, Y => 
                           n850);
   U959 : OAI21X1 port map( A => n1142, B => n213, C => currentPlainKey_24_port
                           , Y => n728);
   U960 : OAI21X1 port map( A => n1144, B => n213, C => n728, Y => n730);
   U961 : NOR2X1 port map( A => n272, B => n31, Y => n729);
   U962 : AOI21X1 port map( A => n788, B => n730, C => n729, Y => n732);
   U963 : NAND2X1 port map( A => n797, B => n281, Y => n731);
   U964 : OAI21X1 port map( A => n809, B => n732, C => n731, Y => n733);
   U965 : NAND2X1 port map( A => n229, B => n733, Y => n735);
   U966 : NAND2X1 port map( A => n809, B => n242, Y => n734);
   U967 : AOI21X1 port map( A => n735, B => n734, C => n747, Y => n736);
   U968 : MUX2X1 port map( B => n736, A => n261, S => n762, Y => n738);
   U969 : NAND2X1 port map( A => n774, B => n253, Y => n737);
   U970 : NAND2X1 port map( A => n738, B => n737, Y => n740);
   U971 : MUX2X1 port map( B => n740, A => n248, S => n739, Y => n742);
   U972 : NAND2X1 port map( A => currentPlainKey_24_port, B => n266, Y => n741)
                           ;
   U973 : NAND3X1 port map( A => n743, B => n742, C => n741, Y => n1810);
   U974 : OAI22X1 port map( A => n251, B => n745, C => n276, D => n744, Y => 
                           n746);
   U975 : AOI21X1 port map( A => currentPlainKey_25_port, B => n266, C => n746,
                           Y => n761);
   U976 : OAI21X1 port map( A => n196, B => n213, C => currentPlainKey_25_port,
                           Y => n749);
   U977 : INVX2 port map( A => n213, Y => n851);
   U978 : NAND2X1 port map( A => n851, B => n1470, Y => n748);
   U979 : NAND2X1 port map( A => n749, B => n748, Y => n751);
   U980 : NAND3X1 port map( A => n228, B => n751, C => n750, Y => n752);
   U981 : NAND2X1 port map( A => n158, B => n178, Y => n847);
   U982 : MUX2X1 port map( B => n752, A => n233, S => n824, Y => n755);
   U983 : OAI22X1 port map( A => n240, B => n815, C => n237, D => n31, Y => 
                           n754);
   U984 : OAI21X1 port map( A => n755, B => n754, C => n753, Y => n758);
   U985 : AOI22X1 port map( A => n756, B => n260, C => n762, D => n253, Y => 
                           n757);
   U986 : NAND2X1 port map( A => n758, B => n757, Y => n759);
   U987 : NAND2X1 port map( A => n678, B => n759, Y => n760);
   U988 : NAND2X1 port map( A => n761, B => n760, Y => n1811);
   U989 : NAND2X1 port map( A => n762, B => n279, Y => n778);
   U990 : NAND2X1 port map( A => n158, B => n1488, Y => n846);
   U991 : OAI21X1 port map( A => n75, B => n213, C => currentPlainKey_26_port, 
                           Y => n763);
   U992 : OAI21X1 port map( A => n1179, B => n213, C => n763, Y => n765);
   U993 : NOR2X1 port map( A => n272, B => n846, Y => n764);
   U994 : AOI21X1 port map( A => n137, B => n765, C => n764, Y => n767);
   U995 : NAND2X1 port map( A => n824, B => n281, Y => n766);
   U996 : OAI21X1 port map( A => n841, B => n767, C => n766, Y => n768);
   U997 : NAND2X1 port map( A => n229, B => n768, Y => n770);
   U998 : NAND2X1 port map( A => n841, B => n243, Y => n769);
   U999 : AOI21X1 port map( A => n770, B => n769, C => n782, Y => n771);
   U1000 : MUX2X1 port map( B => n771, A => n262, S => n797, Y => n773);
   U1001 : NAND2X1 port map( A => n809, B => n254, Y => n772);
   U1002 : NAND2X1 port map( A => n773, B => n772, Y => n775);
   U1003 : MUX2X1 port map( B => n775, A => n248, S => n774, Y => n777);
   U1004 : NAND2X1 port map( A => currentPlainKey_26_port, B => n268, Y => n776
                           );
   U1005 : NAND3X1 port map( A => n778, B => n777, C => n776, Y => n1812);
   U1006 : OAI22X1 port map( A => n251, B => n780, C => n276, D => n37, Y => 
                           n781);
   U1007 : AOI21X1 port map( A => currentPlainKey_27_port, B => n268, C => n781
                           , Y => n796);
   U1008 : OAI21X1 port map( A => n202, B => n213, C => currentPlainKey_27_port
                           , Y => n784);
   U1009 : NAND2X1 port map( A => n851, B => n1357, Y => n783);
   U1010 : NAND2X1 port map( A => n784, B => n783, Y => n786);
   U1011 : NAND3X1 port map( A => n228, B => n786, C => n785, Y => n787);
   U1012 : NAND2X1 port map( A => n158, B => n174, Y => n882);
   U1013 : INVX2 port map( A => n882, Y => n863);
   U1014 : MUX2X1 port map( B => n787, A => n233, S => n863, Y => n790);
   U1015 : OAI22X1 port map( A => n240, B => n847, C => n238, D => n846, Y => 
                           n789);
   U1016 : OAI21X1 port map( A => n790, B => n789, C => n788, Y => n793);
   U1017 : AOI22X1 port map( A => n791, B => n260, C => n797, D => n253, Y => 
                           n792);
   U1018 : NAND2X1 port map( A => n793, B => n792, Y => n794);
   U1019 : NAND2X1 port map( A => n716, B => n794, Y => n795);
   U1020 : NAND2X1 port map( A => n796, B => n795, Y => n1813);
   U1021 : NAND2X1 port map( A => n797, B => n277, Y => n813);
   U1022 : INVX2 port map( A => n846, Y => n876);
   U1023 : NAND2X1 port map( A => n158, B => n175, Y => n881);
   U1024 : OAI21X1 port map( A => n71, B => n213, C => currentPlainKey_28_port,
                           Y => n798);
   U1025 : OAI21X1 port map( A => n1521, B => n213, C => n798, Y => n800);
   U1026 : NOR2X1 port map( A => n272, B => n881, Y => n799);
   U1027 : AOI21X1 port map( A => n139, B => n800, C => n799, Y => n802);
   U1028 : NAND2X1 port map( A => n863, B => n281, Y => n801);
   U1029 : OAI21X1 port map( A => n802, B => n876, C => n801, Y => n803);
   U1030 : NAND2X1 port map( A => n229, B => n803, Y => n805);
   U1031 : NAND2X1 port map( A => n876, B => n243, Y => n804);
   U1032 : AOI21X1 port map( A => n805, B => n804, C => n817, Y => n806);
   U1033 : MUX2X1 port map( B => n806, A => n261, S => n824, Y => n808);
   U1034 : NAND2X1 port map( A => n841, B => n253, Y => n807);
   U1035 : NAND2X1 port map( A => n808, B => n807, Y => n810);
   U1036 : MUX2X1 port map( B => n810, A => n247, S => n809, Y => n812);
   U1037 : NAND2X1 port map( A => currentPlainKey_28_port, B => n266, Y => n811
                           );
   U1038 : NAND3X1 port map( A => n813, B => n812, C => n811, Y => n1814);
   U1039 : OAI22X1 port map( A => n251, B => n815, C => n276, D => n31, Y => 
                           n816);
   U1040 : AOI21X1 port map( A => currentPlainKey_29_port, B => n268, C => n816
                           , Y => n829);
   U1041 : OAI21X1 port map( A => n206, B => n213, C => currentPlainKey_29_port
                           , Y => n819);
   U1042 : NAND2X1 port map( A => n851, B => n1393, Y => n818);
   U1043 : NAND2X1 port map( A => n819, B => n818, Y => n820);
   U1044 : NAND3X1 port map( A => n227, B => n820, C => n896, Y => n821);
   U1045 : NAND2X1 port map( A => n158, B => n173, Y => n916);
   U1046 : MUX2X1 port map( B => n821, A => n234, S => n892, Y => n823);
   U1047 : OAI22X1 port map( A => n240, B => n882, C => n238, D => n11, Y => 
                           n822);
   U1048 : OAI21X1 port map( A => n823, B => n822, C => n785, Y => n826);
   U1049 : AOI22X1 port map( A => n876, B => n260, C => n824, D => n253, Y => 
                           n825);
   U1050 : NAND2X1 port map( A => n826, B => n825, Y => n827);
   U1051 : NAND2X1 port map( A => n750, B => n827, Y => n828);
   U1052 : NAND2X1 port map( A => n829, B => n828, Y => n1815);
   U1053 : NAND2X1 port map( A => n824, B => n279, Y => n845);
   U1054 : NAND2X1 port map( A => n158, B => n176, Y => n915);
   U1055 : OAI21X1 port map( A => n200, B => n213, C => currentPlainKey_30_port
                           , Y => n830);
   U1056 : OAI21X1 port map( A => n1556, B => n213, C => n830, Y => n832);
   U1057 : NOR2X1 port map( A => n272, B => n915, Y => n831);
   U1058 : AOI21X1 port map( A => n149, B => n832, C => n831, Y => n834);
   U1059 : NAND2X1 port map( A => n892, B => n281, Y => n833);
   U1060 : OAI21X1 port map( A => n834, B => n910, C => n833, Y => n835);
   U1061 : NAND2X1 port map( A => n229, B => n835, Y => n837);
   U1062 : NAND2X1 port map( A => n910, B => n244, Y => n836);
   U1063 : AOI21X1 port map( A => n837, B => n836, C => n849, Y => n838);
   U1064 : MUX2X1 port map( B => n838, A => n261, S => n863, Y => n840);
   U1065 : NAND2X1 port map( A => n876, B => n253, Y => n839);
   U1066 : NAND2X1 port map( A => n840, B => n839, Y => n842);
   U1067 : MUX2X1 port map( B => n842, A => n247, S => n841, Y => n844);
   U1068 : NAND2X1 port map( A => currentPlainKey_30_port, B => n268, Y => n843
                           );
   U1069 : NAND3X1 port map( A => n845, B => n844, C => n843, Y => n1816);
   U1070 : OAI22X1 port map( A => n251, B => n847, C => n275, D => n846, Y => 
                           n848);
   U1071 : AOI21X1 port map( A => currentPlainKey_31_port, B => n267, C => n848
                           , Y => n862);
   U1072 : OAI21X1 port map( A => n204, B => n213, C => currentPlainKey_31_port
                           , Y => n853);
   U1073 : NAND2X1 port map( A => n851, B => n1430, Y => n852);
   U1074 : NAND2X1 port map( A => n853, B => n852, Y => n854);
   U1075 : NAND3X1 port map( A => n228, B => n854, C => n931, Y => n855);
   U1076 : NAND2X1 port map( A => n158, B => n1130, Y => n952);
   U1077 : INVX2 port map( A => n952, Y => n934);
   U1078 : MUX2X1 port map( B => n855, A => n234, S => n934, Y => n857);
   U1079 : OAI22X1 port map( A => n240, B => n916, C => n237, D => n6, Y => 
                           n856);
   U1080 : OAI21X1 port map( A => n857, B => n856, C => n896, Y => n859);
   U1081 : AOI22X1 port map( A => n910, B => n259, C => n863, D => n252, Y => 
                           n858);
   U1082 : NAND2X1 port map( A => n859, B => n858, Y => n860);
   U1083 : NAND2X1 port map( A => n785, B => n860, Y => n861);
   U1084 : NAND2X1 port map( A => n862, B => n861, Y => n1817);
   U1085 : NAND2X1 port map( A => n863, B => n280, Y => n880);
   U1086 : INVX2 port map( A => n915, Y => n946);
   U1087 : NAND2X1 port map( A => n158, B => n179, Y => n951);
   U1088 : NAND3X1 port map( A => address_5_port, B => n221, C => n1004, Y => 
                           n989);
   U1089 : OAI21X1 port map( A => n1142, B => n215, C => 
                           currentPlainKey_32_port, Y => n865);
   U1090 : OAI21X1 port map( A => n1144, B => n215, C => n865, Y => n867);
   U1091 : NOR2X1 port map( A => n272, B => n951, Y => n866);
   U1092 : AOI21X1 port map( A => n153, B => n867, C => n866, Y => n869);
   U1093 : NAND2X1 port map( A => n934, B => n281, Y => n868);
   U1094 : OAI21X1 port map( A => n946, B => n869, C => n868, Y => n870);
   U1095 : NAND2X1 port map( A => n229, B => n870, Y => n872);
   U1096 : NAND2X1 port map( A => n946, B => n243, Y => n871);
   U1097 : AOI21X1 port map( A => n872, B => n871, C => n884, Y => n873);
   U1098 : MUX2X1 port map( B => n873, A => n261, S => n892, Y => n875);
   U1099 : NAND2X1 port map( A => n910, B => n253, Y => n874);
   U1100 : NAND2X1 port map( A => n875, B => n874, Y => n877);
   U1101 : MUX2X1 port map( B => n877, A => n247, S => n876, Y => n879);
   U1102 : NAND2X1 port map( A => currentPlainKey_32_port, B => n266, Y => n878
                           );
   U1103 : NAND3X1 port map( A => n880, B => n879, C => n878, Y => n1818);
   U1104 : OAI22X1 port map( A => n251, B => n93, C => n275, D => n11, Y => 
                           n883);
   U1105 : AOI21X1 port map( A => currentPlainKey_33_port, B => n267, C => n883
                           , Y => n898);
   U1106 : OAI21X1 port map( A => n196, B => n215, C => currentPlainKey_33_port
                           , Y => n886);
   U1107 : INVX2 port map( A => n215, Y => n990);
   U1108 : NAND2X1 port map( A => n990, B => n1470, Y => n885);
   U1109 : NAND2X1 port map( A => n886, B => n885, Y => n887);
   U1110 : NAND3X1 port map( A => n227, B => n887, C => n965, Y => n889);
   U1111 : NAND3X1 port map( A => n79, B => address_5_port, C => n1004, Y => 
                           n888);
   U1112 : NAND2X1 port map( A => n182, B => n47, Y => n986);
   U1113 : INVX2 port map( A => n986, Y => n968);
   U1114 : MUX2X1 port map( B => n889, A => n234, S => n968, Y => n891);
   U1115 : OAI22X1 port map( A => n239, B => n45, C => n16, D => n41, Y => n890
                           );
   U1116 : OAI21X1 port map( A => n891, B => n890, C => n931, Y => n894);
   U1117 : AOI22X1 port map( A => n946, B => n259, C => n892, D => n252, Y => 
                           n893);
   U1118 : NAND2X1 port map( A => n894, B => n893, Y => n895);
   U1119 : NAND2X1 port map( A => n896, B => n895, Y => n897);
   U1120 : NAND2X1 port map( A => n898, B => n897, Y => n1819);
   U1121 : NAND2X1 port map( A => n892, B => n279, Y => n914);
   U1122 : NAND2X1 port map( A => n182, B => n195, Y => n985);
   U1123 : NAND2X1 port map( A => n986, B => n985, Y => n988);
   U1124 : INVX2 port map( A => n988, Y => n959);
   U1125 : OAI21X1 port map( A => n75, B => n215, C => currentPlainKey_34_port,
                           Y => n899);
   U1126 : OAI21X1 port map( A => n1179, B => n215, C => n899, Y => n901);
   U1127 : NOR2X1 port map( A => n272, B => n33, Y => n900);
   U1128 : AOI21X1 port map( A => n959, B => n901, C => n900, Y => n903);
   U1129 : NAND2X1 port map( A => n968, B => n281, Y => n902);
   U1130 : OAI21X1 port map( A => n980, B => n903, C => n902, Y => n904);
   U1131 : NAND2X1 port map( A => n229, B => n904, Y => n906);
   U1132 : NAND2X1 port map( A => n980, B => n243, Y => n905);
   U1133 : AOI21X1 port map( A => n906, B => n905, C => n918, Y => n907);
   U1134 : MUX2X1 port map( B => n907, A => n261, S => n934, Y => n909);
   U1135 : NAND2X1 port map( A => n946, B => n254, Y => n908);
   U1136 : NAND2X1 port map( A => n909, B => n908, Y => n911);
   U1137 : MUX2X1 port map( B => n911, A => n247, S => n910, Y => n913);
   U1138 : NAND2X1 port map( A => currentPlainKey_34_port, B => n268, Y => n912
                           );
   U1139 : NAND3X1 port map( A => n914, B => n913, C => n912, Y => n1820);
   U1140 : OAI22X1 port map( A => n251, B => n916, C => n275, D => n6, Y => 
                           n917);
   U1141 : AOI21X1 port map( A => currentPlainKey_35_port, B => n269, C => n917
                           , Y => n933);
   U1142 : OAI21X1 port map( A => n202, B => n215, C => currentPlainKey_35_port
                           , Y => n920);
   U1143 : NAND2X1 port map( A => n990, B => n1357, Y => n919);
   U1144 : NAND2X1 port map( A => n920, B => n919, Y => n922);
   U1145 : NAND3X1 port map( A => n228, B => n922, C => n921, Y => n923);
   U1146 : NAND2X1 port map( A => n182, B => n159, Y => n1022);
   U1147 : INVX2 port map( A => n1022, Y => n1003);
   U1148 : MUX2X1 port map( B => n923, A => n234, S => n1003, Y => n925);
   U1149 : OAI22X1 port map( A => n239, B => n986, C => n237, D => n33, Y => 
                           n924);
   U1150 : OAI21X1 port map( A => n925, B => n924, C => n965, Y => n929);
   U1151 : AOI22X1 port map( A => n927, B => n259, C => n926, D => n252, Y => 
                           n928);
   U1152 : NAND2X1 port map( A => n929, B => n928, Y => n930);
   U1153 : NAND2X1 port map( A => n931, B => n930, Y => n932);
   U1154 : NAND2X1 port map( A => n933, B => n932, Y => n1821);
   U1155 : NAND2X1 port map( A => n934, B => n277, Y => n950);
   U1156 : NAND2X1 port map( A => n182, B => n201, Y => n1021);
   U1157 : OAI21X1 port map( A => n71, B => n215, C => currentPlainKey_36_port,
                           Y => n935);
   U1158 : OAI21X1 port map( A => n1521, B => n215, C => n935, Y => n937);
   U1159 : NOR2X1 port map( A => n272, B => n1021, Y => n936);
   U1160 : AOI21X1 port map( A => n99, B => n937, C => n936, Y => n939);
   U1161 : NAND2X1 port map( A => n1003, B => n281, Y => n938);
   U1162 : OAI21X1 port map( A => n1016, B => n939, C => n938, Y => n940);
   U1163 : NAND2X1 port map( A => n229, B => n940, Y => n942);
   U1164 : NAND2X1 port map( A => n1016, B => n243, Y => n941);
   U1165 : AOI21X1 port map( A => n942, B => n941, C => n954, Y => n943);
   U1166 : NAND2X1 port map( A => n980, B => n254, Y => n944);
   U1167 : NAND2X1 port map( A => n944, B => n945, Y => n947);
   U1168 : MUX2X1 port map( B => n947, A => n247, S => n946, Y => n949);
   U1169 : NAND2X1 port map( A => currentPlainKey_36_port, B => n270, Y => n948
                           );
   U1170 : NAND3X1 port map( A => n950, B => n949, C => n948, Y => n1822);
   U1171 : OAI22X1 port map( A => n251, B => n45, C => n275, D => n41, Y => 
                           n953);
   U1172 : AOI21X1 port map( A => currentPlainKey_37_port, B => n270, C => n953
                           , Y => n967);
   U1173 : OAI21X1 port map( A => n206, B => n215, C => currentPlainKey_37_port
                           , Y => n956);
   U1174 : NAND2X1 port map( A => n990, B => n1393, Y => n955);
   U1175 : NAND2X1 port map( A => n956, B => n955, Y => n957);
   U1176 : NAND3X1 port map( A => n227, B => n957, C => n1036, Y => n958);
   U1177 : NAND2X1 port map( A => n182, B => n1520, Y => n1057);
   U1178 : INVX2 port map( A => n1057, Y => n1039);
   U1179 : MUX2X1 port map( B => n958, A => n234, S => n1039, Y => n961);
   U1180 : OAI22X1 port map( A => n239, B => n1022, C => n237, D => n1021, Y =>
                           n960);
   U1181 : OAI21X1 port map( A => n961, B => n960, C => n959, Y => n963);
   U1182 : AOI22X1 port map( A => n1016, B => n259, C => n968, D => n252, Y => 
                           n962);
   U1183 : NAND2X1 port map( A => n963, B => n962, Y => n964);
   U1184 : NAND2X1 port map( A => n965, B => n964, Y => n966);
   U1185 : NAND2X1 port map( A => n967, B => n966, Y => n1823);
   U1186 : NAND2X1 port map( A => n968, B => n280, Y => n984);
   U1187 : NAND2X1 port map( A => n182, B => n205, Y => n1056);
   U1188 : NAND2X1 port map( A => n1057, B => n1056, Y => n1059);
   U1189 : INVX2 port map( A => n1059, Y => n1029);
   U1190 : OAI21X1 port map( A => n199, B => n215, C => currentPlainKey_38_port
                           , Y => n969);
   U1191 : OAI21X1 port map( A => n1556, B => n215, C => n969, Y => n971);
   U1192 : NOR2X1 port map( A => n272, B => n39, Y => n970);
   U1193 : AOI21X1 port map( A => n1029, B => n971, C => n970, Y => n973);
   U1194 : NAND2X1 port map( A => n1039, B => n281, Y => n972);
   U1195 : OAI21X1 port map( A => n1051, B => n973, C => n972, Y => n974);
   U1196 : NAND2X1 port map( A => n229, B => n974, Y => n976);
   U1197 : NAND2X1 port map( A => n1051, B => n244, Y => n975);
   U1198 : AOI21X1 port map( A => n976, B => n975, C => n988, Y => n977);
   U1199 : MUX2X1 port map( B => n977, A => n261, S => n1003, Y => n979);
   U1200 : NAND2X1 port map( A => n1016, B => n254, Y => n978);
   U1201 : NAND2X1 port map( A => n979, B => n978, Y => n981);
   U1202 : MUX2X1 port map( B => n981, A => n247, S => n980, Y => n983);
   U1203 : NAND2X1 port map( A => currentPlainKey_38_port, B => n268, Y => n982
                           );
   U1204 : NAND3X1 port map( A => n984, B => n983, C => n982, Y => n1824);
   U1205 : OAI22X1 port map( A => n250, B => n986, C => n275, D => n33, Y => 
                           n987);
   U1206 : AOI21X1 port map( A => currentPlainKey_39_port, B => n269, C => n987
                           , Y => n1002);
   U1207 : OAI21X1 port map( A => n204, B => n215, C => currentPlainKey_39_port
                           , Y => n992);
   U1208 : NAND2X1 port map( A => n990, B => n1430, Y => n991);
   U1209 : NAND2X1 port map( A => n992, B => n991, Y => n994);
   U1210 : NAND3X1 port map( A => n227, B => n994, C => n993, Y => n995);
   U1211 : NAND2X1 port map( A => n182, B => n186, Y => n1090);
   U1212 : INVX2 port map( A => n1090, Y => n1072);
   U1213 : MUX2X1 port map( B => n995, A => n234, S => n1072, Y => n997);
   U1214 : OAI22X1 port map( A => n239, B => n1057, C => n238, D => n39, Y => 
                           n996);
   U1215 : OAI21X1 port map( A => n997, B => n996, C => n1036, Y => n999);
   U1216 : AOI22X1 port map( A => n1051, B => n259, C => n1003, D => n252, Y =>
                           n998);
   U1217 : NAND2X1 port map( A => n999, B => n998, Y => n1000);
   U1218 : NAND2X1 port map( A => n921, B => n1000, Y => n1001);
   U1219 : NAND2X1 port map( A => n1002, B => n1001, Y => n1825);
   U1220 : NAND2X1 port map( A => n1003, B => n277, Y => n1020);
   U1221 : NAND2X1 port map( A => n182, B => n191, Y => n1089);
   U1222 : NAND3X1 port map( A => n222, B => address_5_port, C => n1004, Y => 
                           n1125);
   U1223 : OAI21X1 port map( A => n1142, B => n217, C => 
                           currentPlainKey_40_port, Y => n1005);
   U1224 : OAI21X1 port map( A => n1144, B => n217, C => n1005, Y => n1007);
   U1225 : NOR2X1 port map( A => n272, B => n1089, Y => n1006);
   U1226 : AOI21X1 port map( A => n95, B => n1007, C => n1006, Y => n1009);
   U1227 : NAND2X1 port map( A => n1072, B => n281, Y => n1008);
   U1228 : OAI21X1 port map( A => n1084, B => n1009, C => n1008, Y => n1010);
   U1229 : NAND2X1 port map( A => n229, B => n1010, Y => n1012);
   U1230 : NAND2X1 port map( A => n1084, B => n244, Y => n1011);
   U1231 : AOI21X1 port map( A => n1012, B => n1011, C => n1024, Y => n1013);
   U1232 : NAND2X1 port map( A => n1051, B => n254, Y => n1014);
   U1233 : NAND2X1 port map( A => n1014, B => n1015, Y => n1017);
   U1234 : MUX2X1 port map( B => n1017, A => n247, S => n1016, Y => n1019);
   U1235 : NAND2X1 port map( A => currentPlainKey_40_port, B => n266, Y => 
                           n1018);
   U1236 : NAND3X1 port map( A => n1020, B => n1019, C => n1018, Y => n1826);
   U1237 : OAI22X1 port map( A => n250, B => n1022, C => n275, D => n1021, Y =>
                           n1023);
   U1238 : AOI21X1 port map( A => currentPlainKey_41_port, B => n266, C => 
                           n1023, Y => n1038);
   U1239 : OAI21X1 port map( A => n196, B => n217, C => currentPlainKey_41_port
                           , Y => n1026);
   U1240 : INVX2 port map( A => n217, Y => n1126);
   U1241 : NAND2X1 port map( A => n1126, B => n1470, Y => n1025);
   U1242 : NAND2X1 port map( A => n1026, B => n1025, Y => n1027);
   U1243 : NAND3X1 port map( A => n227, B => n1027, C => n1102, Y => n1028);
   U1244 : NAND2X1 port map( A => n1141, B => n178, Y => n1122);
   U1245 : MUX2X1 port map( B => n1028, A => n234, S => n1105, Y => n1031);
   U1246 : OAI22X1 port map( A => n239, B => n1090, C => n16, D => n1089, Y => 
                           n1030);
   U1247 : OAI21X1 port map( A => n1031, B => n1030, C => n1029, Y => n1034);
   U1248 : AOI22X1 port map( A => n1032, B => n259, C => n1039, D => n252, Y =>
                           n1033);
   U1249 : NAND2X1 port map( A => n1034, B => n1033, Y => n1035);
   U1250 : NAND2X1 port map( A => n1036, B => n1035, Y => n1037);
   U1251 : NAND2X1 port map( A => n1038, B => n1037, Y => n1827);
   U1252 : NAND2X1 port map( A => n1039, B => n278, Y => n1055);
   U1253 : NAND2X1 port map( A => n1141, B => n1488, Y => n1121);
   U1254 : OAI21X1 port map( A => n75, B => n217, C => currentPlainKey_42_port,
                           Y => n1040);
   U1255 : OAI21X1 port map( A => n1179, B => n217, C => n1040, Y => n1042);
   U1256 : NOR2X1 port map( A => n272, B => n1121, Y => n1041);
   U1257 : AOI21X1 port map( A => n127, B => n1042, C => n1041, Y => n1044);
   U1258 : NAND2X1 port map( A => n1105, B => n281, Y => n1043);
   U1259 : OAI21X1 port map( A => n1066, B => n1044, C => n1043, Y => n1045);
   U1260 : NAND2X1 port map( A => n229, B => n1045, Y => n1047);
   U1261 : NAND2X1 port map( A => n1066, B => n244, Y => n1046);
   U1262 : AOI21X1 port map( A => n1047, B => n1046, C => n1059, Y => n1048);
   U1263 : MUX2X1 port map( B => n1048, A => n261, S => n1072, Y => n1050);
   U1264 : NAND2X1 port map( A => n1084, B => n254, Y => n1049);
   U1265 : NAND2X1 port map( A => n1050, B => n1049, Y => n1052);
   U1266 : NAND2X1 port map( A => currentPlainKey_42_port, B => n268, Y => 
                           n1053);
   U1267 : NAND3X1 port map( A => n1055, B => n1053, C => n1054, Y => n1828);
   U1268 : OAI22X1 port map( A => n250, B => n1057, C => n275, D => n39, Y => 
                           n1058);
   U1269 : AOI21X1 port map( A => currentPlainKey_43_port, B => n268, C => 
                           n1058, Y => n1071);
   U1270 : OAI21X1 port map( A => n202, B => n217, C => currentPlainKey_43_port
                           , Y => n1061);
   U1271 : NAND2X1 port map( A => n1126, B => n1357, Y => n1060);
   U1272 : NAND2X1 port map( A => n1061, B => n1060, Y => n1062);
   U1273 : NAND3X1 port map( A => n227, B => n1062, C => n1137, Y => n1063);
   U1274 : NAND2X1 port map( A => n1141, B => n174, Y => n1161);
   U1275 : INVX2 port map( A => n1161, Y => n1140);
   U1276 : MUX2X1 port map( B => n1063, A => n234, S => n1140, Y => n1065);
   U1277 : OAI22X1 port map( A => n239, B => n1122, C => n16, D => n9, Y => 
                           n1064);
   U1278 : OAI21X1 port map( A => n1065, B => n1064, C => n1102, Y => n1068);
   U1279 : INVX2 port map( A => n1089, Y => n1066);
   U1280 : AOI22X1 port map( A => n1066, B => n259, C => n1072, D => n252, Y =>
                           n1067);
   U1281 : NAND2X1 port map( A => n1068, B => n1067, Y => n1069);
   U1282 : NAND2X1 port map( A => n993, B => n1069, Y => n1070);
   U1283 : NAND2X1 port map( A => n1071, B => n1070, Y => n1829);
   U1284 : NAND2X1 port map( A => n1072, B => n280, Y => n1088);
   U1285 : NAND2X1 port map( A => n1141, B => n175, Y => n1160);
   U1286 : OAI21X1 port map( A => n71, B => n217, C => currentPlainKey_44_port,
                           Y => n1073);
   U1287 : OAI21X1 port map( A => n1521, B => n217, C => n1073, Y => n1075);
   U1288 : NOR2X1 port map( A => n271, B => n1160, Y => n1074);
   U1289 : AOI21X1 port map( A => n135, B => n1075, C => n1074, Y => n1077);
   U1290 : NAND2X1 port map( A => n1140, B => n281, Y => n1076);
   U1291 : OAI21X1 port map( A => n1077, B => n1155, C => n1076, Y => n1078);
   U1292 : NAND2X1 port map( A => n229, B => n1078, Y => n1080);
   U1293 : NAND2X1 port map( A => n1155, B => n244, Y => n1079);
   U1294 : AOI21X1 port map( A => n1080, B => n1079, C => n1092, Y => n1081);
   U1295 : MUX2X1 port map( B => n1081, A => n261, S => n1105, Y => n1083);
   U1296 : NAND2X1 port map( A => n1066, B => n254, Y => n1082);
   U1297 : NAND2X1 port map( A => n1083, B => n1082, Y => n1085);
   U1298 : MUX2X1 port map( B => n1085, A => n247, S => n1084, Y => n1087);
   U1299 : NAND2X1 port map( A => currentPlainKey_44_port, B => n266, Y => 
                           n1086);
   U1300 : NAND3X1 port map( A => n1088, B => n1087, C => n1086, Y => n1830);
   U1301 : OAI22X1 port map( A => n251, B => n1090, C => n275, D => n1089, Y =>
                           n1091);
   U1302 : AOI21X1 port map( A => currentPlainKey_45_port, B => n266, C => 
                           n1091, Y => n1104);
   U1303 : OAI21X1 port map( A => n206, B => n217, C => currentPlainKey_45_port
                           , Y => n1094);
   U1304 : NAND2X1 port map( A => n1126, B => n1393, Y => n1093);
   U1306 : NAND2X1 port map( A => n1094, B => n1093, Y => n1095);
   U1307 : NAND3X1 port map( A => n227, B => n1095, C => n135, Y => n1096);
   U1308 : NAND2X1 port map( A => n1141, B => n173, Y => n1196);
   U1309 : INVX2 port map( A => n1196, Y => n1175);
   U1310 : MUX2X1 port map( B => n1096, A => n234, S => n1175, Y => n1098);
   U1311 : OAI22X1 port map( A => n239, B => n1161, C => n16, D => n10, Y => 
                           n1097);
   U1312 : OAI21X1 port map( A => n1098, B => n1097, C => n1137, Y => n1100);
   U1313 : AOI22X1 port map( A => n1155, B => n259, C => n1105, D => n252, Y =>
                           n1099);
   U1314 : NAND2X1 port map( A => n1100, B => n1099, Y => n1101);
   U1315 : NAND2X1 port map( A => n1102, B => n1101, Y => n1103);
   U1316 : NAND2X1 port map( A => n1104, B => n1103, Y => n1831);
   U1317 : NAND2X1 port map( A => n1105, B => n280, Y => n1120);
   U1318 : NAND2X1 port map( A => n1141, B => n176, Y => n1195);
   U1319 : OAI21X1 port map( A => n199, B => n217, C => currentPlainKey_46_port
                           , Y => n1106);
   U1320 : OAI21X1 port map( A => n1556, B => n217, C => n1106, Y => n1108);
   U1321 : NOR2X1 port map( A => n271, B => n1195, Y => n1107);
   U1322 : AOI21X1 port map( A => n154, B => n1108, C => n1107, Y => n1110);
   U1323 : NAND2X1 port map( A => n1175, B => n281, Y => n1109);
   U1324 : OAI21X1 port map( A => n1110, B => n1190, C => n1109, Y => n1111);
   U1325 : NAND2X1 port map( A => n229, B => n1111, Y => n1113);
   U1326 : NAND2X1 port map( A => n1190, B => n245, Y => n1112);
   U1327 : AOI21X1 port map( A => n1113, B => n1112, C => n1124, Y => n1114);
   U1328 : MUX2X1 port map( B => n1114, A => n261, S => n1140, Y => n1116);
   U1329 : NAND2X1 port map( A => n1155, B => n254, Y => n1115);
   U1330 : NAND2X1 port map( A => n1116, B => n1115, Y => n1117);
   U1331 : MUX2X1 port map( B => n1117, A => n246, S => n1066, Y => n1119);
   U1332 : NAND2X1 port map( A => currentPlainKey_46_port, B => n268, Y => 
                           n1118);
   U1333 : NAND3X1 port map( A => n1120, B => n1119, C => n1118, Y => n1832);
   U1334 : OAI22X1 port map( A => n249, B => n1122, C => n276, D => n9, Y => 
                           n1123);
   U1335 : AOI21X1 port map( A => currentPlainKey_47_port, B => n268, C => 
                           n1123, Y => n1139);
   U1336 : OAI21X1 port map( A => n204, B => n217, C => currentPlainKey_47_port
                           , Y => n1128);
   U1337 : NAND2X1 port map( A => n1126, B => n1430, Y => n1127);
   U1338 : NAND2X1 port map( A => n1128, B => n1127, Y => n1129);
   U1339 : NAND3X1 port map( A => n227, B => n1129, C => n1368, Y => n1131);
   U1340 : NAND2X1 port map( A => n1141, B => n1130, Y => n1390);
   U1341 : INVX2 port map( A => n1390, Y => n1371);
   U1342 : MUX2X1 port map( B => n1131, A => n234, S => n1371, Y => n1133);
   U1343 : OAI22X1 port map( A => n239, B => n89, C => n237, D => n59, Y => 
                           n1132);
   U1344 : OAI21X1 port map( A => n1133, B => n1132, C => n135, Y => n1135);
   U1345 : AOI22X1 port map( A => n1190, B => n259, C => n1140, D => n252, Y =>
                           n1134);
   U1346 : NAND2X1 port map( A => n1135, B => n1134, Y => n1136);
   U1347 : NAND2X1 port map( A => n1137, B => n1136, Y => n1138);
   U1348 : NAND2X1 port map( A => n1139, B => n1138, Y => n1833);
   U1349 : NAND2X1 port map( A => n1140, B => n279, Y => n1159);
   U1350 : NAND2X1 port map( A => n1141, B => n179, Y => n1389);
   U1351 : OAI21X1 port map( A => n1142, B => n218, C => 
                           currentPlainKey_48_port, Y => n1143);
   U1358 : OAI21X1 port map( A => n1144, B => n218, C => n1143, Y => n1146);
   U1359 : NOR2X1 port map( A => n271, B => n1389, Y => n1145);
   U1360 : AOI21X1 port map( A => n145, B => n1146, C => n1145, Y => n1148);
   U1361 : NAND2X1 port map( A => n1371, B => n281, Y => n1147);
   U1362 : OAI21X1 port map( A => n1384, B => n1148, C => n1147, Y => n1149);
   U1363 : NAND2X1 port map( A => n229, B => n1149, Y => n1151);
   U1364 : NAND2X1 port map( A => n1384, B => n245, Y => n1150);
   U1365 : AOI21X1 port map( A => n1151, B => n1150, C => n1163, Y => n1152);
   U1366 : MUX2X1 port map( B => n1152, A => n261, S => n1175, Y => n1154);
   U1367 : NAND2X1 port map( A => n1190, B => n254, Y => n1153);
   U1368 : NAND2X1 port map( A => n1154, B => n1153, Y => n1156);
   U1369 : MUX2X1 port map( B => n1156, A => n248, S => n1155, Y => n1158);
   U1370 : NAND2X1 port map( A => currentPlainKey_48_port, B => n268, Y => 
                           n1157);
   U1371 : NAND3X1 port map( A => n1159, B => n1158, C => n1157, Y => n1834);
   U1372 : OAI22X1 port map( A => n251, B => n1161, C => n275, D => n10, Y => 
                           n1162);
   U1373 : AOI21X1 port map( A => currentPlainKey_49_port, B => n270, C => 
                           n1162, Y => n1174);
   U1374 : OAI21X1 port map( A => n196, B => n218, C => currentPlainKey_49_port
                           , Y => n1165);
   U1375 : INVX2 port map( A => n218, Y => n1429);
   U1376 : NAND2X1 port map( A => n1429, B => n1470, Y => n1164);
   U1377 : NAND2X1 port map( A => n1165, B => n1164, Y => n1166);
   U1378 : NAND3X1 port map( A => n227, B => n1166, C => n1404, Y => n1167);
   U1379 : NAND2X1 port map( A => n79, B => n188, Y => n1582);
   U1380 : NAND2X1 port map( A => n169, B => n47, Y => n1425);
   U1381 : INVX2 port map( A => n1425, Y => n1407);
   U1382 : MUX2X1 port map( B => n1167, A => n234, S => n1407, Y => n1169);
   U1383 : OAI22X1 port map( A => n239, B => n20, C => n16, D => n51, Y => 
                           n1168);
   U1384 : OAI21X1 port map( A => n1169, B => n1168, C => n1368, Y => n1171);
   U1385 : AOI22X1 port map( A => n1384, B => n259, C => n1175, D => n252, Y =>
                           n1170);
   U1386 : NAND2X1 port map( A => n1171, B => n1170, Y => n1172);
   U1387 : NAND2X1 port map( A => n135, B => n1172, Y => n1173);
   U1388 : NAND2X1 port map( A => n1174, B => n1173, Y => n1835);
   U1389 : NAND2X1 port map( A => n1175, B => n278, Y => n1194);
   U1390 : NAND2X1 port map( A => n169, B => n195, Y => n1424);
   U1391 : OAI21X1 port map( A => n75, B => n218, C => currentPlainKey_50_port,
                           Y => n1177);
   U1392 : OAI21X1 port map( A => n1179, B => n218, C => n1177, Y => n1181);
   U1393 : NOR2X1 port map( A => n271, B => n1424, Y => n1180);
   U1394 : AOI21X1 port map( A => n129, B => n1181, C => n1180, Y => n1183);
   U1395 : NAND2X1 port map( A => n1407, B => n281, Y => n1182);
   U1396 : OAI21X1 port map( A => n1419, B => n1183, C => n1182, Y => n1184);
   U1397 : NAND2X1 port map( A => n229, B => n1184, Y => n1186);
   U1398 : NAND2X1 port map( A => n1419, B => n242, Y => n1185);
   U1399 : AOI21X1 port map( A => n1186, B => n1185, C => n1268, Y => n1187);
   U1400 : MUX2X1 port map( B => n1187, A => n260, S => n1371, Y => n1189);
   U1401 : NAND2X1 port map( A => n1384, B => n254, Y => n1188);
   U1402 : NAND2X1 port map( A => n1189, B => n1188, Y => n1191);
   U1403 : MUX2X1 port map( B => n1191, A => n248, S => n1190, Y => n1193);
   U1404 : NAND2X1 port map( A => currentPlainKey_50_port, B => n270, Y => 
                           n1192);
   U1405 : NAND3X1 port map( A => n1194, B => n1193, C => n1192, Y => n1836);
   U1406 : OAI22X1 port map( A => n251, B => n89, C => n275, D => n59, Y => 
                           n1267);
   U1407 : AOI21X1 port map( A => currentPlainKey_51_port, B => n269, C => 
                           n1267, Y => n1370);
   U1408 : OAI21X1 port map( A => n202, B => n218, C => currentPlainKey_51_port
                           , Y => n1359);
   U1409 : NAND2X1 port map( A => n1357, B => n1429, Y => n1358);
   U1410 : NAND2X1 port map( A => n1359, B => n1358, Y => n1360);
   U1411 : NAND3X1 port map( A => n227, B => n1360, C => n1441, Y => n1361);
   U1412 : NAND2X1 port map( A => n169, B => n159, Y => n1481);
   U1413 : MUX2X1 port map( B => n1361, A => n234, S => n1444, Y => n1363);
   U1414 : OAI22X1 port map( A => n239, B => n43, C => n237, D => n21, Y => 
                           n1362);
   U1415 : OAI21X1 port map( A => n1363, B => n1362, C => n1404, Y => n1366);
   U1416 : AOI22X1 port map( A => n1419, B => n259, C => n1364, D => n252, Y =>
                           n1365);
   U1417 : NAND2X1 port map( A => n1366, B => n1365, Y => n1367);
   U1418 : NAND2X1 port map( A => n1368, B => n1367, Y => n1369);
   U1419 : NAND2X1 port map( A => n1370, B => n1369, Y => n1837);
   U1420 : NAND2X1 port map( A => n1371, B => n278, Y => n1388);
   U1421 : NAND2X1 port map( A => n169, B => n201, Y => n1480);
   U1422 : OAI21X1 port map( A => n71, B => n218, C => currentPlainKey_52_port,
                           Y => n1373);
   U1423 : OAI21X1 port map( A => n1521, B => n218, C => n1373, Y => n1375);
   U1424 : NOR2X1 port map( A => n271, B => n1480, Y => n1374);
   U1425 : AOI21X1 port map( A => n147, B => n1375, C => n1374, Y => n1377);
   U1426 : NAND2X1 port map( A => n1444, B => n281, Y => n1376);
   U1427 : OAI21X1 port map( A => n1460, B => n1377, C => n1376, Y => n1378);
   U1428 : NAND2X1 port map( A => n229, B => n1378, Y => n1380);
   U1429 : NAND2X1 port map( A => n1460, B => n242, Y => n1379);
   U1430 : AOI21X1 port map( A => n1380, B => n1379, C => n1392, Y => n1381);
   U1431 : MUX2X1 port map( B => n1381, A => n260, S => n1407, Y => n1383);
   U1432 : NAND2X1 port map( A => n1419, B => n254, Y => n1382);
   U1433 : NAND2X1 port map( A => n1383, B => n1382, Y => n1385);
   U1434 : MUX2X1 port map( B => n1385, A => n248, S => n1384, Y => n1387);
   U1435 : NAND2X1 port map( A => currentPlainKey_52_port, B => n269, Y => 
                           n1386);
   U1436 : NAND3X1 port map( A => n1388, B => n1387, C => n1386, Y => n1838);
   U1437 : OAI22X1 port map( A => n251, B => n20, C => n275, D => n51, Y => 
                           n1391);
   U1438 : AOI21X1 port map( A => currentPlainKey_53_port, B => n267, C => 
                           n1391, Y => n1406);
   U1439 : OAI21X1 port map( A => n206, B => n218, C => currentPlainKey_53_port
                           , Y => n1395);
   U1440 : NAND2X1 port map( A => n1429, B => n1393, Y => n1394);
   U1441 : NAND2X1 port map( A => n1395, B => n1394, Y => n1396);
   U1442 : NAND3X1 port map( A => n227, B => n1396, C => n147, Y => n1397);
   U1443 : NAND2X1 port map( A => n169, B => n1520, Y => n1465);
   U1444 : INVX2 port map( A => n1465, Y => n1515);
   U1445 : MUX2X1 port map( B => n1397, A => n235, S => n1515, Y => n1399);
   U1446 : OAI22X1 port map( A => n239, B => n27, C => n238, D => n65, Y => 
                           n1398);
   U1447 : OAI21X1 port map( A => n1399, B => n1398, C => n1441, Y => n1402);
   U1448 : AOI22X1 port map( A => n1400, B => n259, C => n1407, D => n252, Y =>
                           n1401);
   U1449 : NAND2X1 port map( A => n1402, B => n1401, Y => n1403);
   U1450 : NAND2X1 port map( A => n1404, B => n1403, Y => n1405);
   U1451 : NAND2X1 port map( A => n1406, B => n1405, Y => n1839);
   U1452 : NAND2X1 port map( A => n1407, B => n278, Y => n1423);
   U1453 : NAND2X1 port map( A => n169, B => n205, Y => n1453);
   U1454 : OAI21X1 port map( A => n199, B => n218, C => currentPlainKey_54_port
                           , Y => n1408);
   U1455 : OAI21X1 port map( A => n218, B => n1556, C => n1408, Y => n1410);
   U1456 : NOR2X1 port map( A => n271, B => n1453, Y => n1409);
   U1457 : AOI21X1 port map( A => n119, B => n1410, C => n1409, Y => n1412);
   U1458 : NAND2X1 port map( A => n1515, B => n281, Y => n1411);
   U1459 : OAI21X1 port map( A => n1437, B => n1412, C => n1411, Y => n1413);
   U1460 : NAND2X1 port map( A => n229, B => n1413, Y => n1415);
   U1461 : NAND2X1 port map( A => n1437, B => n242, Y => n1414);
   U1462 : AOI21X1 port map( A => n1415, B => n1414, C => n1427, Y => n1416);
   U1463 : MUX2X1 port map( B => n1416, A => n260, S => n1444, Y => n1418);
   U1464 : NAND2X1 port map( A => n1460, B => n254, Y => n1417);
   U1465 : NAND2X1 port map( A => n1418, B => n1417, Y => n1420);
   U1466 : MUX2X1 port map( B => n1420, A => n248, S => n1419, Y => n1422);
   U1467 : NAND2X1 port map( A => currentPlainKey_54_port, B => n268, Y => 
                           n1421);
   U1468 : NAND3X1 port map( A => n1423, B => n1422, C => n1421, Y => n1840);
   U1469 : OAI22X1 port map( A => n251, B => n43, C => n275, D => n21, Y => 
                           n1426);
   U1470 : AOI21X1 port map( A => currentPlainKey_55_port, B => n268, C => 
                           n1426, Y => n1443);
   U1471 : OAI21X1 port map( A => n204, B => n218, C => currentPlainKey_55_port
                           , Y => n1432);
   U1472 : NAND2X1 port map( A => n1430, B => n1429, Y => n1431);
   U1473 : NAND2X1 port map( A => n1432, B => n1431, Y => n1433);
   U1474 : NAND3X1 port map( A => n227, B => n1433, C => n119, Y => n1434);
   U1475 : NAND2X1 port map( A => n169, B => n186, Y => n1504);
   U1476 : INVX2 port map( A => n1504, Y => n1552);
   U1477 : MUX2X1 port map( B => n1434, A => n235, S => n1552, Y => n1436);
   U1478 : OAI22X1 port map( A => n5, B => n239, C => n1453, D => n237, Y => 
                           n1435);
   U1479 : OAI21X1 port map( A => n1436, B => n1435, C => n147, Y => n1439);
   U1480 : AOI22X1 port map( A => n1437, B => n259, C => n1444, D => n252, Y =>
                           n1438);
   U1481 : NAND2X1 port map( A => n1439, B => n1438, Y => n1440);
   U1482 : NAND2X1 port map( A => n1441, B => n1440, Y => n1442);
   U1483 : NAND2X1 port map( A => n1443, B => n1442, Y => n1841);
   U1484 : NAND2X1 port map( A => n1444, B => n280, Y => n1464);
   U1485 : NAND2X1 port map( A => n1552, B => n281, Y => n1451);
   U1486 : NAND2X1 port map( A => n223, B => n188, Y => n1578);
   U1487 : NAND2X1 port map( A => n1557, B => n47, Y => n1446);
   U1488 : AOI22X1 port map( A => currentPlainKey_56_port, B => n1446, C => 
                           n1445, D => n1557, Y => n1448);
   U1489 : NAND2X1 port map( A => n169, B => n191, Y => n1503);
   U1490 : NAND2X1 port map( A => n1504, B => n1503, Y => n1467);
   U1491 : NAND2X1 port map( A => n1571, B => RCV_DATA(1), Y => n1447);
   U1492 : OAI21X1 port map( A => n1448, B => n1467, C => n1447, Y => n1449);
   U1493 : NAND2X1 port map( A => n1449, B => n1453, Y => n1450);
   U1494 : NAND2X1 port map( A => n1451, B => n1450, Y => n1452);
   U1495 : NAND2X1 port map( A => n229, B => n1452, Y => n1456);
   U1496 : NAND2X1 port map( A => n244, B => n1534, Y => n1455);
   U1497 : AOI21X1 port map( A => n1456, B => n1455, C => n1454, Y => n1457);
   U1498 : MUX2X1 port map( B => n1457, A => n260, S => n1515, Y => n1459);
   U1499 : NAND2X1 port map( A => n1437, B => n254, Y => n1458);
   U1500 : NAND2X1 port map( A => n1459, B => n1458, Y => n1461);
   U1501 : MUX2X1 port map( B => n1461, A => n248, S => n1460, Y => n1463);
   U1502 : NAND2X1 port map( A => currentPlainKey_56_port, B => n267, Y => 
                           n1462);
   U1503 : NOR2X1 port map( A => n257, B => n5, Y => n1479);
   U1504 : OAI22X1 port map( A => n7, B => n167, C => n63, D => n236, Y => 
                           n1475);
   U1505 : NAND2X1 port map( A => n1561, B => n178, Y => n1529);
   U1506 : INVX2 port map( A => n1467, Y => n1468);
   U1507 : NOR2X1 port map( A => n111, B => n113, Y => n1474);
   U1508 : OAI21X1 port map( A => n196, B => n61, C => currentPlainKey_57_port,
                           Y => n1472);
   U1509 : NAND2X1 port map( A => n1470, B => n1557, Y => n1471);
   U1510 : NAND2X1 port map( A => n168, B => n1529, Y => n1519);
   U1511 : AOI21X1 port map( A => n1472, B => n1471, C => n1519, Y => n1473);
   U1512 : NOR3X1 port map( A => n1473, B => n1474, C => n1475, Y => n1477);
   U1513 : NAND2X1 port map( A => n1534, B => n262, Y => n1476);
   U1514 : OAI21X1 port map( A => n1493, B => n1477, C => n1476, Y => n1478);
   U1515 : OAI21X1 port map( A => n1479, B => n1478, C => n147, Y => n1485);
   U1516 : OAI22X1 port map( A => n251, B => n27, C => n275, D => n65, Y => 
                           n1483);
   U1517 : AOI21X1 port map( A => currentPlainKey_57_port, B => n266, C => 
                           n1483, Y => n1484);
   U1518 : NAND2X1 port map( A => n1485, B => n1484, Y => n1843);
   U1519 : NAND2X1 port map( A => n1515, B => n279, Y => n1502);
   U1520 : NAND2X1 port map( A => n244, B => n1571, Y => n1495);
   U1521 : NAND2X1 port map( A => n159, B => n1557, Y => n1487);
   U1522 : AOI22X1 port map( A => currentPlainKey_58_port, B => n1487, C => 
                           n1557, D => n1486, Y => n1489);
   U1523 : NAND2X1 port map( A => n1488, B => n1561, Y => n1524);
   U1524 : NAND2X1 port map( A => n1490, B => n63, Y => n1491);
   U1525 : NAND2X1 port map( A => n229, B => n1492, Y => n1494);
   U1526 : AOI21X1 port map( A => n1495, B => n1494, C => n1493, Y => n1496);
   U1527 : MUX2X1 port map( B => n1496, A => n260, S => n1552, Y => n1498);
   U1528 : NAND2X1 port map( A => n1534, B => n254, Y => n1497);
   U1529 : NAND2X1 port map( A => n1498, B => n1497, Y => n1499);
   U1530 : MUX2X1 port map( B => n1499, A => n248, S => n1437, Y => n1501);
   U1531 : NAND2X1 port map( A => currentPlainKey_58_port, B => n270, Y => 
                           n1500);
   U1532 : NAND3X1 port map( A => n1502, B => n1501, C => n1500, Y => n1844);
   U1533 : NAND2X1 port map( A => n1534, B => n278, Y => n1518);
   U1534 : OAI22X1 port map( A => n256, B => n7, C => n264, D => n63, Y => 
                           n1514);
   U1535 : NOR2X1 port map( A => n283, B => n1524, Y => n1511);
   U1536 : NOR2X1 port map( A => n61, B => n202, Y => n1507);
   U1537 : MUX2X1 port map( B => n1700, A => n1761, S => n1507, Y => n1508);
   U1538 : NAND2X1 port map( A => n1508, B => n1524, Y => n1509);
   U1539 : NAND2X1 port map( A => n174, B => n1561, Y => n1568);
   U1540 : INVX2 port map( A => n1568, Y => n1592);
   U1541 : MUX2X1 port map( B => n1509, A => n271, S => n1592, Y => n1510);
   U1542 : NOR2X1 port map( A => n1511, B => n1510, Y => n1512);
   U1543 : OAI22X1 port map( A => n1512, B => n143, C => n1589, D => n17, Y => 
                           n1513);
   U1544 : OAI21X1 port map( A => n1514, B => n1513, C => n119, Y => n1517);
   U1545 : AOI22X1 port map( A => n1515, B => n246, C => 
                           currentPlainKey_59_port, D => n267, Y => n1516);
   U1546 : NAND3X1 port map( A => n1518, B => n1517, C => n1516, Y => n1845);
   U1547 : AOI22X1 port map( A => n1552, B => n279, C => 
                           currentPlainKey_60_port, D => n270, Y => n1537);
   U1548 : AOI22X1 port map( A => n1592, B => n281, C => n1596, D => 
                           RCV_DATA(3), Y => n1528);
   U1549 : NAND2X1 port map( A => n162, B => n1557, Y => n1523);
   U1550 : INVX2 port map( A => n1521, Y => n1522);
   U1551 : AOI22X1 port map( A => currentPlainKey_60_port, B => n1523, C => 
                           n1522, D => n1557, Y => n1525);
   U1552 : NAND2X1 port map( A => n1568, B => n1524, Y => n1538);
   U1553 : NOR2X1 port map( A => n1525, B => n1538, Y => n1526);
   U1554 : NAND2X1 port map( A => n175, B => n1561, Y => n1540);
   U1555 : INVX2 port map( A => n1540, Y => n1590);
   U1556 : MUX2X1 port map( B => n1526, A => RCV_DATA(1), S => n1590, Y => 
                           n1527);
   U1557 : NAND2X1 port map( A => n1528, B => n1527, Y => n1531);
   U1558 : NOR2X1 port map( A => n265, B => n1529, Y => n1530);
   U1559 : AOI21X1 port map( A => n1551, B => n1531, C => n1530, Y => n1533);
   U1560 : NAND2X1 port map( A => n255, B => n1571, Y => n1532);
   U1561 : NAND2X1 port map( A => n1533, B => n1532, Y => n1535);
   U1562 : MUX2X1 port map( B => n1535, A => n248, S => n1534, Y => n1536);
   U1563 : NAND2X1 port map( A => n1537, B => n1536, Y => n1846);
   U1564 : NAND2X1 port map( A => n157, B => n1561, Y => n1587);
   U1565 : INVX2 port map( A => n1538, Y => n1539);
   U1566 : NAND3X1 port map( A => n1587, B => n1540, C => n1539, Y => n1541);
   U1567 : INVX2 port map( A => n1541, Y => n1565);
   U1568 : OAI21X1 port map( A => n61, B => n206, C => currentPlainKey_61_port,
                           Y => n1543);
   U1569 : OAI21X1 port map( A => n61, B => n1544, C => n1543, Y => n1546);
   U1570 : NOR2X1 port map( A => n271, B => n1587, Y => n1545);
   U1571 : AOI21X1 port map( A => n1565, B => n1546, C => n1545, Y => n1549);
   U1572 : NAND2X1 port map( A => n1590, B => n281, Y => n1548);
   U1573 : AOI22X1 port map( A => n1592, B => RCV_DATA(3), C => n1596, D => 
                           RCV_DATA(4), Y => n1547);
   U1574 : NAND3X1 port map( A => n1549, B => n1548, C => n1547, Y => n1550);
   U1575 : AOI22X1 port map( A => n115, B => RCV_DATA(5), C => n1551, D => 
                           n1550, Y => n1555);
   U1576 : NAND2X1 port map( A => n280, B => n1571, Y => n1554);
   U1577 : AOI22X1 port map( A => n1552, B => n246, C => 
                           currentPlainKey_61_port, D => n267, Y => n1553);
   U1578 : NAND3X1 port map( A => n1555, B => n1554, C => n1553, Y => n1847);
   U1579 : AOI22X1 port map( A => n246, B => n1571, C => n269, D => 
                           currentPlainKey_62_port, Y => n1576);
   U1580 : INVX2 port map( A => n1556, Y => n1560);
   U1581 : AOI21X1 port map( A => n186, B => n1557, C => n1685, Y => n1559);
   U1582 : NAND2X1 port map( A => n61, B => n1685, Y => n1558);
   U1583 : OAI21X1 port map( A => n1560, B => n1559, C => n1558, Y => n1562);
   U1584 : MUX2X1 port map( B => n1562, A => n271, S => n170, Y => n1564);
   U1585 : NOR2X1 port map( A => n283, B => n1587, Y => n1563);
   U1586 : AOI21X1 port map( A => n1565, B => n1564, C => n1563, Y => n1567);
   U1587 : NAND2X1 port map( A => n1590, B => RCV_DATA(3), Y => n1566);
   U1588 : NAND2X1 port map( A => n1567, B => n1566, Y => n1570);
   U1589 : NOR2X1 port map( A => n265, B => n1568, Y => n1569);
   U1590 : AOI21X1 port map( A => n227, B => n1570, C => n1569, Y => n1573);
   U1591 : NAND2X1 port map( A => n1596, B => n254, Y => n1572);
   U1592 : AOI21X1 port map( A => n1573, B => n1572, C => n1571, Y => n1574);
   U1593 : MUX2X1 port map( B => n1574, A => n278, S => n1598, Y => n1575);
   U1594 : NAND2X1 port map( A => n1576, B => n1575, Y => n1848);
   U1595 : NAND2X1 port map( A => n266, B => currentPlainKey_63_port, Y => 
                           n1601);
   U1596 : INVX2 port map( A => n1761, Y => n1580);
   U1597 : NOR2X1 port map( A => n1578, B => n204, Y => n1579);
   U1598 : MUX2X1 port map( B => currentPlainKey_63_port, A => n1580, S => 
                           n1579, Y => n1585);
   U1599 : NOR2X1 port map( A => n1582, B => n1581, Y => n1583);
   U1600 : MUX2X1 port map( B => n1585, A => n271, S => n1583, Y => n1586);
   U1601 : MUX2X1 port map( B => n1586, A => n281, S => n170, Y => n1588);
   U1602 : MUX2X1 port map( B => n1589, A => n1588, S => n1587, Y => n1591);
   U1603 : MUX2X1 port map( B => n1591, A => RCV_DATA(4), S => n1590, Y => 
                           n1594);
   U1604 : INVX2 port map( A => RCV_DATA(5), Y => n1593);
   U1605 : MUX2X1 port map( B => n1594, A => n1593, S => n1592, Y => n1595);
   U1606 : NAND2X1 port map( A => n229, B => n1595, Y => n1597);
   U1607 : MUX2X1 port map( B => n1597, A => n276, S => n1596, Y => n1599);
   U1608 : MUX2X1 port map( B => n1599, A => n247, S => n1598, Y => n1600);
   U1609 : NAND2X1 port map( A => n1601, B => n1600, Y => n1849);
   U1610 : NAND2X1 port map( A => n1669, B => n1602, Y => n1614);
   U1611 : INVX2 port map( A => n1614, Y => n1603);
   U1612 : NAND3X1 port map( A => n1603, B => n292, C => n1663, Y => n1612);
   U1613 : NAND2X1 port map( A => n160, B => n166, Y => n1604);
   U1614 : NAND2X1 port map( A => n1613, B => n1604, Y => n1785);
   U1615 : NAND2X1 port map( A => n151, B => n166, Y => n1605);
   U1616 : NAND2X1 port map( A => n1613, B => n1605, Y => n1784);
   U1617 : NAND2X1 port map( A => n105, B => n166, Y => n1606);
   U1618 : NAND2X1 port map( A => n1613, B => n1606, Y => n1783);
   U1619 : MUX2X1 port map( B => n222, A => keyCount_0_port, S => n1609, Y => 
                           n1607);
   U1620 : NAND2X1 port map( A => n1613, B => n1607, Y => n1782);
   U1621 : MUX2X1 port map( B => address_4_port, A => keyCount_1_port, S => 
                           n1609, Y => n1608);
   U1622 : NAND2X1 port map( A => n1613, B => n1608, Y => n1781);
   U1623 : MUX2X1 port map( B => address_5_port, A => keyCount_2_port, S => 
                           n1609, Y => n1610);
   U1624 : NAND2X1 port map( A => n1613, B => n1610, Y => n1780);
   U1625 : OAI21X1 port map( A => n1696, B => n1611, C => n1613, Y => n1779);
   U1626 : OAI21X1 port map( A => n1695, B => n1611, C => n1613, Y => n1778);
   U1627 : OAI21X1 port map( A => n1615, B => n1614, C => parityError, Y => 
                           n1618);
   U1628 : INVX2 port map( A => n1663, Y => n1616);
   U1629 : OAI21X1 port map( A => n1988, B => n1987, C => n1616, Y => n1617);
   U1630 : NAND2X1 port map( A => n1618, B => n1617, Y => nextParityError);
   U1631 : OAI21X1 port map( A => keyCount_0_port, B => n198, C => n1683, Y => 
                           n1619);
   U1632 : INVX2 port map( A => n1619, Y => n1671);
   U1633 : NAND2X1 port map( A => n1660, B => n1683, Y => n1684);
   U1634 : INVX2 port map( A => n1684, Y => n1674);
   U1635 : NAND2X1 port map( A => keyCount_0_port, B => n1674, Y => n1679);
   U1636 : MUX2X1 port map( B => n1671, A => n1679, S => n1694, Y => n1768);
   U1637 : NAND3X1 port map( A => n1661, B => n23, C => n1663, Y => n1622);
   U1638 : NAND3X1 port map( A => n1620, B => n292, C => n1657, Y => n1621);
   U1639 : OR2X2 port map( A => n1622, B => n1621, Y => n1635);
   U1640 : NAND2X1 port map( A => n1638, B => CLR_RBUFF_port, Y => n1637);
   U1641 : INVX2 port map( A => n1637, Y => n1633);
   U1642 : NAND2X1 port map( A => N1799, B => n1633, Y => n1624);
   U1643 : NAND2X1 port map( A => parityAccumulator_7_port, B => n1635, Y => 
                           n1623);
   U1644 : NAND2X1 port map( A => n1624, B => n1623, Y => n1777);
   U1645 : NAND2X1 port map( A => N1798, B => n1633, Y => n1626);
   U1646 : NAND2X1 port map( A => parityAccumulator_6_port, B => n1635, Y => 
                           n1625);
   U1647 : NAND2X1 port map( A => n1626, B => n1625, Y => n1776);
   U1648 : NAND2X1 port map( A => N1797, B => n1633, Y => n1628);
   U1649 : NAND2X1 port map( A => n1635, B => parityAccumulator_5_port, Y => 
                           n1627);
   U1650 : NAND2X1 port map( A => n1628, B => n1627, Y => n1775);
   U1651 : NAND2X1 port map( A => N1796, B => n1633, Y => n1630);
   U1652 : NAND2X1 port map( A => n1635, B => parityAccumulator_4_port, Y => 
                           n1629);
   U1653 : NAND2X1 port map( A => n1630, B => n1629, Y => n1774);
   U1654 : NAND2X1 port map( A => N1795, B => n1633, Y => n1631);
   U1655 : OAI21X1 port map( A => n1691, B => n1638, C => n1631, Y => n1773);
   U1656 : NAND2X1 port map( A => N1794, B => n1633, Y => n1632);
   U1657 : OAI21X1 port map( A => n1690, B => n1638, C => n1632, Y => n1772);
   U1658 : NAND2X1 port map( A => N1793, B => n1633, Y => n1634);
   U1659 : OAI21X1 port map( A => n1689, B => n1638, C => n1634, Y => n1771);
   U1660 : INVX2 port map( A => n1635, Y => n1638);
   U1661 : INVX2 port map( A => N1792, Y => n1636);
   U1662 : OAI22X1 port map( A => n1688, B => n1638, C => n1637, D => n1636, Y 
                           => n1770);
   U1663 : AOI21X1 port map( A => n1644, B => RBUF_FULL, C => n1920, Y => n1639
                           );
   U1664 : NAND2X1 port map( A => n1639, B => n1651, Y => n1640);
   U1665 : OAI21X1 port map( A => n224, B => n193, C => n1662, Y => n1645);
   U1666 : NAND2X1 port map( A => n1640, B => n1645, Y => n1655);
   U1667 : NAND2X1 port map( A => n224, B => n1655, Y => n1641);
   U1668 : NAND2X1 port map( A => n1642, B => n1641, Y => n1764);
   U1669 : INVX2 port map( A => keyCount_3_port, Y => n1644);
   U1670 : AND2X2 port map( A => keyCount_2_port, B => keyCount_0_port, Y => 
                           n1643);
   U1671 : NAND3X1 port map( A => keyCount_1_port, B => n1644, C => n1643, Y =>
                           n1659);
   U1672 : INVX2 port map( A => n1659, Y => n1675);
   U1673 : INVX2 port map( A => n1645, Y => n1658);
   U1674 : AOI22X1 port map( A => n1675, B => n1660, C => n1658, D => n225, Y 
                           => n1654);
   U1675 : INVX2 port map( A => RBUF_FULL, Y => n1646);
   U1676 : NAND2X1 port map( A => n1647, B => n1646, Y => n1653);
   U1677 : INVX2 port map( A => OE, Y => n1648);
   U1678 : NAND2X1 port map( A => n1760, B => n1648, Y => n1650);
   U1679 : NAND2X1 port map( A => n1661, B => n1663, Y => n1649);
   U1680 : AOI21X1 port map( A => n1651, B => n1650, C => n1649, Y => n1652);
   U1681 : NAND3X1 port map( A => n1654, B => n1653, C => n1652, Y => n1766);
   U1682 : AOI21X1 port map( A => n226, B => n1655, C => n1660, Y => n1656);
   U1683 : NAND3X1 port map( A => n1661, B => n1657, C => n1656, Y => n1767);
   U1684 : AOI22X1 port map( A => n1660, B => n1659, C => n1658, D => n164, Y 
                           => n1670);
   U1685 : NAND2X1 port map( A => n1662, B => n1661, Y => n1667);
   U1686 : NAND2X1 port map( A => n1760, B => n1648, Y => n1665);
   U1687 : OAI21X1 port map( A => n1665, B => n23, C => n1663, Y => n1666);
   U1688 : AOI21X1 port map( A => RBUF_FULL, B => n1667, C => n1666, Y => n1668
                           );
   U1689 : NAND3X1 port map( A => n1670, B => n1669, C => n1668, Y => n1765);
   U1690 : NOR2X1 port map( A => keyCount_2_port, B => n198, Y => n1673);
   U1691 : OAI21X1 port map( A => keyCount_1_port, B => n198, C => n1671, Y => 
                           n1678);
   U1692 : OAI21X1 port map( A => n1673, B => n1678, C => keyCount_3_port, Y =>
                           n1677);
   U1693 : NAND2X1 port map( A => n1675, B => n1674, Y => n1676);
   U1694 : NAND2X1 port map( A => n1677, B => n1676, Y => n1763);
   U1695 : INVX2 port map( A => n1678, Y => n1682);
   U1696 : INVX2 port map( A => n1679, Y => n1680);
   U1697 : NAND2X1 port map( A => n1680, B => keyCount_1_port, Y => n1681);
   U1698 : MUX2X1 port map( B => n1682, A => n1681, S => n1686, Y => n1769);
   U1699 : MUX2X1 port map( B => n1684, A => n1683, S => keyCount_0_port, Y => 
                           n1762);
   U1700 : INVX2 port map( A => keyCount_2_port, Y => n1686);
   U1701 : INVX2 port map( A => parityAccumulator_0_port, Y => n1688);
   U1702 : INVX2 port map( A => parityAccumulator_1_port, Y => n1689);
   U1703 : INVX2 port map( A => parityAccumulator_2_port, Y => n1690);
   U1704 : INVX2 port map( A => parityAccumulator_3_port, Y => n1691);
   U1705 : INVX2 port map( A => keyCount_1_port, Y => n1694);
   U1706 : INVX2 port map( A => address_7_port, Y => n1695);
   U1707 : INVX2 port map( A => currentPlainKey_61_port, Y => n1698);
   U1708 : INVX2 port map( A => currentPlainKey_60_port, Y => n1699);
   U1709 : INVX2 port map( A => currentPlainKey_59_port, Y => n1700);
   U1710 : INVX2 port map( A => currentPlainKey_58_port, Y => n1701);
   U1711 : INVX2 port map( A => currentPlainKey_57_port, Y => n1702);
   U1712 : INVX2 port map( A => currentPlainKey_56_port, Y => n1703);
   U1713 : INVX2 port map( A => currentPlainKey_55_port, Y => n1704);
   U1714 : INVX2 port map( A => currentPlainKey_54_port, Y => n1705);
   U1715 : INVX2 port map( A => currentPlainKey_53_port, Y => n1706);
   U1716 : INVX2 port map( A => currentPlainKey_52_port, Y => n1707);
   U1717 : INVX2 port map( A => currentPlainKey_51_port, Y => n1708);
   U1718 : INVX2 port map( A => currentPlainKey_50_port, Y => n1709);
   U1719 : INVX2 port map( A => currentPlainKey_49_port, Y => n1710);
   U1720 : INVX2 port map( A => currentPlainKey_48_port, Y => n1711);
   U1721 : INVX2 port map( A => currentPlainKey_47_port, Y => n1712);
   U1722 : INVX2 port map( A => currentPlainKey_46_port, Y => n1713);
   U1723 : INVX2 port map( A => currentPlainKey_45_port, Y => n1714);
   U1724 : INVX2 port map( A => currentPlainKey_44_port, Y => n1715);
   U1725 : INVX2 port map( A => currentPlainKey_43_port, Y => n1716);
   U1726 : INVX2 port map( A => currentPlainKey_42_port, Y => n1717);
   U1727 : INVX2 port map( A => currentPlainKey_41_port, Y => n1718);
   U1728 : INVX2 port map( A => currentPlainKey_40_port, Y => n1719);
   U1729 : INVX2 port map( A => currentPlainKey_39_port, Y => n1720);
   U1730 : INVX2 port map( A => currentPlainKey_38_port, Y => n1721);
   U1731 : INVX2 port map( A => currentPlainKey_37_port, Y => n1722);
   U1732 : INVX2 port map( A => currentPlainKey_36_port, Y => n1723);
   U1733 : INVX2 port map( A => currentPlainKey_35_port, Y => n1724);
   U1734 : INVX2 port map( A => currentPlainKey_34_port, Y => n1725);
   U1735 : INVX2 port map( A => currentPlainKey_33_port, Y => n1726);
   U1736 : INVX2 port map( A => currentPlainKey_32_port, Y => n1727);
   U1737 : INVX2 port map( A => currentPlainKey_31_port, Y => n1728);
   U1738 : INVX2 port map( A => currentPlainKey_30_port, Y => n1729);
   U1739 : INVX2 port map( A => currentPlainKey_29_port, Y => n1730);
   U1740 : INVX2 port map( A => currentPlainKey_28_port, Y => n1731);
   U1741 : INVX2 port map( A => currentPlainKey_27_port, Y => n1732);
   U1742 : INVX2 port map( A => currentPlainKey_26_port, Y => n1733);
   U1743 : INVX2 port map( A => currentPlainKey_25_port, Y => n1734);
   U1744 : INVX2 port map( A => currentPlainKey_24_port, Y => n1735);
   U1745 : INVX2 port map( A => currentPlainKey_23_port, Y => n1736);
   U1746 : INVX2 port map( A => currentPlainKey_22_port, Y => n1737);
   U1747 : INVX2 port map( A => currentPlainKey_21_port, Y => n1738);
   U1748 : INVX2 port map( A => currentPlainKey_20_port, Y => n1739);
   U1749 : INVX2 port map( A => currentPlainKey_19_port, Y => n1740);
   U1750 : INVX2 port map( A => currentPlainKey_18_port, Y => n1741);
   U1751 : INVX2 port map( A => currentPlainKey_17_port, Y => n1742);
   U1752 : INVX2 port map( A => currentPlainKey_16_port, Y => n1743);
   U1753 : INVX2 port map( A => currentPlainKey_15_port, Y => n1744);
   U1754 : INVX2 port map( A => currentPlainKey_14_port, Y => n1745);
   U1755 : INVX2 port map( A => currentPlainKey_13_port, Y => n1746);
   U1756 : INVX2 port map( A => currentPlainKey_12_port, Y => n1747);
   U1757 : INVX2 port map( A => currentPlainKey_11_port, Y => n1748);
   U1758 : INVX2 port map( A => currentPlainKey_10_port, Y => n1749);
   U1759 : INVX2 port map( A => currentPlainKey_9_port, Y => n1750);
   U1760 : INVX2 port map( A => currentPlainKey_8_port, Y => n1751);
   U1761 : INVX2 port map( A => currentPlainKey_7_port, Y => n1752);
   U1762 : INVX2 port map( A => currentPlainKey_6_port, Y => n1753);
   U1763 : INVX2 port map( A => currentPlainKey_5_port, Y => n1754);
   U1764 : INVX2 port map( A => currentPlainKey_4_port, Y => n1755);
   U1765 : INVX2 port map( A => SBE, Y => n1760);
   U1766 : INVX2 port map( A => n220, Y => n1761);

end SYN_keyb;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_sr_10bit_0 is

   port( CLK, RST, SHIFT_STROBE, SERIAL_IN : in std_logic;  LOAD_DATA : out 
         std_logic_vector (7 downto 0);  STOP_DATA : out std_logic_vector (1 
         downto 0));

end uart_sr_10bit_0;

architecture SYN_dataflow of uart_sr_10bit_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal LOAD_DATA_7_port, LOAD_DATA_6_port, LOAD_DATA_5_port, 
      LOAD_DATA_4_port, LOAD_DATA_3_port, LOAD_DATA_2_port, LOAD_DATA_1_port, 
      LOAD_DATA_0_port, STOP_DATA_1_port, STOP_DATA_0_port, n1, n2, n4, n5, n6,
      n7, n8, n9, n10, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48
      : std_logic;

begin
   LOAD_DATA <= ( LOAD_DATA_7_port, LOAD_DATA_6_port, LOAD_DATA_5_port, 
      LOAD_DATA_4_port, LOAD_DATA_3_port, LOAD_DATA_2_port, LOAD_DATA_1_port, 
      LOAD_DATA_0_port );
   STOP_DATA <= ( STOP_DATA_1_port, STOP_DATA_0_port );
   
   present_val_reg_9_inst : DFFSR port map( D => n36, CLK => CLK, R => n15, S 
                           => n37, Q => STOP_DATA_1_port);
   U2 : OAI21X1 port map( A => n35, B => n17, C => n48, Y => n46);
   U3 : NAND2X1 port map( A => LOAD_DATA_0_port, B => n17, Y => n48);
   U4 : OAI22X1 port map( A => n17, B => n34, C => n13, D => n35, Y => n45);
   U6 : OAI22X1 port map( A => n17, B => n31, C => n13, D => n34, Y => n44);
   U8 : OAI22X1 port map( A => n17, B => n29, C => n13, D => n31, Y => n43);
   U10 : OAI22X1 port map( A => n17, B => n27, C => n13, D => n29, Y => n42);
   U12 : OAI22X1 port map( A => n17, B => n25, C => n13, D => n27, Y => n41);
   U14 : OAI22X1 port map( A => n17, B => n23, C => n13, D => n25, Y => n40);
   U16 : OAI22X1 port map( A => n17, B => n21, C => n13, D => n23, Y => n39);
   U18 : OAI22X1 port map( A => n17, B => n19, C => n13, D => n21, Y => n38);
   U22 : OAI21X1 port map( A => n13, B => n19, C => n47, Y => n36);
   U23 : NAND2X1 port map( A => SERIAL_IN, B => n13, Y => n47);
   n37 <= '1';
   present_val_reg_8_inst : DFFSR port map( D => n38, CLK => CLK, R => n15, S 
                           => n10, Q => STOP_DATA_0_port);
   present_val_reg_7_inst : DFFSR port map( D => n39, CLK => CLK, R => n15, S 
                           => n9, Q => LOAD_DATA_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n40, CLK => CLK, R => n15, S 
                           => n8, Q => LOAD_DATA_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n41, CLK => CLK, R => n15, S 
                           => n7, Q => LOAD_DATA_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n42, CLK => CLK, R => n15, S 
                           => n6, Q => LOAD_DATA_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n43, CLK => CLK, R => n15, S 
                           => n5, Q => LOAD_DATA_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n44, CLK => CLK, R => n15, S 
                           => n4, Q => LOAD_DATA_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n45, CLK => CLK, R => n15, S 
                           => n2, Q => LOAD_DATA_1_port);
   present_val_reg_0_inst : DFFSR port map( D => n46, CLK => CLK, R => n15, S 
                           => n1, Q => LOAD_DATA_0_port);
   n1 <= '1';
   n2 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   U21 : INVX2 port map( A => RST, Y => n15);
   U24 : INVX2 port map( A => n13, Y => n17);
   U25 : INVX4 port map( A => n11, Y => n13);
   U26 : INVX2 port map( A => SHIFT_STROBE, Y => n11);
   U27 : INVX2 port map( A => STOP_DATA_1_port, Y => n19);
   U28 : INVX2 port map( A => STOP_DATA_0_port, Y => n21);
   U29 : INVX2 port map( A => LOAD_DATA_7_port, Y => n23);
   U30 : INVX2 port map( A => LOAD_DATA_6_port, Y => n25);
   U31 : INVX2 port map( A => LOAD_DATA_5_port, Y => n27);
   U32 : INVX2 port map( A => LOAD_DATA_4_port, Y => n29);
   U33 : INVX2 port map( A => LOAD_DATA_3_port, Y => n31);
   U35 : INVX2 port map( A => LOAD_DATA_2_port, Y => n34);
   U36 : INVX2 port map( A => LOAD_DATA_1_port, Y => n35);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_sb_check_0 is

   port( RST, CLK, SBC_CLR, SBC_EN : in std_logic;  STOP_DATA : in 
         std_logic_vector (1 downto 0);  SB_DETECT, SBE : out std_logic);

end uart_sb_check_0;

architecture SYN_behavioral of uart_sb_check_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal SBE_prime, sb_detect_flag, n2, n4, n5, n6, n10, n11, n12, n13, n14 : 
      std_logic;

begin
   
   SB_DETECT_reg : DFFSR port map( D => sb_detect_flag, CLK => CLK, R => n2, S 
                           => n13, Q => SB_DETECT);
   SBE_reg : DFFSR port map( D => SBE_prime, CLK => CLK, R => n2, S => n14, Q 
                           => SBE);
   n14 <= '1';
   n13 <= '1';
   U6 : OR2X2 port map( A => SBC_CLR, B => STOP_DATA(0), Y => n12);
   U10 : NOR2X1 port map( A => n12, B => n11, Y => sb_detect_flag);
   U11 : NAND2X1 port map( A => STOP_DATA(1), B => SBC_EN, Y => n11);
   U12 : NOR2X1 port map( A => n6, B => n10, Y => SBE_prime);
   U13 : OAI21X1 port map( A => STOP_DATA(0), B => n4, C => n5, Y => n10);
   U4 : INVX2 port map( A => RST, Y => n2);
   U7 : INVX2 port map( A => STOP_DATA(1), Y => n4);
   U8 : INVX2 port map( A => SBC_CLR, Y => n5);
   U9 : INVX2 port map( A => SBC_EN, Y => n6);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_buf_full_0 is

   port( CLK, RST, CLR_RBUF, SET_RBUF_FULL : in std_logic;  RBUF_FULL : out 
         std_logic);

end uart_rcv_buf_full_0;

architecture SYN_Behavioral of uart_rcv_buf_full_0 is

   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal RBUF_FULL_port, n4, n5, n6 : std_logic;

begin
   RBUF_FULL <= RBUF_FULL_port;
   
   Q_int_reg : DFFSR port map( D => n4, CLK => CLK, R => n6, S => n5, Q => 
                           RBUF_FULL_port);
   U3 : NOR2X1 port map( A => RST, B => CLR_RBUF, Y => n6);
   n5 <= '1';
   U4 : OR2X2 port map( A => RBUF_FULL_port, B => SET_RBUF_FULL, Y => n4);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_buf_0 is

   port( CLK, RST, LOAD_RBUF : in std_logic;  LOAD_DATA : in std_logic_vector 
         (7 downto 0);  RCV_DATA : out std_logic_vector (7 downto 0));

end uart_rcv_buf_0;

architecture SYN_Behavioral of uart_rcv_buf_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, n2, 
      n11, n12, n13, n15, n17, n19, n21, n23, n24, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41 : std_logic;

begin
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   Q_int_reg_7_inst : DFFSR port map( D => n12, CLK => CLK, R => n11, S => n27,
                           Q => RCV_DATA_7_port);
   Q_int_reg_6_inst : DFFSR port map( D => n13, CLK => CLK, R => n11, S => n28,
                           Q => RCV_DATA_6_port);
   Q_int_reg_5_inst : DFFSR port map( D => n15, CLK => CLK, R => n11, S => n29,
                           Q => RCV_DATA_5_port);
   Q_int_reg_4_inst : DFFSR port map( D => n17, CLK => CLK, R => n11, S => n30,
                           Q => RCV_DATA_4_port);
   Q_int_reg_3_inst : DFFSR port map( D => n19, CLK => CLK, R => n11, S => n31,
                           Q => RCV_DATA_3_port);
   Q_int_reg_2_inst : DFFSR port map( D => n21, CLK => CLK, R => n11, S => n32,
                           Q => RCV_DATA_2_port);
   Q_int_reg_0_inst : DFFSR port map( D => n24, CLK => CLK, R => n11, S => n33,
                           Q => RCV_DATA_0_port);
   U3 : AOI22X1 port map( A => LOAD_RBUF, B => LOAD_DATA(0), C => 
                           RCV_DATA_0_port, D => n26, Y => n41);
   U5 : AOI22X1 port map( A => LOAD_DATA(1), B => LOAD_RBUF, C => 
                           RCV_DATA_1_port, D => n26, Y => n40);
   U7 : AOI22X1 port map( A => LOAD_DATA(2), B => LOAD_RBUF, C => 
                           RCV_DATA_2_port, D => n26, Y => n39);
   U9 : AOI22X1 port map( A => LOAD_DATA(3), B => LOAD_RBUF, C => 
                           RCV_DATA_3_port, D => n26, Y => n38);
   U11 : AOI22X1 port map( A => LOAD_DATA(4), B => LOAD_RBUF, C => 
                           RCV_DATA_4_port, D => n26, Y => n37);
   U13 : AOI22X1 port map( A => LOAD_DATA(5), B => LOAD_RBUF, C => 
                           RCV_DATA_5_port, D => n26, Y => n36);
   U15 : AOI22X1 port map( A => LOAD_DATA(6), B => LOAD_RBUF, C => 
                           RCV_DATA_6_port, D => n26, Y => n35);
   U18 : AOI22X1 port map( A => LOAD_DATA(7), B => LOAD_RBUF, C => 
                           RCV_DATA_7_port, D => n26, Y => n34);
   n33 <= '1';
   n32 <= '1';
   n31 <= '1';
   n30 <= '1';
   n29 <= '1';
   n28 <= '1';
   n27 <= '1';
   Q_int_reg_1_inst : DFFSR port map( D => n23, CLK => CLK, R => n11, S => n2, 
                           Q => RCV_DATA_1_port);
   n2 <= '1';
   U4 : INVX2 port map( A => RST, Y => n11);
   U6 : INVX2 port map( A => n34, Y => n12);
   U8 : INVX2 port map( A => n35, Y => n13);
   U10 : INVX2 port map( A => n36, Y => n15);
   U12 : INVX2 port map( A => n37, Y => n17);
   U14 : INVX2 port map( A => n38, Y => n19);
   U16 : INVX2 port map( A => n39, Y => n21);
   U17 : INVX2 port map( A => n40, Y => n23);
   U19 : INVX2 port map( A => n41, Y => n24);
   U21 : INVX2 port map( A => LOAD_RBUF, Y => n26);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcu_0 is

   port( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT : in std_logic;  RBUF_LOAD
         , TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR : out 
         std_logic);

end uart_rcu_0;

architecture SYN_rcub of uart_rcu_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal RBUF_LOAD_port, TIMER_TRIG_port, CHK_ERROR_port, SET_RBUF_FULL_port, 
      SBC_EN_port, SBC_CLR_port, state_2_port, state_1_port, state_0_port, 
      timerRunning, count_7_port, count_6_port, count_5_port, count_4_port, 
      count_3_port, count_2_port, count_1_port, count_0_port, nextCount_7_port,
      nextCount_6_port, nextCount_5_port, nextCount_4_port, nextCount_3_port, 
      nextCount_2_port, nextCount_1_port, nextCount_0_port, nextState_1_port, 
      nextState_0_port, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, 
      N35, N36, N37, N38, N99, add_46_carry_3_port, add_46_carry_4_port, 
      add_46_carry_5_port, add_46_carry_6_port, n1, n2, n3, n4, n5, n6, n7, 
      n25_port, n32_port, n34_port, n35_port, n36_port, n37_port, n38_port, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99_port, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139 : std_logic;

begin
   RBUF_LOAD <= RBUF_LOAD_port;
   TIMER_TRIG <= TIMER_TRIG_port;
   CHK_ERROR <= CHK_ERROR_port;
   SET_RBUF_FULL <= SET_RBUF_FULL_port;
   SBC_EN <= SBC_EN_port;
   SBC_CLR <= SBC_CLR_port;
   
   count_reg_0_inst : DFFSR port map( D => nextCount_0_port, CLK => CLK, R => 
                           n5, S => n116, Q => count_0_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n4, S => n117, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => n43, CLK => CLK, R => n4, S => n118,
                           Q => state_2_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n4, S => n119, Q => state_0_port);
   SBC_CLR_reg : DFFSR port map( D => n85, CLK => CLK, R => n4, S => n120, Q =>
                           SBC_CLR_port);
   TIMER_TRIG_reg : DFFSR port map( D => n84, CLK => CLK, R => n4, S => n121, Q
                           => TIMER_TRIG_port);
   RBUF_LOAD_reg : DFFSR port map( D => n83, CLK => CLK, R => n4, S => n122, Q 
                           => RBUF_LOAD_port);
   timerRunning_reg : DFFSR port map( D => n89, CLK => CLK, R => n4, S => n123,
                           Q => timerRunning);
   nextCount_reg_1_inst : DFFSR port map( D => N32, CLK => CLK, R => n4, S => 
                           n124, Q => nextCount_1_port);
   count_reg_1_inst : DFFSR port map( D => nextCount_1_port, CLK => CLK, R => 
                           n4, S => n125, Q => count_1_port);
   nextCount_reg_0_inst : DFFSR port map( D => N31, CLK => CLK, R => n126, S =>
                           n5, Q => nextCount_0_port);
   nextCount_reg_2_inst : DFFSR port map( D => N33, CLK => CLK, R => n4, S => 
                           n127, Q => nextCount_2_port);
   count_reg_2_inst : DFFSR port map( D => nextCount_2_port, CLK => CLK, R => 
                           n5, S => n128, Q => count_2_port);
   nextCount_reg_3_inst : DFFSR port map( D => N34, CLK => CLK, R => n5, S => 
                           n129, Q => nextCount_3_port);
   count_reg_3_inst : DFFSR port map( D => nextCount_3_port, CLK => CLK, R => 
                           n5, S => n130, Q => count_3_port);
   nextCount_reg_4_inst : DFFSR port map( D => N35, CLK => CLK, R => n5, S => 
                           n131, Q => nextCount_4_port);
   count_reg_4_inst : DFFSR port map( D => nextCount_4_port, CLK => CLK, R => 
                           n5, S => n132, Q => count_4_port);
   nextCount_reg_5_inst : DFFSR port map( D => N36, CLK => CLK, R => n5, S => 
                           n133, Q => nextCount_5_port);
   count_reg_5_inst : DFFSR port map( D => nextCount_5_port, CLK => CLK, R => 
                           n5, S => n134, Q => count_5_port);
   nextCount_reg_6_inst : DFFSR port map( D => N37, CLK => CLK, R => n5, S => 
                           n135, Q => nextCount_6_port);
   count_reg_6_inst : DFFSR port map( D => nextCount_6_port, CLK => CLK, R => 
                           n5, S => n136, Q => count_6_port);
   nextCount_reg_7_inst : DFFSR port map( D => N38, CLK => CLK, R => n5, S => 
                           n137, Q => nextCount_7_port);
   count_reg_7_inst : DFFSR port map( D => nextCount_7_port, CLK => CLK, R => 
                           n5, S => n138, Q => count_7_port);
   SBC_EN_reg : DFFSR port map( D => n87, CLK => CLK, R => n4, S => n139, Q => 
                           SBC_EN_port);
   n139 <= '1';
   n138 <= '1';
   n137 <= '1';
   n136 <= '1';
   n135 <= '1';
   n134 <= '1';
   n133 <= '1';
   n132 <= '1';
   n131 <= '1';
   n130 <= '1';
   n129 <= '1';
   n128 <= '1';
   n127 <= '1';
   n126 <= '1';
   n125 <= '1';
   n124 <= '1';
   n123 <= '1';
   n122 <= '1';
   n121 <= '1';
   n120 <= '1';
   n119 <= '1';
   n118 <= '1';
   n117 <= '1';
   n116 <= '1';
   U33 : AND2X2 port map( A => N30, B => timerRunning, Y => N38);
   U34 : AND2X2 port map( A => N29, B => timerRunning, Y => N37);
   U35 : AND2X2 port map( A => N28, B => timerRunning, Y => N36);
   U36 : AND2X2 port map( A => N27, B => timerRunning, Y => N35);
   U37 : AND2X2 port map( A => N26, B => timerRunning, Y => N34);
   U38 : AND2X2 port map( A => N25, B => timerRunning, Y => N33);
   U39 : AND2X2 port map( A => N24, B => timerRunning, Y => N32);
   U54 : OAI21X1 port map( A => n114, B => n45, C => n113, Y => n115);
   U55 : OAI21X1 port map( A => n46, B => n44, C => n45, Y => n113);
   U56 : NAND2X1 port map( A => n112, B => n111, Y => n89);
   U57 : OAI21X1 port map( A => n110, B => n109, C => timerRunning, Y => n111);
   U58 : NAND2X1 port map( A => n108, B => n107, Y => n109);
   U59 : NAND2X1 port map( A => n106, B => n107, Y => n88);
   U60 : NAND3X1 port map( A => n37_port, B => n112, C => CHK_ERROR_port, Y => 
                           n106);
   U61 : OAI21X1 port map( A => n105, B => n82, C => n104, Y => n87);
   U62 : NAND2X1 port map( A => n107, B => n103, Y => n105);
   U63 : NAND2X1 port map( A => n102, B => n40, Y => n107);
   U64 : NAND3X1 port map( A => n101, B => n100, C => n99_port, Y => n86);
   U65 : NAND3X1 port map( A => n36_port, B => n112, C => SET_RBUF_FULL_port, Y
                           => n99_port);
   U66 : NAND2X1 port map( A => n103, B => n100, Y => n110);
   U67 : NAND3X1 port map( A => nextState_0_port, B => nextState_1_port, C => 
                           n102, Y => n100);
   U68 : NAND3X1 port map( A => n38_port, B => n40, C => n102, Y => n101);
   U69 : OAI21X1 port map( A => n98, B => n47, C => n112, Y => n85);
   U70 : OAI21X1 port map( A => n98, B => n81, C => n112, Y => n84);
   U71 : NAND2X1 port map( A => n103, B => n104, Y => n98);
   U72 : NAND3X1 port map( A => nextState_1_port, B => n38_port, C => n41, Y =>
                           n104);
   U73 : NAND2X1 port map( A => n97, B => n108, Y => n83);
   U74 : NAND3X1 port map( A => nextState_1_port, B => n38_port, C => n102, Y 
                           => n108);
   U75 : NAND3X1 port map( A => n103, B => n112, C => RBUF_LOAD_port, Y => n97)
                           ;
   U76 : NAND3X1 port map( A => nextState_0_port, B => n40, C => n41, Y => n112
                           );
   U77 : NAND3X1 port map( A => n38_port, B => n40, C => n41, Y => n103);
   U78 : OAI21X1 port map( A => n42, B => n45, C => n96, Y => n102);
   U79 : NAND3X1 port map( A => state_0_port, B => n45, C => state_1_port, Y =>
                           n96);
   U80 : NAND2X1 port map( A => n95, B => n94, Y => n114);
   U81 : OAI21X1 port map( A => n93, B => n94, C => n95, Y => nextState_1_port)
                           ;
   U82 : NOR2X1 port map( A => N99, B => state_2_port, Y => n93);
   U83 : OAI21X1 port map( A => state_2_port, B => n92, C => n95, Y => 
                           nextState_0_port);
   U84 : NAND2X1 port map( A => state_1_port, B => n46, Y => n95);
   U85 : AOI21X1 port map( A => START_BIT, B => n46, C => n91, Y => n92);
   U86 : OAI21X1 port map( A => N99, B => n94, C => n90, Y => n91);
   U87 : NAND2X1 port map( A => SB_DETECT, B => state_1_port, Y => n90);
   U88 : NAND2X1 port map( A => state_0_port, B => n44, Y => n94);
   U89 : NAND2X1 port map( A => n39, B => timerRunning, Y => N31);
   SET_RBUF_FULL_reg : DFFSR port map( D => n86, CLK => CLK, R => n4, S => n2, 
                           Q => SET_RBUF_FULL_port);
   CHK_ERROR_reg : DFFSR port map( D => n88, CLK => CLK, R => n4, S => n1, Q =>
                           CHK_ERROR_port);
   n1 <= '1';
   n2 <= '1';
   U7 : INVX2 port map( A => RST, Y => n4);
   U8 : INVX2 port map( A => RST, Y => n5);
   U24 : XNOR2X1 port map( A => count_7_port, B => n3, Y => N30);
   U31 : NAND2X1 port map( A => count_6_port, B => add_46_carry_6_port, Y => n3
                           );
   U40 : XOR2X1 port map( A => add_46_carry_6_port, B => count_6_port, Y => N29
                           );
   U41 : AND2X1 port map( A => count_5_port, B => add_46_carry_5_port, Y => 
                           add_46_carry_6_port);
   U42 : XOR2X1 port map( A => add_46_carry_5_port, B => count_5_port, Y => N28
                           );
   U43 : AND2X1 port map( A => count_4_port, B => add_46_carry_4_port, Y => 
                           add_46_carry_5_port);
   U44 : XOR2X1 port map( A => add_46_carry_4_port, B => count_4_port, Y => N27
                           );
   U45 : AND2X1 port map( A => count_3_port, B => add_46_carry_3_port, Y => 
                           add_46_carry_4_port);
   U46 : XOR2X1 port map( A => add_46_carry_3_port, B => count_3_port, Y => N26
                           );
   U47 : AND2X1 port map( A => count_2_port, B => count_1_port, Y => 
                           add_46_carry_3_port);
   U48 : XOR2X1 port map( A => count_1_port, B => count_2_port, Y => N25);
   U49 : INVX2 port map( A => count_1_port, Y => N24);
   U50 : OAI21X1 port map( A => count_0_port, B => count_1_port, C => 
                           count_2_port, Y => n6);
   U51 : NOR2X1 port map( A => n35_port, B => n6, Y => n7);
   U52 : OAI21X1 port map( A => n7, B => count_4_port, C => count_6_port, Y => 
                           n25_port);
   U53 : OAI21X1 port map( A => n34_port, B => n25_port, C => n32_port, Y => 
                           N99);
   U90 : INVX2 port map( A => count_7_port, Y => n32_port);
   U91 : INVX2 port map( A => count_5_port, Y => n34_port);
   U92 : INVX2 port map( A => count_3_port, Y => n35_port);
   U93 : INVX2 port map( A => n110, Y => n36_port);
   U94 : INVX2 port map( A => n105, Y => n37_port);
   U95 : INVX2 port map( A => nextState_0_port, Y => n38_port);
   U96 : INVX2 port map( A => count_0_port, Y => n39);
   U97 : INVX2 port map( A => nextState_1_port, Y => n40);
   U98 : INVX2 port map( A => n102, Y => n41);
   U99 : INVX2 port map( A => n114, Y => n42);
   U100 : INVX2 port map( A => n115, Y => n43);
   U101 : INVX2 port map( A => state_1_port, Y => n44);
   U102 : INVX2 port map( A => state_2_port, Y => n45);
   U103 : INVX2 port map( A => state_0_port, Y => n46);
   U104 : INVX2 port map( A => SBC_CLR_port, Y => n47);
   U105 : INVX2 port map( A => TIMER_TRIG_port, Y => n81);
   U106 : INVX2 port map( A => SBC_EN_port, Y => n82);

end SYN_rcub;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_error_0 is

   port( RST, CLK, RBUF_FULL, CHK_ERROR : in std_logic;  OE : out std_logic);

end uart_error_0;

architecture SYN_behavioral of uart_error_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal OE_prime, n1, n3 : std_logic;

begin
   
   OE_reg : DFFSR port map( D => OE_prime, CLK => CLK, R => n1, S => n3, Q => 
                           OE);
   n3 <= '1';
   U5 : AND2X2 port map( A => RBUF_FULL, B => CHK_ERROR, Y => OE_prime);
   U3 : INVX2 port map( A => RST, Y => n1);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_edge_detector_0 is

   port( CLK, RST, SERIAL_IN : in std_logic;  START_BIT : out std_logic);

end uart_edge_detector_0;

architecture SYN_Behavioral of uart_edge_detector_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal Q_int, Q_int2, n2, n4, n5, n6 : std_logic;

begin
   
   Q_int_reg : DFFSR port map( D => SERIAL_IN, CLK => CLK, R => n2, S => n5, Q 
                           => Q_int);
   Q_int2_reg : DFFSR port map( D => Q_int, CLK => CLK, R => n2, S => n6, Q => 
                           Q_int2);
   n6 <= '1';
   n5 <= '1';
   U7 : NOR2X1 port map( A => Q_int, B => n4, Y => START_BIT);
   U4 : INVX2 port map( A => RST, Y => n2);
   U6 : INVX2 port map( A => Q_int2, Y => n4);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_timer_0 is

   port( CLK, RST, SENDING : in std_logic;  SHIFT_ENABLE_R, SHIFT_ENABLE_E : 
         out std_logic);

end tx_timer_0;

architecture SYN_moore of tx_timer_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal count_3_port, count_2_port, count_1_port, count_0_port, state, 
      nextcount_3_port, nextcount_2_port, nextcount_1_port, nextcount_0_port, 
      nxt_SHIFT_ENABLE_E, n6, n8, n9, n10, n11, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34 : std_logic;

begin
   SHIFT_ENABLE_R <= nxt_SHIFT_ENABLE_E;
   
   state_reg : DFFSR port map( D => SENDING, CLK => CLK, R => n6, S => n29, Q 
                           => state);
   count_reg_0_inst : DFFSR port map( D => nextcount_0_port, CLK => CLK, R => 
                           n6, S => n30, Q => count_0_port);
   count_reg_2_inst : DFFSR port map( D => nextcount_2_port, CLK => CLK, R => 
                           n6, S => n31, Q => count_2_port);
   count_reg_1_inst : DFFSR port map( D => nextcount_1_port, CLK => CLK, R => 
                           n6, S => n32, Q => count_1_port);
   count_reg_3_inst : DFFSR port map( D => nextcount_3_port, CLK => CLK, R => 
                           n6, S => n33, Q => count_3_port);
   SHIFT_ENABLE_E_reg : DFFSR port map( D => nxt_SHIFT_ENABLE_E, CLK => CLK, R 
                           => n6, S => n34, Q => SHIFT_ENABLE_E);
   n34 <= '1';
   n33 <= '1';
   n32 <= '1';
   n31 <= '1';
   n30 <= '1';
   n29 <= '1';
   U14 : NOR2X1 port map( A => n28, B => n27, Y => nextcount_3_port);
   U15 : XNOR2X1 port map( A => count_3_port, B => n26, Y => n28);
   U16 : NOR2X1 port map( A => n25, B => n20, Y => n26);
   U17 : AOI21X1 port map( A => n24, B => state, C => n21, Y => 
                           nextcount_2_port);
   U18 : XNOR2X1 port map( A => n25, B => n20, Y => n24);
   U19 : NAND2X1 port map( A => count_1_port, B => count_0_port, Y => n25);
   U20 : NOR2X1 port map( A => n23, B => n27, Y => nextcount_1_port);
   U21 : NAND3X1 port map( A => SENDING, B => n22, C => state, Y => n27);
   U22 : XNOR2X1 port map( A => count_0_port, B => count_1_port, Y => n23);
   U23 : OAI21X1 port map( A => count_0_port, B => n21, C => state, Y => 
                           nextcount_0_port);
   U8 : INVX1 port map( A => SENDING, Y => n21);
   U10 : INVX2 port map( A => RST, Y => n6);
   U11 : NOR2X1 port map( A => count_0_port, B => count_2_port, Y => n9);
   U12 : INVX2 port map( A => count_1_port, Y => n8);
   U13 : NAND2X1 port map( A => n9, B => n8, Y => n22);
   U24 : INVX2 port map( A => n22, Y => n11);
   U25 : AND2X2 port map( A => count_3_port, B => state, Y => n10);
   U26 : NAND3X1 port map( A => SENDING, B => n11, C => n10, Y => n19);
   U27 : INVX2 port map( A => n19, Y => nxt_SHIFT_ENABLE_E);
   U28 : INVX2 port map( A => count_2_port, Y => n20);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_tcu_0 is

   port( clk, rst, p_ready, t_bitstuff : in std_logic;  PRGA_OUT : in 
         std_logic_vector (7 downto 0);  prga_opcode : in std_logic_vector (1 
         downto 0);  t_crc : in std_logic_vector (15 downto 0);  sending, EOP, 
         next_byte : out std_logic;  send_data : out std_logic_vector (7 downto
         0);  t_strobe : out std_logic);

end tx_tcu_0;

architecture SYN_behavioral of tx_tcu_0 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component tx_tcu_0_DW01_inc_0
      port( A : in std_logic_vector (6 downto 0);  SUM : out std_logic_vector 
            (6 downto 0));
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal send_data_7_port, send_data_6_port, send_data_5_port, 
      send_data_4_port, send_data_3_port, send_data_2_port, send_data_1_port, 
      send_data_0_port, state_2_port, state_1_port, state_0_port, count_5_port,
      count_4_port, count_3_port, count_2_port, count_1_port, count_0_port, 
      nextstate_2_port, nextstate_1_port, nextstate_0_port, flop_data_7_port, 
      flop_data_6_port, flop_data_5_port, flop_data_4_port, flop_data_3_port, 
      flop_data_2_port, flop_data_1_port, flop_data_0_port, 
      current_send_data_7_port, current_send_data_6_port, 
      current_send_data_5_port, current_send_data_4_port, 
      current_send_data_3_port, current_send_data_2_port, 
      current_send_data_1_port, current_send_data_0_port, N59, N60, N61, N62, 
      N63, N64, N65, N188, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59_port, n60_port, n61_port, n62_port, n63_port, n64_port, 
      n65_port, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n175, n177, n179, n184, n185, n186, n187, 
      n188_port, n189, n190, n191, n192, n193, n201, n202, n203, n204, n205, 
      n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
      n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
      n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290 : std_logic;

begin
   send_data <= ( send_data_7_port, send_data_6_port, send_data_5_port, 
      send_data_4_port, send_data_3_port, send_data_2_port, send_data_1_port, 
      send_data_0_port );
   
   count_reg_0_inst : DFFSR port map( D => n261, CLK => clk, R => n29, S => 
                           n268, Q => count_0_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n29, S => n269, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n29, S => n270, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n29, S => n271, Q => state_2_port);
   count_reg_1_inst : DFFSR port map( D => n267, CLK => clk, R => n29, S => 
                           n272, Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n266, CLK => clk, R => n29, S => 
                           n273, Q => count_2_port);
   count_reg_4_inst : DFFSR port map( D => n264, CLK => clk, R => n29, S => 
                           n274, Q => count_4_port);
   flop_data_reg_7_inst : DFFPOSX1 port map( D => n253, CLK => clk, Q => 
                           flop_data_7_port);
   current_send_data_reg_7_inst : DFFPOSX1 port map( D => n275, CLK => clk, Q 
                           => current_send_data_7_port);
   flop_data_reg_6_inst : DFFPOSX1 port map( D => n254, CLK => clk, Q => 
                           flop_data_6_port);
   current_send_data_reg_6_inst : DFFPOSX1 port map( D => n276, CLK => clk, Q 
                           => current_send_data_6_port);
   flop_data_reg_5_inst : DFFPOSX1 port map( D => n255, CLK => clk, Q => 
                           flop_data_5_port);
   current_send_data_reg_5_inst : DFFPOSX1 port map( D => n277, CLK => clk, Q 
                           => current_send_data_5_port);
   flop_data_reg_4_inst : DFFPOSX1 port map( D => n256, CLK => clk, Q => 
                           flop_data_4_port);
   current_send_data_reg_4_inst : DFFPOSX1 port map( D => n278, CLK => clk, Q 
                           => current_send_data_4_port);
   flop_data_reg_3_inst : DFFPOSX1 port map( D => n257, CLK => clk, Q => 
                           flop_data_3_port);
   current_send_data_reg_3_inst : DFFPOSX1 port map( D => n279, CLK => clk, Q 
                           => current_send_data_3_port);
   flop_data_reg_2_inst : DFFPOSX1 port map( D => n258, CLK => clk, Q => 
                           flop_data_2_port);
   current_send_data_reg_2_inst : DFFPOSX1 port map( D => n280, CLK => clk, Q 
                           => current_send_data_2_port);
   flop_data_reg_1_inst : DFFPOSX1 port map( D => n259, CLK => clk, Q => 
                           flop_data_1_port);
   current_send_data_reg_1_inst : DFFPOSX1 port map( D => n281, CLK => clk, Q 
                           => current_send_data_1_port);
   flop_data_reg_0_inst : DFFPOSX1 port map( D => n260, CLK => clk, Q => 
                           flop_data_0_port);
   current_send_data_reg_0_inst : DFFPOSX1 port map( D => n282, CLK => clk, Q 
                           => current_send_data_0_port);
   send_data_reg_7_inst : DFFPOSX1 port map( D => n283, CLK => clk, Q => 
                           send_data_7_port);
   send_data_reg_6_inst : DFFPOSX1 port map( D => n284, CLK => clk, Q => 
                           send_data_6_port);
   send_data_reg_5_inst : DFFPOSX1 port map( D => n285, CLK => clk, Q => 
                           send_data_5_port);
   send_data_reg_4_inst : DFFPOSX1 port map( D => n286, CLK => clk, Q => 
                           send_data_4_port);
   send_data_reg_3_inst : DFFPOSX1 port map( D => n287, CLK => clk, Q => 
                           send_data_3_port);
   send_data_reg_2_inst : DFFPOSX1 port map( D => n288, CLK => clk, Q => 
                           send_data_2_port);
   send_data_reg_1_inst : DFFPOSX1 port map( D => n289, CLK => clk, Q => 
                           send_data_1_port);
   send_data_reg_0_inst : DFFPOSX1 port map( D => n290, CLK => clk, Q => 
                           send_data_0_port);
   n274 <= '1';
   n273 <= '1';
   n272 <= '1';
   n271 <= '1';
   n270 <= '1';
   n269 <= '1';
   n268 <= '1';
   r80 : tx_tcu_0_DW01_inc_0 port map( A(6) => n27, A(5) => n7, A(4) => n8, 
                           A(3) => n9, A(2) => n6, A(1) => n13, A(0) => 
                           count_0_port, SUM(6) => N65, SUM(5) => N64, SUM(4) 
                           => N63, SUM(3) => N62, SUM(2) => N61, SUM(1) => N60,
                           SUM(0) => N59);
   count_reg_6_inst : DFFSR port map( D => n262, CLK => clk, R => n29, S => n4,
                           Q => N188);
   count_reg_3_inst : DFFSR port map( D => n265, CLK => clk, R => n29, S => n3,
                           Q => count_3_port);
   count_reg_5_inst : DFFSR port map( D => n263, CLK => clk, R => n29, S => n2,
                           Q => count_5_port);
   U3 : INVX2 port map( A => n11, Y => n13);
   U4 : INVX4 port map( A => n28, Y => n36);
   U5 : INVX2 port map( A => n187, Y => n19);
   U6 : INVX2 port map( A => count_0_port, Y => n175);
   U7 : NAND2X1 port map( A => n14, B => n112, Y => n1);
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   U11 : INVX2 port map( A => n125, Y => n5);
   U12 : INVX1 port map( A => n191, Y => n6);
   U13 : INVX2 port map( A => n154, Y => n7);
   U14 : BUFX4 port map( A => count_4_port, Y => n8);
   U15 : BUFX4 port map( A => count_3_port, Y => n9);
   U16 : INVX1 port map( A => n147, Y => n10);
   U17 : INVX2 port map( A => count_1_port, Y => n11);
   U18 : INVX1 port map( A => n11, Y => n12);
   U19 : INVX1 port map( A => n20, Y => n137);
   U20 : AND2X2 port map( A => n120, B => n112, Y => n15);
   U21 : INVX2 port map( A => n111, Y => n14);
   U22 : NAND2X1 port map( A => n9, B => count_0_port, Y => n16);
   U23 : NAND2X1 port map( A => n201, B => n17, Y => n192);
   U24 : INVX2 port map( A => n16, Y => n17);
   U25 : INVX2 port map( A => count_3_port, Y => n190);
   U26 : INVX1 port map( A => n248, Y => n62_port);
   U27 : AND2X2 port map( A => n132, B => n94, Y => n18);
   U28 : INVX4 port map( A => n18, Y => n147);
   U29 : INVX1 port map( A => n109, Y => n110);
   U30 : OR2X2 port map( A => n20, B => n19, Y => n140);
   U31 : INVX2 port map( A => n20, Y => n186);
   U32 : INVX1 port map( A => n127, Y => n138);
   U33 : INVX1 port map( A => n65_port, Y => n34);
   U34 : AND2X2 port map( A => n6, B => n24, Y => n25);
   U35 : OR2X2 port map( A => n192, B => n193, Y => n20);
   U36 : INVX1 port map( A => n141, Y => n90);
   U37 : AND2X1 port map( A => n13, B => n22, Y => n24);
   U38 : INVX1 port map( A => n93, Y => n125);
   U39 : INVX2 port map( A => count_2_port, Y => n191);
   U40 : INVX1 port map( A => n140, Y => n126);
   U41 : AND2X1 port map( A => n185, B => n125, Y => n21);
   U42 : INVX2 port map( A => rst, Y => n29);
   U43 : NOR2X1 port map( A => t_bitstuff, B => n175, Y => n22);
   U44 : BUFX4 port map( A => N188, Y => n27);
   U45 : BUFX4 port map( A => state_0_port, Y => n28);
   U46 : AND2X2 port map( A => state_2_port, B => n26, Y => n23);
   U47 : XOR2X1 port map( A => n22, B => n13, Y => n116);
   U48 : XOR2X1 port map( A => n25, B => n9, Y => n99);
   U49 : XOR2X1 port map( A => n24, B => n6, Y => n105);
   U50 : BUFX4 port map( A => state_1_port, Y => n26);
   U51 : INVX2 port map( A => n27, Y => n153);
   U52 : INVX2 port map( A => state_2_port, Y => n64_port);
   U53 : INVX2 port map( A => n26, Y => n30);
   U54 : NAND3X1 port map( A => n28, B => n64_port, C => n30, Y => n88);
   U55 : NAND3X1 port map( A => n26, B => n64_port, C => n36, Y => n93);
   U56 : NAND2X1 port map( A => n88, B => n93, Y => n69);
   U57 : NAND2X1 port map( A => n69, B => n29, Y => n56);
   U58 : NAND2X1 port map( A => state_2_port, B => n30, Y => n35);
   U59 : NOR2X1 port map( A => n36, B => n35, Y => n32);
   U60 : INVX2 port map( A => n222, Y => n31);
   U61 : NAND2X1 port map( A => n32, B => n31, Y => n33);
   U62 : OAI21X1 port map( A => n189, B => n56, C => n33, Y => n220);
   U63 : NAND2X1 port map( A => n23, B => n36, Y => n65_port);
   U64 : NAND2X1 port map( A => n34, B => n29, Y => n39);
   U65 : INVX2 port map( A => n35, Y => n68);
   U66 : NAND2X1 port map( A => n68, B => n36, Y => n127);
   U67 : NAND2X1 port map( A => n138, B => n29, Y => n38);
   U68 : INVX2 port map( A => t_crc(15), Y => n37);
   U69 : OAI22X1 port map( A => n188_port, B => n39, C => n38, D => n37, Y => 
                           n221);
   U70 : INVX2 port map( A => n38, Y => n53);
   U71 : INVX2 port map( A => n39, Y => n52);
   U72 : AOI22X1 port map( A => t_crc(14), B => n53, C => PRGA_OUT(6), D => n52
                           , Y => n225);
   U73 : INVX2 port map( A => flop_data_6_port, Y => n86);
   U74 : NAND3X1 port map( A => n245, B => n28, C => n68, Y => n55);
   U75 : INVX2 port map( A => t_crc(6), Y => n40);
   U76 : OAI22X1 port map( A => n56, B => n86, C => n55, D => n40, Y => n41);
   U77 : INVX2 port map( A => n41, Y => n226);
   U78 : AOI22X1 port map( A => t_crc(13), B => n53, C => PRGA_OUT(5), D => n52
                           , Y => n228);
   U79 : INVX2 port map( A => flop_data_5_port, Y => n84);
   U80 : INVX2 port map( A => t_crc(5), Y => n42);
   U81 : OAI22X1 port map( A => n56, B => n84, C => n55, D => n42, Y => n43);
   U82 : INVX2 port map( A => n43, Y => n229);
   U83 : AOI22X1 port map( A => t_crc(12), B => n53, C => PRGA_OUT(4), D => n52
                           , Y => n231);
   U84 : INVX2 port map( A => flop_data_4_port, Y => n82);
   U85 : INVX2 port map( A => t_crc(4), Y => n44);
   U86 : OAI22X1 port map( A => n56, B => n82, C => n55, D => n44, Y => n45);
   U87 : INVX2 port map( A => n45, Y => n232);
   U88 : AOI22X1 port map( A => t_crc(11), B => n53, C => PRGA_OUT(3), D => n52
                           , Y => n234);
   U89 : INVX2 port map( A => flop_data_3_port, Y => n80);
   U90 : INVX2 port map( A => t_crc(3), Y => n46);
   U91 : OAI22X1 port map( A => n56, B => n80, C => n55, D => n46, Y => n47);
   U92 : INVX2 port map( A => n47, Y => n235);
   U93 : AOI22X1 port map( A => t_crc(10), B => n53, C => PRGA_OUT(2), D => n52
                           , Y => n237);
   U94 : INVX2 port map( A => flop_data_2_port, Y => n78);
   U95 : INVX2 port map( A => t_crc(2), Y => n48);
   U96 : OAI22X1 port map( A => n56, B => n78, C => n55, D => n48, Y => n49);
   U97 : INVX2 port map( A => n49, Y => n238);
   U98 : AOI22X1 port map( A => t_crc(9), B => n53, C => PRGA_OUT(1), D => n52,
                           Y => n240);
   U99 : INVX2 port map( A => flop_data_1_port, Y => n76);
   U100 : INVX2 port map( A => t_crc(1), Y => n50);
   U101 : OAI22X1 port map( A => n56, B => n76, C => n55, D => n50, Y => n51);
   U102 : INVX2 port map( A => n51, Y => n241);
   U103 : AOI22X1 port map( A => t_crc(8), B => n53, C => PRGA_OUT(0), D => n52
                           , Y => n243);
   U104 : INVX2 port map( A => flop_data_0_port, Y => n74);
   U105 : INVX2 port map( A => t_crc(0), Y => n54);
   U106 : OAI22X1 port map( A => n56, B => n74, C => n55, D => n54, Y => n57);
   U107 : INVX2 port map( A => n57, Y => n244);
   U108 : INVX2 port map( A => count_4_port, Y => n155);
   U109 : INVX2 port map( A => count_5_port, Y => n154);
   U110 : INVX2 port map( A => n88, Y => n139);
   U111 : NAND2X1 port map( A => n157, B => n139, Y => n58);
   U112 : NOR2X1 port map( A => n156, B => n58, Y => t_strobe);
   U113 : NOR3X1 port map( A => n26, B => n28, C => state_2_port, Y => n131);
   U114 : INVX2 port map( A => p_ready, Y => n59_port);
   U115 : NAND2X1 port map( A => n131, B => n59_port, Y => n70);
   U116 : OAI21X1 port map( A => n187, B => n5, C => n70, Y => n60_port);
   U117 : AOI21X1 port map( A => n23, B => n28, C => n60_port, Y => n61_port);
   U118 : INVX2 port map( A => n61_port, Y => next_byte);
   U119 : NAND2X1 port map( A => n247, B => n27, Y => n63_port);
   U120 : NAND2X1 port map( A => n68, B => n62_port, Y => n141);
   U121 : OAI22X1 port map( A => n63_port, B => n141, C => n185, D => n93, Y =>
                           EOP);
   U122 : NAND2X1 port map( A => n68, B => n153, Y => n67);
   U123 : NAND3X1 port map( A => n28, B => n26, C => n64_port, Y => n92);
   U124 : NAND2X1 port map( A => n65_port, B => n92, Y => n142);
   U125 : NOR2X1 port map( A => n142, B => n69, Y => n66);
   U126 : NAND3X1 port map( A => n127, B => n66, C => n67, Y => sending);
   U127 : INVX2 port map( A => PRGA_OUT(0), Y => n73);
   U128 : NOR3X1 port map( A => n69, B => n23, C => n68, Y => n72);
   U129 : AND2X2 port map( A => n70, B => n29, Y => n71);
   U130 : AND2X2 port map( A => n72, B => n71, Y => n87);
   U131 : MUX2X1 port map( B => n74, A => n73, S => n87, Y => n260);
   U132 : INVX2 port map( A => PRGA_OUT(1), Y => n75);
   U133 : MUX2X1 port map( B => n76, A => n75, S => n87, Y => n259);
   U134 : INVX2 port map( A => PRGA_OUT(2), Y => n77);
   U135 : MUX2X1 port map( B => n78, A => n77, S => n87, Y => n258);
   U136 : INVX2 port map( A => PRGA_OUT(3), Y => n79);
   U137 : MUX2X1 port map( B => n80, A => n79, S => n87, Y => n257);
   U138 : INVX2 port map( A => PRGA_OUT(4), Y => n81);
   U139 : MUX2X1 port map( B => n82, A => n81, S => n87, Y => n256);
   U140 : INVX2 port map( A => PRGA_OUT(5), Y => n83);
   U141 : MUX2X1 port map( B => n84, A => n83, S => n87, Y => n255);
   U142 : INVX2 port map( A => PRGA_OUT(6), Y => n85);
   U143 : MUX2X1 port map( B => n86, A => n85, S => n87, Y => n254);
   U144 : MUX2X1 port map( B => n189, A => n188_port, S => n87, Y => n253);
   U145 : OAI21X1 port map( A => n186, B => n127, C => n88, Y => n89);
   U146 : NAND2X1 port map( A => t_bitstuff, B => n139, Y => n100);
   U147 : OAI21X1 port map( A => n90, B => n89, C => n100, Y => n91);
   U148 : INVX2 port map( A => n91, Y => n146);
   U149 : NAND2X1 port map( A => N63, B => n146, Y => n98);
   U150 : NAND2X1 port map( A => n9, B => n25, Y => n109);
   U151 : OR2X2 port map( A => n186, B => n92, Y => n132);
   U152 : NAND2X1 port map( A => n125, B => n140, Y => n94);
   U153 : NOR2X1 port map( A => n109, B => n10, Y => n96);
   U154 : NAND2X1 port map( A => n109, B => n147, Y => n95);
   U155 : NAND2X1 port map( A => n100, B => n95, Y => n111);
   U156 : MUX2X1 port map( B => n96, A => n111, S => n8, Y => n97);
   U157 : NAND2X1 port map( A => n98, B => n97, Y => n264);
   U158 : NAND2X1 port map( A => N62, B => n146, Y => n104);
   U159 : NAND2X1 port map( A => n99, B => n147, Y => n103);
   U160 : INVX2 port map( A => n100, Y => n150);
   U161 : INVX2 port map( A => n190, Y => n101);
   U162 : NAND2X1 port map( A => n150, B => n101, Y => n102);
   U163 : NAND3X1 port map( A => n104, B => n103, C => n102, Y => n265);
   U164 : NAND2X1 port map( A => N61, B => n146, Y => n108);
   U165 : NAND2X1 port map( A => n105, B => n147, Y => n107);
   U166 : NAND2X1 port map( A => n150, B => n6, Y => n106);
   U167 : NAND3X1 port map( A => n108, B => n107, C => n106, Y => n266);
   U168 : NAND2X1 port map( A => N64, B => n146, Y => n115);
   U169 : NAND3X1 port map( A => n110, B => n8, C => n147, Y => n119);
   U170 : INVX2 port map( A => n119, Y => n113);
   U171 : NAND2X1 port map( A => n147, B => n155, Y => n112);
   U172 : MUX2X1 port map( B => n113, A => n1, S => n7, Y => n114);
   U173 : NAND2X1 port map( A => n115, B => n114, Y => n263);
   U174 : AOI22X1 port map( A => n116, B => n147, C => N60, D => n146, Y => 
                           n118);
   U175 : NAND2X1 port map( A => n150, B => n13, Y => n117);
   U176 : NAND2X1 port map( A => n118, B => n117, Y => n267);
   U177 : NAND2X1 port map( A => N65, B => n146, Y => n124);
   U178 : NOR2X1 port map( A => n154, B => n119, Y => n122);
   U179 : NAND2X1 port map( A => n147, B => n154, Y => n120);
   U180 : NAND2X1 port map( A => n15, B => n14, Y => n121);
   U181 : MUX2X1 port map( B => n122, A => n121, S => n27, Y => n123);
   U182 : NAND2X1 port map( A => n124, B => n123, Y => n262);
   U183 : NAND2X1 port map( A => n177, B => p_ready, Y => n130);
   U184 : NAND2X1 port map( A => n126, B => n21, Y => n129);
   U185 : AND2X2 port map( A => n127, B => n141, Y => n128);
   U186 : NAND3X1 port map( A => n130, B => n129, C => n128, Y => 
                           nextstate_2_port);
   U187 : NAND2X1 port map( A => n131, B => p_ready, Y => n136);
   U188 : NAND2X1 port map( A => n21, B => n140, Y => n135);
   U189 : INVX2 port map( A => n132, Y => n133);
   U190 : AOI21X1 port map( A => n179, B => n139, C => n133, Y => n134);
   U191 : NAND3X1 port map( A => n136, B => n135, C => n134, Y => 
                           nextstate_1_port);
   U192 : AOI22X1 port map( A => n184, B => n139, C => n138, D => n137, Y => 
                           n145);
   U194 : NAND3X1 port map( A => n21, B => n140, C => p_ready, Y => n144);
   U196 : NOR2X1 port map( A => n142, B => n90, Y => n143);
   U198 : NAND3X1 port map( A => n145, B => n144, C => n143, Y => 
                           nextstate_0_port);
   U203 : XOR2X1 port map( A => n175, B => t_bitstuff, Y => n148);
   U204 : AOI22X1 port map( A => n148, B => n147, C => N59, D => n146, Y => 
                           n152);
   U205 : INVX2 port map( A => n175, Y => n149);
   U206 : NAND2X1 port map( A => n150, B => n149, Y => n151);
   U207 : NAND2X1 port map( A => n152, B => n151, Y => n261);
   U208 : NAND2X1 port map( A => n153, B => n175, Y => n156);
   U209 : NOR2X1 port map( A => n26, B => n28, Y => n177);
   U210 : INVX1 port map( A => n184, Y => n179);
   U211 : NAND3X1 port map( A => n157, B => n153, C => count_0_port, Y => n184)
                           ;
   U212 : AND2X1 port map( A => prga_opcode(1), B => prga_opcode(0), Y => n187)
                           ;
   U213 : NAND3X1 port map( A => n8, B => n13, C => n7, Y => n193);
   U214 : NOR2X1 port map( A => n27, B => n191, Y => n201);
   U215 : OAI21X1 port map( A => n202, B => n203, C => n204, Y => n275);
   U216 : INVX1 port map( A => current_send_data_7_port, Y => n203);
   U217 : OAI21X1 port map( A => n202, B => n205, C => n206, Y => n276);
   U218 : INVX1 port map( A => current_send_data_6_port, Y => n205);
   U219 : OAI21X1 port map( A => n202, B => n207, C => n208, Y => n277);
   U220 : INVX1 port map( A => current_send_data_5_port, Y => n207);
   U221 : OAI21X1 port map( A => n202, B => n209, C => n210, Y => n278);
   U222 : INVX1 port map( A => current_send_data_4_port, Y => n209);
   U223 : OAI21X1 port map( A => n202, B => n211, C => n212, Y => n279);
   U224 : INVX1 port map( A => current_send_data_3_port, Y => n211);
   U225 : OAI21X1 port map( A => n202, B => n213, C => n214, Y => n280);
   U226 : INVX1 port map( A => current_send_data_2_port, Y => n213);
   U227 : OAI21X1 port map( A => n202, B => n215, C => n216, Y => n281);
   U228 : INVX1 port map( A => current_send_data_1_port, Y => n215);
   U229 : OAI21X1 port map( A => n202, B => n217, C => n218, Y => n282);
   U230 : INVX1 port map( A => current_send_data_0_port, Y => n217);
   U231 : AOI21X1 port map( A => n28, B => n26, C => rst, Y => n202);
   U232 : NAND2X1 port map( A => n219, B => n204, Y => n283);
   U233 : NOR2X1 port map( A => n220, B => n221, Y => n204);
   U234 : INVX1 port map( A => PRGA_OUT(7), Y => n188_port);
   U235 : OAI21X1 port map( A => n27, B => t_crc(7), C => n29, Y => n222);
   U236 : INVX1 port map( A => flop_data_7_port, Y => n189);
   U237 : AOI22X1 port map( A => n223, B => current_send_data_7_port, C => 
                           send_data_7_port, D => rst, Y => n219);
   U238 : NAND2X1 port map( A => n224, B => n206, Y => n284);
   U239 : AND2X1 port map( A => n225, B => n226, Y => n206);
   U240 : AOI22X1 port map( A => n223, B => current_send_data_6_port, C => 
                           send_data_6_port, D => rst, Y => n224);
   U241 : NAND2X1 port map( A => n227, B => n208, Y => n285);
   U242 : AND2X1 port map( A => n228, B => n229, Y => n208);
   U243 : AOI22X1 port map( A => n223, B => current_send_data_5_port, C => 
                           send_data_5_port, D => rst, Y => n227);
   U244 : NAND2X1 port map( A => n230, B => n210, Y => n286);
   U245 : AND2X1 port map( A => n231, B => n232, Y => n210);
   U246 : AOI22X1 port map( A => n223, B => current_send_data_4_port, C => 
                           send_data_4_port, D => rst, Y => n230);
   U247 : NAND2X1 port map( A => n233, B => n212, Y => n287);
   U248 : AND2X1 port map( A => n234, B => n235, Y => n212);
   U249 : AOI22X1 port map( A => n223, B => current_send_data_3_port, C => 
                           send_data_3_port, D => rst, Y => n233);
   U250 : NAND2X1 port map( A => n236, B => n214, Y => n288);
   U251 : AND2X1 port map( A => n237, B => n238, Y => n214);
   U252 : AOI22X1 port map( A => n223, B => current_send_data_2_port, C => 
                           send_data_2_port, D => rst, Y => n236);
   U253 : NAND2X1 port map( A => n239, B => n216, Y => n289);
   U254 : AND2X1 port map( A => n240, B => n241, Y => n216);
   U255 : AOI22X1 port map( A => n223, B => current_send_data_1_port, C => 
                           send_data_1_port, D => rst, Y => n239);
   U256 : NAND2X1 port map( A => n242, B => n218, Y => n290);
   U257 : AND2X1 port map( A => n243, B => n244, Y => n218);
   U258 : NOR2X1 port map( A => rst, B => n27, Y => n245);
   U259 : AOI22X1 port map( A => n223, B => current_send_data_0_port, C => 
                           send_data_0_port, D => rst, Y => n242);
   U260 : INVX1 port map( A => n246, Y => n223);
   U261 : NAND3X1 port map( A => n28, B => n29, C => n26, Y => n246);
   U262 : OAI21X1 port map( A => n249, B => n250, C => n28, Y => n248);
   U263 : NAND3X1 port map( A => count_2_port, B => n27, C => n9, Y => n250);
   U264 : NAND3X1 port map( A => n155, B => n154, C => n251, Y => n249);
   U265 : NOR2X1 port map( A => n12, B => count_0_port, Y => n251);
   U266 : NAND3X1 port map( A => n157, B => n175, C => n27, Y => n185);
   U267 : NOR2X1 port map( A => n247, B => n13, Y => n157);
   U268 : NAND3X1 port map( A => n191, B => n190, C => n252, Y => n247);
   U269 : NOR2X1 port map( A => count_5_port, B => count_4_port, Y => n252);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_shiftreg_0 is

   port( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe : in std_logic;  
         send_data : in std_logic_vector (7 downto 0);  d_encode : out 
         std_logic);

end tx_shiftreg_0;

architecture SYN_dataflow of tx_shiftreg_0 is

   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal d_encode_port, present_val_7_port, present_val_6_port, 
      present_val_5_port, present_val_4_port, present_val_3_port, 
      present_val_2_port, present_val_1_port, count_2_port, count_1_port, 
      count_0_port, n1, n2, n3, n4, n5, n6, n7, n11, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83 : std_logic;

begin
   d_encode <= d_encode_port;
   
   count_reg_0_inst : DFFSR port map( D => n69, CLK => clk, R => n80, S => n17,
                           Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => n71, CLK => clk, R => n81, S => n17,
                           Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n70, CLK => clk, R => n82, S => n17,
                           Q => count_2_port);
   present_val_reg_7_inst : DFFSR port map( D => n78, CLK => clk, R => n17, S 
                           => n83, Q => present_val_7_port);
   n83 <= '1';
   n82 <= '1';
   n81 <= '1';
   n80 <= '1';
   present_val_reg_6_inst : DFFSR port map( D => n77, CLK => clk, R => n17, S 
                           => n11, Q => present_val_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n76, CLK => clk, R => n17, S 
                           => n7, Q => present_val_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n75, CLK => clk, R => n17, S 
                           => n6, Q => present_val_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n74, CLK => clk, R => n17, S 
                           => n5, Q => present_val_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n73, CLK => clk, R => n17, S 
                           => n4, Q => present_val_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n72, CLK => clk, R => n17, S 
                           => n3, Q => present_val_1_port);
   present_val_reg_0_inst : DFFSR port map( D => n79, CLK => clk, R => n17, S 
                           => n2, Q => d_encode_port);
   U3 : AND2X2 port map( A => n19, B => count_2_port, Y => n1);
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n11 <= '1';
   U15 : INVX2 port map( A => n20, Y => n13);
   U16 : OR2X2 port map( A => n13, B => n15, Y => n67);
   U17 : INVX2 port map( A => n15, Y => n16);
   U18 : INVX1 port map( A => t_bitstuff, Y => n18);
   U19 : AND2X2 port map( A => n67, B => n16, Y => n14);
   U20 : INVX2 port map( A => n14, Y => n68);
   U21 : AND2X2 port map( A => n1, B => SHIFT_ENABLE_R, Y => n15);
   U22 : INVX2 port map( A => rst, Y => n17);
   U23 : INVX1 port map( A => n67, Y => n56);
   U24 : NAND2X1 port map( A => SHIFT_ENABLE_R, B => n18, Y => n20);
   U25 : NAND2X1 port map( A => count_1_port, B => count_0_port, Y => n64);
   U26 : INVX2 port map( A => n64, Y => n19);
   U27 : NAND2X1 port map( A => d_encode_port, B => n56, Y => n24);
   U28 : NAND2X1 port map( A => present_val_1_port, B => n14, Y => n23);
   U29 : INVX2 port map( A => send_data(0), Y => n21);
   U30 : OR2X2 port map( A => n16, B => n21, Y => n22);
   U31 : NAND3X1 port map( A => n24, B => n23, C => n22, Y => n79);
   U32 : NAND2X1 port map( A => present_val_1_port, B => n56, Y => n28);
   U33 : NAND2X1 port map( A => present_val_2_port, B => n14, Y => n27);
   U34 : INVX2 port map( A => send_data(1), Y => n25);
   U35 : OR2X2 port map( A => n16, B => n25, Y => n26);
   U36 : NAND3X1 port map( A => n28, B => n27, C => n26, Y => n72);
   U37 : NAND2X1 port map( A => present_val_2_port, B => n56, Y => n32);
   U38 : NAND2X1 port map( A => present_val_3_port, B => n14, Y => n31);
   U39 : INVX2 port map( A => send_data(2), Y => n29);
   U40 : OR2X2 port map( A => n16, B => n29, Y => n30);
   U41 : NAND3X1 port map( A => n32, B => n31, C => n30, Y => n73);
   U42 : NAND2X1 port map( A => present_val_3_port, B => n56, Y => n36);
   U43 : NAND2X1 port map( A => present_val_4_port, B => n14, Y => n35);
   U44 : INVX2 port map( A => send_data(3), Y => n33);
   U45 : OR2X2 port map( A => n16, B => n33, Y => n34);
   U46 : NAND3X1 port map( A => n36, B => n35, C => n34, Y => n74);
   U47 : NAND2X1 port map( A => present_val_4_port, B => n56, Y => n40);
   U48 : NAND2X1 port map( A => present_val_5_port, B => n14, Y => n39);
   U49 : INVX2 port map( A => send_data(4), Y => n37);
   U50 : OR2X2 port map( A => n16, B => n37, Y => n38);
   U51 : NAND3X1 port map( A => n40, B => n39, C => n38, Y => n75);
   U52 : NAND2X1 port map( A => present_val_5_port, B => n56, Y => n55);
   U53 : NAND2X1 port map( A => present_val_6_port, B => n14, Y => n54);
   U54 : INVX2 port map( A => send_data(5), Y => n41);
   U55 : OR2X2 port map( A => n16, B => n41, Y => n42);
   U56 : NAND3X1 port map( A => n55, B => n54, C => n42, Y => n76);
   U57 : NAND2X1 port map( A => present_val_6_port, B => n56, Y => n60);
   U58 : NAND2X1 port map( A => present_val_7_port, B => n14, Y => n59);
   U59 : INVX2 port map( A => send_data(6), Y => n57);
   U60 : OR2X2 port map( A => n16, B => n57, Y => n58);
   U61 : NAND3X1 port map( A => n60, B => n59, C => n58, Y => n77);
   U62 : INVX2 port map( A => present_val_7_port, Y => n62);
   U63 : INVX2 port map( A => send_data(7), Y => n61);
   U64 : OAI22X1 port map( A => n67, B => n62, C => n16, D => n61, Y => n78);
   U65 : NAND2X1 port map( A => count_2_port, B => n16, Y => n63);
   U66 : OAI21X1 port map( A => n64, B => n68, C => n63, Y => n70);
   U67 : NAND2X1 port map( A => n14, B => count_0_port, Y => n66);
   U68 : AND2X2 port map( A => count_0_port, B => n67, Y => n65);
   U69 : MUX2X1 port map( B => n66, A => n65, S => count_1_port, Y => n71);
   U70 : MUX2X1 port map( B => n68, A => n67, S => count_0_port, Y => n69);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_encode_0 is

   port( clk, rst, SHIFT_ENABLE_E, d_encode, EOP : in std_logic;  t_bitstuff, 
         dp_tx_out, dm_tx_out : out std_logic);

end tx_encode_0;

architecture SYN_moore of tx_encode_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal DE_holdout, DE_holdout_BS, state_3_port, state_2_port, state_1_port, 
      state_0_port, nextstate_3_port, nextstate_2_port, nextstate_1_port, 
      nextstate_0_port, DE_holdout_last, DE_holdout_nxt, dm_tx_nxt, n1, n2, n3,
      n5, n6, n7, n8, n10, n11, n16, n17, n21, n22, n23, n24, n25, n28, n29, 
      n30, n31, n33, n34, n35, n36, n38, n42, n45, n46, n47, n48, n51, n52, n53
      , n56, n57, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97 : std_logic;

begin
   
   DE_holdout_reg : DFFSR port map( D => DE_holdout_nxt, CLK => clk, R => n72, 
                           S => n11, Q => DE_holdout);
   DE_holdout_last_reg : DFFPOSX1 port map( D => n73, CLK => clk, Q => 
                           DE_holdout_last);
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => clk, R => 
                           n11, S => n74, Q => state_3_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n11, S => n75, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n11, S => n76, Q => state_1_port);
   dp_tx_out_reg : DFFSR port map( D => DE_holdout_nxt, CLK => clk, R => n77, S
                           => n11, Q => dp_tx_out);
   dm_tx_out_reg : DFFSR port map( D => dm_tx_nxt, CLK => clk, R => n11, S => 
                           n78, Q => dm_tx_out);
   U9 : OAI21X1 port map( A => n3, B => n7, C => n95, Y => nextstate_1_port);
   U11 : OAI21X1 port map( A => n6, B => n8, C => n53, Y => n94);
   U12 : NAND3X1 port map( A => SHIFT_ENABLE_E, B => n65, C => n6, Y => n97);
   U14 : OAI21X1 port map( A => n5, B => n53, C => n92, Y => nextstate_0_port);
   U15 : OAI21X1 port map( A => n91, B => n90, C => SHIFT_ENABLE_E, Y => n92);
   U18 : NOR2X1 port map( A => n6, B => n93, Y => n91);
   U19 : NAND3X1 port map( A => d_encode, B => n89, C => n88, Y => n93);
   U20 : XNOR2X1 port map( A => n68, B => n67, Y => n88);
   U22 : NOR2X1 port map( A => n63, B => SHIFT_ENABLE_E, Y => n96);
   U23 : OAI22X1 port map( A => n11, B => n68, C => rst, D => n67, Y => n73);
   U26 : OAI22X1 port map( A => n10, B => n69, C => n67, D => n87, Y => n71);
   U36 : NOR2X1 port map( A => EOP, B => state_3_port, Y => n89);
   U37 : NOR2X1 port map( A => EOP, B => n84, Y => n86);
   U38 : AOI22X1 port map( A => n6, B => n83, C => n56, D => n5, Y => n84);
   U40 : XNOR2X1 port map( A => DE_holdout_BS, B => n81, Y => n83);
   U46 : XOR2X1 port map( A => DE_holdout, B => SHIFT_ENABLE_E, Y => n82);
   U47 : XNOR2X1 port map( A => n80, B => n67, Y => n85);
   U49 : NAND2X1 port map( A => SHIFT_ENABLE_E, B => n66, Y => n80);
   U55 : NAND2X1 port map( A => n81, B => n69, Y => n79);
   U57 : NAND2X1 port map( A => SHIFT_ENABLE_E, B => d_encode, Y => n81);
   n78 <= '1';
   n77 <= '1';
   n76 <= '1';
   n75 <= '1';
   n74 <= '1';
   n72 <= '1';
   DE_holdout_BS_reg : DFFSR port map( D => n71, CLK => clk, R => n11, S => n2,
                           Q => DE_holdout_BS);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n11, S => n1, Q => state_2_port);
   U3 : INVX2 port map( A => n38, Y => n3);
   U4 : INVX2 port map( A => state_0_port, Y => n5);
   U5 : INVX2 port map( A => n5, Y => n6);
   U6 : INVX1 port map( A => state_1_port, Y => n38);
   n1 <= '1';
   n2 <= '1';
   U10 : BUFX4 port map( A => n70, Y => t_bitstuff);
   U13 : INVX1 port map( A => n89, Y => n63);
   U16 : INVX1 port map( A => n52, Y => n7);
   U17 : INVX1 port map( A => n65, Y => n8);
   U21 : INVX2 port map( A => rst, Y => n11);
   U24 : NOR2X1 port map( A => n48, B => n17, Y => n10);
   U25 : INVX1 port map( A => n10, Y => n87);
   U27 : NAND2X1 port map( A => state_2_port, B => state_1_port, Y => n16);
   U28 : NOR3X1 port map( A => state_3_port, B => n16, C => n5, Y => n70);
   U29 : INVX2 port map( A => n16, Y => n31);
   U30 : NAND3X1 port map( A => n89, B => n5, C => n31, Y => n48);
   U31 : INVX2 port map( A => SHIFT_ENABLE_E, Y => n17);
   U32 : NAND2X1 port map( A => n66, B => n31, Y => n21);
   U33 : OAI21X1 port map( A => n63, B => n21, C => n48, Y => n90);
   U34 : INVX2 port map( A => n48, Y => n22);
   U35 : AOI21X1 port map( A => n94, B => n3, C => n22, Y => n95);
   U39 : INVX2 port map( A => state_2_port, Y => n23);
   U41 : NAND3X1 port map( A => n5, B => n23, C => n38, Y => n51);
   U42 : NAND2X1 port map( A => n51, B => state_3_port, Y => n36);
   U43 : INVX2 port map( A => n85, Y => n24);
   U44 : NOR2X1 port map( A => n63, B => n24, Y => n25);
   U45 : MUX2X1 port map( B => n25, A => n86, S => n31, Y => n28);
   U48 : NAND2X1 port map( A => n36, B => n28, Y => dm_tx_nxt);
   U50 : OAI21X1 port map( A => n69, B => n81, C => n79, Y => n30);
   U51 : AND2X2 port map( A => n82, B => n5, Y => n29);
   U52 : AOI21X1 port map( A => n6, B => n30, C => n29, Y => n33);
   U53 : MUX2X1 port map( B => n85, A => n33, S => n31, Y => n34);
   U54 : OAI21X1 port map( A => state_3_port, B => n34, C => n57, Y => n35);
   U56 : NAND2X1 port map( A => n36, B => n35, Y => DE_holdout_nxt);
   U58 : NAND2X1 port map( A => n52, B => n3, Y => n45);
   U59 : AOI21X1 port map( A => n65, B => n38, C => n96, Y => n42);
   U60 : MUX2X1 port map( B => n45, A => n42, S => state_2_port, Y => n46);
   U61 : INVX2 port map( A => n46, Y => n47);
   U62 : NAND2X1 port map( A => n48, B => n47, Y => nextstate_2_port);
   U63 : AOI21X1 port map( A => state_3_port, B => n51, C => n57, Y => 
                           nextstate_3_port);
   U64 : INVX2 port map( A => n97, Y => n52);
   U65 : INVX2 port map( A => n96, Y => n53);
   U68 : INVX2 port map( A => n82, Y => n56);
   U69 : INVX2 port map( A => EOP, Y => n57);
   U74 : INVX2 port map( A => n93, Y => n65);
   U75 : INVX2 port map( A => d_encode, Y => n66);
   U76 : INVX2 port map( A => DE_holdout, Y => n67);
   U77 : INVX2 port map( A => DE_holdout_last, Y => n68);
   U78 : INVX2 port map( A => DE_holdout_BS, Y => n69);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_CRC_CALC_0 is

   port( CLK, RST, EOP, T_STROBE : in std_logic;  PRGA_OPCODE : in 
         std_logic_vector (1 downto 0);  PRGA_OUT : in std_logic_vector (7 
         downto 0);  TX_CRC : out std_logic_vector (15 downto 0));

end tx_CRC_CALC_0;

architecture SYN_txcrcm of tx_CRC_CALC_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal TX_CRC_15_port, TX_CRC_14_port, TX_CRC_13_port, TX_CRC_12_port, 
      TX_CRC_11_port, TX_CRC_10_port, TX_CRC_9_port, TX_CRC_8_port, 
      TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port, TX_CRC_4_port, TX_CRC_3_port
      , TX_CRC_2_port, TX_CRC_1_port, TX_CRC_0_port, n1, n2, n3, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22
      , n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
      n37, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121 : std_logic;

begin
   TX_CRC <= ( TX_CRC_15_port, TX_CRC_14_port, TX_CRC_13_port, TX_CRC_12_port, 
      TX_CRC_11_port, TX_CRC_10_port, TX_CRC_9_port, TX_CRC_8_port, 
      TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port, TX_CRC_4_port, TX_CRC_3_port
      , TX_CRC_2_port, TX_CRC_1_port, TX_CRC_0_port );
   
   U39 : OAI22X1 port map( A => n25, B => n20, C => n121, D => n19, Y => n96);
   U40 : XNOR2X1 port map( A => n119, B => n79, Y => n121);
   U41 : OAI22X1 port map( A => n37, B => n20, C => n19, D => n36, Y => n95);
   U42 : OAI22X1 port map( A => n35, B => n20, C => n19, D => n34, Y => n94);
   U43 : OAI22X1 port map( A => n33, B => n20, C => n19, D => n32, Y => n93);
   U44 : OAI22X1 port map( A => n31, B => n20, C => n19, D => n30, Y => n92);
   U45 : OAI22X1 port map( A => n29, B => n20, C => n19, D => n28, Y => n91);
   U46 : OAI22X1 port map( A => n27, B => n20, C => n118, D => n19, Y => n90);
   U47 : XNOR2X1 port map( A => TX_CRC_1_port, B => n117, Y => n118);
   U48 : OAI22X1 port map( A => n24, B => n20, C => n116, D => n19, Y => n89);
   U49 : XOR2X1 port map( A => n115, B => n114, Y => n116);
   U50 : XNOR2X1 port map( A => TX_CRC_0_port, B => n117, Y => n115);
   U51 : OAI22X1 port map( A => n79, B => n20, C => n113, D => n19, Y => n88);
   U52 : OAI22X1 port map( A => n20, B => n36, C => n112, D => n19, Y => n87);
   U53 : XNOR2X1 port map( A => n111, B => n110, Y => n112);
   U54 : OAI22X1 port map( A => n20, B => n34, C => n109, D => n19, Y => n86);
   U55 : OAI22X1 port map( A => n20, B => n32, C => n108, D => n19, Y => n85);
   U56 : XNOR2X1 port map( A => n107, B => n106, Y => n108);
   U57 : OAI22X1 port map( A => n20, B => n30, C => n105, D => n19, Y => n84);
   U58 : OAI22X1 port map( A => n20, B => n28, C => n104, D => n19, Y => n83);
   U59 : XOR2X1 port map( A => n103, B => n102, Y => n104);
   U60 : OAI22X1 port map( A => n20, B => n26, C => n101, D => n19, Y => n82);
   U61 : XOR2X1 port map( A => n100, B => n99, Y => n101);
   U62 : XOR2X1 port map( A => n117, B => n113, Y => n100);
   U63 : OAI22X1 port map( A => n20, B => n23, C => n119, D => n19, Y => n81);
   U64 : XOR2X1 port map( A => n98, B => n97, Y => n119);
   U65 : XOR2X1 port map( A => n102, B => n117, Y => n97);
   U66 : XNOR2X1 port map( A => n25, B => PRGA_OUT(7), Y => n117);
   U67 : XNOR2X1 port map( A => n24, B => PRGA_OUT(0), Y => n102);
   U68 : XOR2X1 port map( A => n113, B => n99, Y => n98);
   U69 : XOR2X1 port map( A => n105, B => n109, Y => n99);
   U70 : XNOR2X1 port map( A => n106, B => n111, Y => n109);
   U71 : XOR2X1 port map( A => TX_CRC_12_port, B => PRGA_OUT(4), Y => n111);
   U72 : XOR2X1 port map( A => TX_CRC_11_port, B => PRGA_OUT(3), Y => n106);
   U74 : XOR2X1 port map( A => TX_CRC_10_port, B => PRGA_OUT(2), Y => n107);
   U75 : XNOR2X1 port map( A => TX_CRC_9_port, B => PRGA_OUT(1), Y => n103);
   U76 : XNOR2X1 port map( A => n110, B => n114, Y => n113);
   U77 : XNOR2X1 port map( A => n37, B => PRGA_OUT(6), Y => n114);
   U78 : XOR2X1 port map( A => TX_CRC_13_port, B => PRGA_OUT(5), Y => n110);
   U80 : NAND3X1 port map( A => PRGA_OPCODE(0), B => n80, C => T_STROBE, Y => 
                           n120);
   current_crc_reg_6_inst : DFFSR port map( D => n87, CLK => CLK, R => n21, S 
                           => n16, Q => TX_CRC_6_port);
   current_crc_reg_5_inst : DFFSR port map( D => n86, CLK => CLK, R => n21, S 
                           => n15, Q => TX_CRC_5_port);
   current_crc_reg_4_inst : DFFSR port map( D => n85, CLK => CLK, R => n21, S 
                           => n14, Q => TX_CRC_4_port);
   current_crc_reg_3_inst : DFFSR port map( D => n84, CLK => CLK, R => n21, S 
                           => n13, Q => TX_CRC_3_port);
   current_crc_reg_2_inst : DFFSR port map( D => n83, CLK => CLK, R => n21, S 
                           => n12, Q => TX_CRC_2_port);
   current_crc_reg_1_inst : DFFSR port map( D => n82, CLK => CLK, R => n21, S 
                           => n11, Q => TX_CRC_1_port);
   current_crc_reg_0_inst : DFFSR port map( D => n81, CLK => CLK, R => n21, S 
                           => n10, Q => TX_CRC_0_port);
   current_crc_reg_15_inst : DFFSR port map( D => n96, CLK => CLK, R => n21, S 
                           => n9, Q => TX_CRC_15_port);
   current_crc_reg_9_inst : DFFSR port map( D => n90, CLK => CLK, R => n21, S 
                           => n8, Q => TX_CRC_9_port);
   current_crc_reg_8_inst : DFFSR port map( D => n89, CLK => CLK, R => n21, S 
                           => n7, Q => TX_CRC_8_port);
   current_crc_reg_14_inst : DFFSR port map( D => n95, CLK => CLK, R => n21, S 
                           => n6, Q => TX_CRC_14_port);
   current_crc_reg_13_inst : DFFSR port map( D => n94, CLK => CLK, R => n21, S 
                           => n5, Q => TX_CRC_13_port);
   current_crc_reg_12_inst : DFFSR port map( D => n93, CLK => CLK, R => n21, S 
                           => n4, Q => TX_CRC_12_port);
   current_crc_reg_11_inst : DFFSR port map( D => n92, CLK => CLK, R => n21, S 
                           => n3, Q => TX_CRC_11_port);
   current_crc_reg_10_inst : DFFSR port map( D => n91, CLK => CLK, R => n21, S 
                           => n2, Q => TX_CRC_10_port);
   current_crc_reg_7_inst : DFFSR port map( D => n88, CLK => CLK, R => n21, S 
                           => n1, Q => TX_CRC_7_port);
   U3 : INVX2 port map( A => n17, Y => n20);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   U20 : INVX1 port map( A => EOP, Y => n22);
   U21 : INVX2 port map( A => n120, Y => n18);
   U22 : AND2X2 port map( A => n120, B => n22, Y => n17);
   U23 : INVX2 port map( A => RST, Y => n21);
   U24 : XOR2X1 port map( A => n103, B => n107, Y => n105);
   U25 : INVX2 port map( A => n18, Y => n19);
   U26 : INVX2 port map( A => TX_CRC_0_port, Y => n23);
   U27 : INVX2 port map( A => TX_CRC_8_port, Y => n24);
   U28 : INVX2 port map( A => TX_CRC_15_port, Y => n25);
   U29 : INVX2 port map( A => TX_CRC_1_port, Y => n26);
   U30 : INVX2 port map( A => TX_CRC_9_port, Y => n27);
   U31 : INVX2 port map( A => TX_CRC_2_port, Y => n28);
   U32 : INVX2 port map( A => TX_CRC_10_port, Y => n29);
   U33 : INVX2 port map( A => TX_CRC_3_port, Y => n30);
   U34 : INVX2 port map( A => TX_CRC_11_port, Y => n31);
   U35 : INVX2 port map( A => TX_CRC_4_port, Y => n32);
   U36 : INVX2 port map( A => TX_CRC_12_port, Y => n33);
   U37 : INVX2 port map( A => TX_CRC_5_port, Y => n34);
   U38 : INVX2 port map( A => TX_CRC_13_port, Y => n35);
   U73 : INVX2 port map( A => TX_CRC_6_port, Y => n36);
   U79 : INVX2 port map( A => TX_CRC_14_port, Y => n37);
   U81 : INVX2 port map( A => TX_CRC_7_port, Y => n79);
   U82 : INVX2 port map( A => PRGA_OPCODE(1), Y => n80);

end SYN_txcrcm;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_timer_0 is

   port( CLK, RST, D_EDGE, RCVING : in std_logic;  SHIFT_ENABLE : out std_logic
         );

end rx_timer_0;

architecture SYN_moore of rx_timer_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal count_3_port, count_2_port, count_1_port, count_0_port, state, 
      nextcount_3_port, nextcount_2_port, nextcount_1_port, nextcount_0_port, 
      n5, n7, n9, n10, n11, n12, n13, n14, n16, n19, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41 : 
      std_logic;

begin
   
   state_reg : DFFSR port map( D => n7, CLK => CLK, R => n12, S => n37, Q => 
                           state);
   count_reg_0_inst : DFFSR port map( D => nextcount_0_port, CLK => CLK, R => 
                           n12, S => n38, Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => nextcount_1_port, CLK => CLK, R => 
                           n12, S => n39, Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => nextcount_2_port, CLK => CLK, R => 
                           n12, S => n40, Q => count_2_port);
   count_reg_3_inst : DFFSR port map( D => nextcount_3_port, CLK => CLK, R => 
                           n12, S => n41, Q => count_3_port);
   n41 <= '1';
   n40 <= '1';
   n39 <= '1';
   n38 <= '1';
   n37 <= '1';
   U19 : XOR2X1 port map( A => n34, B => n27, Y => n35);
   U20 : NOR2X1 port map( A => count_3_port, B => n28, Y => n36);
   U22 : XOR2X1 port map( A => n32, B => count_2_port, Y => n33);
   U24 : NAND2X1 port map( A => state, B => n30, Y => nextcount_0_port);
   U25 : OAI21X1 port map( A => D_EDGE, B => n29, C => n7, Y => n30);
   U30 : NAND2X1 port map( A => count_0_port, B => count_1_port, Y => n32);
   U32 : XNOR2X1 port map( A => count_0_port, B => count_1_port, Y => n31);
   U7 : INVX1 port map( A => RCVING, Y => n5);
   U9 : INVX2 port map( A => n5, Y => n7);
   U10 : NOR2X1 port map( A => n24, B => n19, Y => SHIFT_ENABLE);
   U11 : INVX2 port map( A => n9, Y => nextcount_2_port);
   U12 : INVX2 port map( A => RST, Y => n12);
   U13 : OAI21X1 port map( A => n10, B => D_EDGE, C => n7, Y => n9);
   U14 : NAND2X1 port map( A => n33, B => state, Y => n10);
   U15 : NOR2X1 port map( A => D_EDGE, B => n16, Y => n11);
   U16 : INVX2 port map( A => count_2_port, Y => n13);
   U17 : OAI21X1 port map( A => n31, B => n13, C => n32, Y => n34);
   U18 : XOR2X1 port map( A => n13, B => n31, Y => n27);
   U21 : INVX2 port map( A => n27, Y => n14);
   U23 : NAND2X1 port map( A => RCVING, B => n14, Y => n24);
   U26 : INVX2 port map( A => state, Y => n16);
   U27 : INVX2 port map( A => n34, Y => n28);
   U28 : NAND3X1 port map( A => count_3_port, B => n11, C => n28, Y => n19);
   U29 : AOI22X1 port map( A => n36, B => n27, C => n35, D => count_3_port, Y 
                           => n25);
   U31 : NAND2X1 port map( A => n7, B => n11, Y => n26);
   U33 : NOR2X1 port map( A => n25, B => n26, Y => nextcount_3_port);
   U34 : NOR2X1 port map( A => n31, B => n26, Y => nextcount_1_port);
   U35 : INVX2 port map( A => count_0_port, Y => n29);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_shift_reg_0 is

   port( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF : in std_logic;  RCV_DATA : 
         out std_logic_vector (7 downto 0));

end rx_shift_reg_0;

architecture SYN_dataflow of rx_shift_reg_0 is

   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      present_val_7_port, present_val_6_port, present_val_5_port, 
      present_val_4_port, present_val_3_port, present_val_2_port, 
      present_val_1_port, present_val_0_port, n1, n3, n4, n5, n7, n9, n11, n13,
      n15, n17, n19, n20, n22, n25, n28, n31, n34, n37, n40, n43, n45, n46, n47
      , n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   RCV_DATA_reg_7_inst : DFFPOSX1 port map( D => n49, CLK => CLK, Q => 
                           RCV_DATA_7_port);
   RCV_DATA_reg_6_inst : DFFPOSX1 port map( D => n51, CLK => CLK, Q => 
                           RCV_DATA_6_port);
   RCV_DATA_reg_5_inst : DFFPOSX1 port map( D => n53, CLK => CLK, Q => 
                           RCV_DATA_5_port);
   RCV_DATA_reg_4_inst : DFFPOSX1 port map( D => n55, CLK => CLK, Q => 
                           RCV_DATA_4_port);
   RCV_DATA_reg_3_inst : DFFPOSX1 port map( D => n57, CLK => CLK, Q => 
                           RCV_DATA_3_port);
   RCV_DATA_reg_2_inst : DFFPOSX1 port map( D => n59, CLK => CLK, Q => 
                           RCV_DATA_2_port);
   RCV_DATA_reg_1_inst : DFFPOSX1 port map( D => n61, CLK => CLK, Q => 
                           RCV_DATA_1_port);
   RCV_DATA_reg_0_inst : DFFPOSX1 port map( D => n63, CLK => CLK, Q => 
                           RCV_DATA_0_port);
   U2 : OAI21X1 port map( A => RST, B => n47, C => n71, Y => n63);
   U3 : NAND2X1 port map( A => RCV_DATA_0_port, B => RST, Y => n71);
   U6 : OAI21X1 port map( A => RST, B => n46, C => n70, Y => n61);
   U7 : NAND2X1 port map( A => RCV_DATA_1_port, B => RST, Y => n70);
   U10 : OAI21X1 port map( A => RST, B => n45, C => n69, Y => n59);
   U11 : NAND2X1 port map( A => RCV_DATA_2_port, B => RST, Y => n69);
   U14 : OAI21X1 port map( A => RST, B => n43, C => n68, Y => n57);
   U15 : NAND2X1 port map( A => RCV_DATA_3_port, B => RST, Y => n68);
   U18 : OAI21X1 port map( A => RST, B => n40, C => n67, Y => n55);
   U19 : NAND2X1 port map( A => RCV_DATA_4_port, B => RST, Y => n67);
   U22 : OAI21X1 port map( A => RST, B => n37, C => n66, Y => n53);
   U23 : NAND2X1 port map( A => RCV_DATA_5_port, B => RST, Y => n66);
   U26 : OAI21X1 port map( A => RST, B => n34, C => n65, Y => n51);
   U27 : NAND2X1 port map( A => n1, B => RST, Y => n65);
   U30 : OAI21X1 port map( A => RST, B => n31, C => n64, Y => n49);
   U31 : NAND2X1 port map( A => n19, B => RST, Y => n64);
   present_val_reg_0_inst : DFFSR port map( D => n62, CLK => CLK, R => n22, S 
                           => n15, Q => present_val_0_port);
   present_val_reg_7_inst : DFFSR port map( D => n48, CLK => CLK, R => n22, S 
                           => n13, Q => present_val_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n50, CLK => CLK, R => n22, S 
                           => n11, Q => present_val_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n52, CLK => CLK, R => n22, S 
                           => n9, Q => present_val_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n54, CLK => CLK, R => n22, S 
                           => n7, Q => present_val_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n56, CLK => CLK, R => n22, S 
                           => n5, Q => present_val_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n58, CLK => CLK, R => n22, S 
                           => n4, Q => present_val_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n60, CLK => CLK, R => n22, S 
                           => n3, Q => present_val_1_port);
   U4 : BUFX2 port map( A => RCV_DATA_6_port, Y => n1);
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n7 <= '1';
   n9 <= '1';
   n11 <= '1';
   n13 <= '1';
   n15 <= '1';
   U21 : INVX1 port map( A => RCV_DATA_7_port, Y => n17);
   U24 : INVX2 port map( A => n17, Y => n19);
   U25 : INVX2 port map( A => RST, Y => n22);
   U28 : AND2X2 port map( A => SHIFT_ENABLE, B => n25, Y => n20);
   U29 : INVX2 port map( A => present_val_7_port, Y => n31);
   U32 : INVX2 port map( A => present_val_6_port, Y => n34);
   U33 : INVX2 port map( A => present_val_5_port, Y => n37);
   U34 : INVX2 port map( A => present_val_4_port, Y => n40);
   U35 : INVX2 port map( A => present_val_3_port, Y => n43);
   U36 : INVX2 port map( A => present_val_2_port, Y => n45);
   U37 : INVX2 port map( A => present_val_1_port, Y => n46);
   U38 : INVX2 port map( A => present_val_0_port, Y => n47);
   U39 : INVX2 port map( A => BITSTUFF, Y => n25);
   U40 : MUX2X1 port map( B => n47, A => n46, S => n20, Y => n62);
   U41 : MUX2X1 port map( B => n46, A => n45, S => n20, Y => n60);
   U42 : MUX2X1 port map( B => n45, A => n43, S => n20, Y => n58);
   U43 : MUX2X1 port map( B => n43, A => n40, S => n20, Y => n56);
   U44 : MUX2X1 port map( B => n40, A => n37, S => n20, Y => n54);
   U45 : MUX2X1 port map( B => n37, A => n34, S => n20, Y => n52);
   U46 : MUX2X1 port map( B => n34, A => n31, S => n20, Y => n50);
   U47 : INVX2 port map( A => D_ORIG, Y => n28);
   U48 : MUX2X1 port map( B => n31, A => n28, S => n20, Y => n48);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_rcu_0 is

   port( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR : in std_logic
         ;  RX_CRC, RX_CHECK_CRC : in std_logic_vector (15 downto 0);  RCV_DATA
         : in std_logic_vector (7 downto 0);  RCVING, W_ENABLE, R_ERROR, 
         CRC_ERROR : out std_logic;  OPCODE : out std_logic_vector (1 downto 0)
         );

end rx_rcu_0;

architecture SYN_moore of rx_rcu_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal CRC_ERROR_port, state_3_port, state_2_port, state_1_port, 
      state_0_port, count_3_port, count_2_port, count_1_port, count_0_port, 
      nextstate_3_port, nextstate_2_port, nextstate_1_port, nextstate_0_port, 
      nxtR_ERROR, curR_ERROR, curCRC_ERROR, n1, n2, n3, n4, n5, n6, n7, n8, n9,
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n39, n40, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84, n85, n86, n89
      , n90, n91, n92, n93, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n152, n153, n154, 
      n155, n160, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244 : std_logic;

begin
   CRC_ERROR <= CRC_ERROR_port;
   
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => CLK, R => 
                           n43, S => n230, Q => state_3_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => CLK, R => 
                           n43, S => n231, Q => state_0_port);
   count_reg_0_inst : DFFSR port map( D => n221, CLK => CLK, R => n43, S => 
                           n232, Q => count_0_port);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => CLK, R => 
                           n43, S => n233, Q => state_2_port);
   curCRC_ERROR_reg : DFFPOSX1 port map( D => n234, CLK => CLK, Q => 
                           curCRC_ERROR);
   curR_ERROR_reg : DFFPOSX1 port map( D => n235, CLK => CLK, Q => curR_ERROR);
   R_ERROR_reg : DFFSR port map( D => nxtR_ERROR, CLK => CLK, R => n43, S => 
                           n236, Q => R_ERROR);
   CRC_ERROR_reg : DFFPOSX1 port map( D => n222, CLK => CLK, Q => 
                           CRC_ERROR_port);
   U16 : NAND2X1 port map( A => n244, B => n243, Y => nextstate_2_port);
   U19 : OAI21X1 port map( A => n5, B => n241, C => n35, Y => n242);
   U20 : NAND2X1 port map( A => n188, B => n189, Y => n241);
   U52 : AOI21X1 port map( A => CRC_ERROR_port, B => RST, C => n238, Y => n239)
                           ;
   U56 : OAI21X1 port map( A => n43, B => n224, C => n237, Y => n235);
   U79 : NOR2X1 port map( A => D_EDGE, B => n23, Y => n240);
   n236 <= '1';
   n233 <= '1';
   n232 <= '1';
   n231 <= '1';
   n230 <= '1';
   count_reg_2_inst : DFFSR port map( D => n228, CLK => CLK, R => n43, S => n12
                           , Q => count_2_port);
   count_reg_1_inst : DFFSR port map( D => n229, CLK => CLK, R => n43, S => n11
                           , Q => count_1_port);
   count_reg_3_inst : DFFSR port map( D => n227, CLK => CLK, R => n43, S => n10
                           , Q => count_3_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => CLK, R => 
                           n43, S => n9, Q => state_1_port);
   U3 : INVX2 port map( A => n117, Y => n119);
   U4 : AND2X2 port map( A => n56, B => n55, Y => n1);
   U5 : INVX1 port map( A => n1, Y => n136);
   U6 : AND2X2 port map( A => n62, B => n180, Y => n29);
   U7 : INVX4 port map( A => n40, Y => n58);
   U8 : BUFX4 port map( A => state_3_port, Y => n33);
   U9 : BUFX2 port map( A => n24, Y => n2);
   U10 : BUFX2 port map( A => n24, Y => n3);
   U11 : BUFX2 port map( A => n24, Y => n4);
   U12 : NAND2X1 port map( A => n217, B => n216, Y => n5);
   U13 : AND2X2 port map( A => n40, B => n170, Y => n6);
   U14 : AND2X2 port map( A => n119, B => n116, Y => n7);
   U15 : AND2X2 port map( A => n67, B => n39, Y => n8);
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   U23 : INVX2 port map( A => n15, Y => n13);
   U24 : INVX2 port map( A => n153, Y => n14);
   U25 : INVX1 port map( A => n6, Y => n15);
   U26 : NAND2X1 port map( A => n34, B => n4, Y => n16);
   U27 : NAND2X1 port map( A => n6, B => n3, Y => n17);
   U28 : BUFX2 port map( A => n33, Y => n18);
   U29 : INVX1 port map( A => n173, Y => n19);
   U30 : INVX2 port map( A => n19, Y => n20);
   U31 : INVX2 port map( A => n36, Y => n39);
   U32 : BUFX2 port map( A => n62, Y => n21);
   U33 : INVX2 port map( A => n36, Y => n23);
   U34 : BUFX2 port map( A => state_1_port, Y => n35);
   U35 : MUX2X1 port map( B => n111, A => n112, S => n189, Y => n227);
   U36 : INVX1 port map( A => n104, Y => n60);
   U37 : AND2X2 port map( A => n119, B => n110, Y => n22);
   U38 : NOR2X1 port map( A => n22, B => n109, Y => n111);
   U39 : INVX2 port map( A => state_2_port, Y => n36);
   U40 : AND2X2 port map( A => state_1_port, B => n36, Y => n24);
   U41 : INVX1 port map( A => n4, Y => n172);
   U42 : NAND2X1 port map( A => n105, B => n7, Y => n114);
   U43 : BUFX2 port map( A => n104, Y => n25);
   U44 : BUFX2 port map( A => n29, Y => n26);
   U45 : NAND2X1 port map( A => n8, B => n173, Y => n62);
   U46 : INVX1 port map( A => n180, Y => n184);
   U47 : INVX1 port map( A => n58, Y => n27);
   U48 : INVX1 port map( A => n114, Y => n106);
   U49 : INVX4 port map( A => n32, Y => n170);
   U50 : INVX1 port map( A => state_1_port, Y => n67);
   U51 : INVX2 port map( A => n126, Y => n28);
   U53 : INVX2 port map( A => RST, Y => n43);
   U54 : INVX1 port map( A => state_1_port, Y => n178);
   U55 : AND2X2 port map( A => SHIFT_ENABLE, B => n102, Y => n30);
   U57 : NOR2X1 port map( A => n40, B => n33, Y => n31);
   U58 : BUFX2 port map( A => state_3_port, Y => n32);
   U59 : AND2X2 port map( A => n33, B => n40, Y => n34);
   U60 : INVX1 port map( A => n34, Y => n153);
   U61 : BUFX4 port map( A => state_0_port, Y => n40);
   U62 : INVX1 port map( A => n108, Y => n105);
   U63 : INVX1 port map( A => n113, Y => n109);
   U64 : INVX1 port map( A => n182, Y => n126);
   U65 : NAND2X1 port map( A => n39, B => n170, Y => n65);
   U66 : INVX2 port map( A => n65, Y => n146);
   U67 : NAND2X1 port map( A => n35, B => n146, Y => n57);
   U68 : INVX2 port map( A => n57, Y => OPCODE(0));
   U69 : NAND2X1 port map( A => n33, B => n39, Y => n44);
   U70 : NOR2X1 port map( A => n40, B => n44, Y => n46);
   U71 : AOI21X1 port map( A => n23, B => n58, C => n18, Y => n45);
   U72 : MUX2X1 port map( B => n46, A => n45, S => n35, Y => n47);
   U73 : NAND2X1 port map( A => n6, B => n4, Y => n124);
   U74 : NAND2X1 port map( A => n34, B => n3, Y => n182);
   U75 : NAND2X1 port map( A => n124, B => n182, Y => n89);
   U76 : OR2X2 port map( A => n89, B => n47, Y => OPCODE(1));
   U77 : NAND2X1 port map( A => n33, B => n58, Y => n85);
   U78 : INVX2 port map( A => n85, Y => n173);
   U80 : INVX2 port map( A => RCV_DATA(1), Y => n49);
   U81 : INVX2 port map( A => RCV_DATA(2), Y => n48);
   U82 : NAND2X1 port map( A => n49, B => n48, Y => n52);
   U83 : INVX2 port map( A => RCV_DATA(0), Y => n50);
   U84 : NAND2X1 port map( A => RCV_DATA(7), B => n50, Y => n51);
   U85 : NOR2X1 port map( A => n52, B => n51, Y => n56);
   U86 : NOR2X1 port map( A => RCV_DATA(4), B => RCV_DATA(3), Y => n54);
   U87 : NOR2X1 port map( A => RCV_DATA(6), B => RCV_DATA(5), Y => n53);
   U88 : AND2X2 port map( A => n54, B => n53, Y => n55);
   U89 : NAND3X1 port map( A => n1, B => n2, C => n31, Y => n180);
   U90 : NAND2X1 port map( A => n29, B => n57, Y => W_ENABLE);
   U91 : NAND2X1 port map( A => n146, B => n58, Y => n166);
   U92 : NAND3X1 port map( A => n34, B => n23, C => n178, Y => n181);
   U93 : OAI21X1 port map( A => n35, B => n166, C => n181, Y => n122);
   U94 : INVX2 port map( A => n122, Y => n64);
   U95 : NAND2X1 port map( A => n4, B => n170, Y => n61);
   U96 : NOR2X1 port map( A => n33, B => n39, Y => n59);
   U97 : NAND3X1 port map( A => n40, B => n67, C => n59, Y => n171);
   U98 : NAND3X1 port map( A => n17, B => n16, C => n171, Y => n104);
   U99 : NAND3X1 port map( A => n21, B => n61, C => n60, Y => n63);
   U100 : INVX2 port map( A => n63, Y => n91);
   U101 : NAND3X1 port map( A => n35, B => n23, C => n6, Y => n130);
   U102 : NAND3X1 port map( A => n64, B => n91, C => n130, Y => RCVING);
   U103 : NAND2X1 port map( A => n240, B => n20, Y => n75);
   U104 : NAND2X1 port map( A => n75, B => n65, Y => n66);
   U105 : NAND3X1 port map( A => curR_ERROR, B => n178, C => n66, Y => n73);
   U106 : NOR2X1 port map( A => n27, B => n172, Y => n69);
   U107 : NAND2X1 port map( A => n1, B => n170, Y => n68);
   U108 : NAND2X1 port map( A => n69, B => n68, Y => n95);
   U109 : NAND2X1 port map( A => n28, B => n171, Y => n71);
   U110 : INVX2 port map( A => n166, Y => n145);
   U111 : NOR2X1 port map( A => count_3_port, B => n178, Y => n70);
   U112 : NOR3X1 port map( A => count_0_port, B => count_1_port, C => 
                           count_2_port, Y => n188);
   U113 : NAND2X1 port map( A => n70, B => n188, Y => n77);
   U114 : AOI22X1 port map( A => EOP, B => n71, C => n145, D => n77, Y => n72);
   U115 : NAND3X1 port map( A => n73, B => n95, C => n72, Y => nxtR_ERROR);
   U116 : INVX2 port map( A => n73, Y => n74);
   U117 : OAI21X1 port map( A => n43, B => n74, C => nxtR_ERROR, Y => n237);
   U118 : NAND2X1 port map( A => curCRC_ERROR, B => n43, Y => n80);
   U119 : NAND2X1 port map( A => n13, B => n23, Y => n81);
   U120 : NAND2X1 port map( A => n81, B => n75, Y => n76);
   U121 : NAND2X1 port map( A => n76, B => n178, Y => n98);
   U122 : INVX2 port map( A => n77, Y => n78);
   U123 : NAND2X1 port map( A => n145, B => n78, Y => n176);
   U124 : INVX2 port map( A => n176, Y => n79);
   U125 : NAND3X1 port map( A => n5, B => n43, C => n79, Y => n101);
   U126 : OAI21X1 port map( A => n80, B => n98, C => n101, Y => n238);
   U127 : INVX2 port map( A => count_3_port, Y => n189);
   U128 : INVX2 port map( A => n81, Y => n84);
   U129 : INVX2 port map( A => D_EDGE, Y => n82);
   U130 : AOI22X1 port map( A => n84, B => n82, C => n226, D => n145, Y => n86)
                           ;
   U131 : MUX2X1 port map( B => n86, A => n19, S => n35, Y => n93);
   U132 : NAND2X1 port map( A => n188, B => count_3_port, Y => n125);
   U133 : INVX2 port map( A => n125, Y => n123);
   U134 : NAND2X1 port map( A => n123, B => n89, Y => n90);
   U135 : OAI21X1 port map( A => n225, B => n91, C => n90, Y => n92);
   U136 : NOR2X1 port map( A => n93, B => n92, Y => n244);
   U137 : OAI21X1 port map( A => n242, B => n166, C => n95, Y => n97);
   U138 : NAND2X1 port map( A => EOP, B => n25, Y => n116);
   U139 : NAND2X1 port map( A => n116, B => n181, Y => n96);
   U140 : NOR2X1 port map( A => n97, B => n96, Y => n243);
   U141 : INVX2 port map( A => n98, Y => n99);
   U142 : OAI21X1 port map( A => RST, B => n99, C => curCRC_ERROR, Y => n100);
   U143 : NAND2X1 port map( A => n101, B => n100, Y => n234);
   U144 : AND2X2 port map( A => count_1_port, B => count_0_port, Y => n103);
   U145 : INVX2 port map( A => BITSTUFF, Y => n102);
   U146 : NAND2X1 port map( A => n103, B => n30, Y => n108);
   U147 : NAND2X1 port map( A => n25, B => n125, Y => n117);
   U148 : NAND2X1 port map( A => count_2_port, B => n106, Y => n112);
   U149 : INVX2 port map( A => count_2_port, Y => n110);
   U150 : INVX2 port map( A => n116, Y => n107);
   U151 : AOI21X1 port map( A => n119, B => n108, C => n107, Y => n113);
   U152 : MUX2X1 port map( B => n114, A => n113, S => count_2_port, Y => n228);
   U153 : NAND3X1 port map( A => n30, B => n119, C => n116, Y => n135);
   U154 : INVX2 port map( A => n135, Y => n115);
   U155 : NAND2X1 port map( A => count_0_port, B => n115, Y => n121);
   U156 : INVX2 port map( A => count_0_port, Y => n118);
   U157 : OAI21X1 port map( A => n30, B => n117, C => n116, Y => n133);
   U158 : AOI21X1 port map( A => n119, B => n118, C => n133, Y => n120);
   U159 : MUX2X1 port map( B => n121, A => n120, S => count_1_port, Y => n229);
   U161 : NAND2X1 port map( A => n122, B => EOP, Y => n132);
   U162 : NAND2X1 port map( A => n123, B => n226, Y => n141);
   U163 : OAI21X1 port map( A => n141, B => n171, C => n17, Y => n129);
   U164 : NAND3X1 port map( A => n226, B => n126, C => n125, Y => n127);
   U169 : NAND2X1 port map( A => n26, B => n127, Y => n128);
   U170 : OAI21X1 port map( A => n129, B => n128, C => n225, Y => n131);
   U171 : NAND3X1 port map( A => n132, B => n131, C => n130, Y => 
                           nextstate_1_port);
   U172 : INVX2 port map( A => n133, Y => n134);
   U173 : MUX2X1 port map( B => n135, A => n134, S => count_0_port, Y => n221);
   U174 : NOR2X1 port map( A => n226, B => n15, Y => n139);
   U175 : NAND2X1 port map( A => n31, B => n136, Y => n137);
   U176 : OAI21X1 port map( A => n153, B => n141, C => n137, Y => n138);
   U177 : OAI21X1 port map( A => n139, B => n138, C => n225, Y => n140);
   U178 : NAND2X1 port map( A => n3, B => n140, Y => n164);
   U179 : NOR2X1 port map( A => n141, B => BS_ERROR, Y => n142);
   U180 : AOI22X1 port map( A => n142, B => n13, C => n14, D => D_EDGE, Y => 
                           n144);
   U181 : NAND2X1 port map( A => EOP, B => n14, Y => n143);
   U182 : MUX2X1 port map( B => n144, A => n143, S => n23, Y => n152);
   U183 : AOI21X1 port map( A => D_EDGE, B => n146, C => n145, Y => n147);
   U184 : OAI21X1 port map( A => n27, B => n223, C => n147, Y => n148);
   U185 : NOR2X1 port map( A => n152, B => n148, Y => n155);
   U186 : AND2X2 port map( A => n23, B => n153, Y => n154);
   U187 : MUX2X1 port map( B => n155, A => n154, S => n35, Y => n160);
   U188 : NAND2X1 port map( A => n164, B => n160, Y => nextstate_0_port);
   U189 : NAND2X1 port map( A => D_EDGE, B => n27, Y => n165);
   U190 : OAI21X1 port map( A => n225, B => n170, C => n165, Y => n168);
   U191 : NOR2X1 port map( A => n226, B => n166, Y => n167);
   U192 : AOI21X1 port map( A => n23, B => n168, C => n167, Y => n169);
   U193 : OAI21X1 port map( A => n223, B => n170, C => n169, Y => n179);
   U194 : OAI21X1 port map( A => n20, B => n172, C => n171, Y => n174);
   U195 : NAND2X1 port map( A => BS_ERROR, B => n174, Y => n175);
   U196 : OAI21X1 port map( A => n5, B => n176, C => n175, Y => n177);
   U197 : AOI21X1 port map( A => n179, B => n178, C => n177, Y => n186);
   U198 : OAI21X1 port map( A => EOP, B => n28, C => n181, Y => n183);
   U199 : NOR2X1 port map( A => n184, B => n183, Y => n185);
   U200 : NAND2X1 port map( A => n186, B => n185, Y => nextstate_3_port);
   U201 : XNOR2X1 port map( A => RX_CHECK_CRC(10), B => RX_CRC(10), Y => n194);
   U202 : XNOR2X1 port map( A => RX_CHECK_CRC(9), B => RX_CRC(9), Y => n193);
   U203 : XOR2X1 port map( A => RX_CHECK_CRC(7), B => RX_CRC(7), Y => n191);
   U204 : XOR2X1 port map( A => RX_CHECK_CRC(8), B => RX_CRC(8), Y => n190);
   U205 : NOR2X1 port map( A => n191, B => n190, Y => n192);
   U206 : NAND3X1 port map( A => n194, B => n193, C => n192, Y => n201);
   U207 : XNOR2X1 port map( A => RX_CHECK_CRC(14), B => RX_CRC(14), Y => n199);
   U208 : XNOR2X1 port map( A => RX_CHECK_CRC(13), B => RX_CRC(13), Y => n198);
   U209 : XOR2X1 port map( A => RX_CHECK_CRC(11), B => RX_CRC(11), Y => n196);
   U210 : XOR2X1 port map( A => RX_CHECK_CRC(12), B => RX_CRC(12), Y => n195);
   U211 : NOR2X1 port map( A => n196, B => n195, Y => n197);
   U212 : NAND3X1 port map( A => n199, B => n198, C => n197, Y => n200);
   U213 : NOR2X1 port map( A => n201, B => n200, Y => n217);
   U214 : NOR2X1 port map( A => n218, B => RX_CHECK_CRC(0), Y => n202);
   U215 : OAI22X1 port map( A => RX_CRC(1), B => n202, C => n202, D => n220, Y 
                           => n208);
   U216 : AND2X1 port map( A => RX_CHECK_CRC(0), B => n218, Y => n203);
   U217 : OAI22X1 port map( A => n203, B => n219, C => RX_CHECK_CRC(1), D => 
                           n203, Y => n207);
   U218 : XOR2X1 port map( A => RX_CHECK_CRC(15), B => RX_CRC(15), Y => n205);
   U219 : XOR2X1 port map( A => RX_CHECK_CRC(2), B => RX_CRC(2), Y => n204);
   U220 : NOR2X1 port map( A => n205, B => n204, Y => n206);
   U221 : NAND3X1 port map( A => n208, B => n207, C => n206, Y => n215);
   U222 : XNOR2X1 port map( A => RX_CHECK_CRC(6), B => RX_CRC(6), Y => n213);
   U223 : XNOR2X1 port map( A => RX_CHECK_CRC(5), B => RX_CRC(5), Y => n212);
   U224 : XOR2X1 port map( A => RX_CHECK_CRC(3), B => RX_CRC(3), Y => n210);
   U225 : XOR2X1 port map( A => RX_CHECK_CRC(4), B => RX_CRC(4), Y => n209);
   U226 : NOR2X1 port map( A => n210, B => n209, Y => n211);
   U227 : NAND3X1 port map( A => n213, B => n212, C => n211, Y => n214);
   U228 : NOR2X1 port map( A => n215, B => n214, Y => n216);
   U229 : INVX2 port map( A => RX_CRC(0), Y => n218);
   U230 : INVX2 port map( A => RX_CRC(1), Y => n219);
   U231 : INVX2 port map( A => RX_CHECK_CRC(1), Y => n220);
   U232 : INVX2 port map( A => n239, Y => n222);
   U233 : INVX2 port map( A => n240, Y => n223);
   U234 : INVX2 port map( A => curR_ERROR, Y => n224);
   U235 : INVX2 port map( A => BS_ERROR, Y => n225);
   U236 : INVX2 port map( A => EOP, Y => n226);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_eopdetect_0 is

   port( DP1_RX, DM1_RX : in std_logic;  EOP : out std_logic);

end rx_eopdetect_0;

architecture SYN_Behavioral of rx_eopdetect_0 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;

begin
   
   U1 : NOR2X1 port map( A => DP1_RX, B => DM1_RX, Y => EOP);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_edgedetect_0 is

   port( CLK, RST, DP1_RX : in std_logic;  D_EDGE : out std_logic);

end rx_edgedetect_0;

architecture SYN_Behavioral of rx_edgedetect_0 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal DP_hold1, DP_hold2, n2, n4, n5, n6 : std_logic;

begin
   
   DP_hold1_reg : DFFSR port map( D => DP1_RX, CLK => CLK, R => n5, S => n2, Q 
                           => DP_hold1);
   DP_hold2_reg : DFFSR port map( D => DP_hold1, CLK => CLK, R => n6, S => n2, 
                           Q => DP_hold2);
   n6 <= '1';
   n5 <= '1';
   U4 : INVX2 port map( A => RST, Y => n2);
   U6 : XNOR2X1 port map( A => DP_hold2, B => DP_hold1, Y => n4);
   U7 : NOR2X1 port map( A => RST, B => n4, Y => D_EDGE);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_decode_0 is

   port( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP : in std_logic;  D_ORIG, BITSTUFF,
         BS_ERROR : out std_logic);

end rx_decode_0;

architecture SYN_moore of rx_decode_0 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal DP_hold1, DP_hold2, state_3_port, state_2_port, state_1_port, 
      state_0_port, N29, N30, N31, N32, n2, n3, n5, n6, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n18, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29_port, n30_port, n31_port, n32_port, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, BS_ERROR_port, n48, n49, n50, n51, n52, n53, n54 : 
      std_logic;

begin
   BS_ERROR <= BS_ERROR_port;
   
   DP_hold2_reg : DFFSR port map( D => n48, CLK => CLK, R => n52, S => n9, Q =>
                           DP_hold2);
   state_reg_3_inst : DFFSR port map( D => N32, CLK => CLK, R => n9, S => n53, 
                           Q => state_3_port);
   DP_hold1_reg : DFFSR port map( D => n49, CLK => CLK, R => n54, S => n9, Q =>
                           DP_hold1);
   n54 <= '1';
   n53 <= '1';
   n52 <= '1';
   U20 : NAND2X1 port map( A => n51, B => n41, Y => n49);
   U21 : AOI22X1 port map( A => DP_hold1, B => n42, C => DP1_RX, D => n50, Y =>
                           n51);
   U25 : XNOR2X1 port map( A => DP_hold1, B => DP_hold2, Y => D_ORIG);
   state_reg_0_inst : DFFSR port map( D => N29, CLK => CLK, R => n9, S => n5, Q
                           => state_0_port);
   state_reg_2_inst : DFFSR port map( D => N31, CLK => CLK, R => n9, S => n3, Q
                           => state_2_port);
   state_reg_1_inst : DFFSR port map( D => N30, CLK => CLK, R => n9, S => n2, Q
                           => state_1_port);
   n2 <= '1';
   n3 <= '1';
   n5 <= '1';
   U8 : INVX2 port map( A => RST, Y => n9);
   U10 : AND2X2 port map( A => state_1_port, B => state_2_port, Y => n6);
   U11 : MUX2X1 port map( B => DP_hold1, A => DP_hold2, S => n8, Y => n40);
   U12 : NAND2X1 port map( A => SHIFT_ENABLE, B => n50, Y => n8);
   U13 : INVX1 port map( A => SHIFT_ENABLE, Y => n31_port);
   U14 : AND2X1 port map( A => SHIFT_ENABLE, B => state_0_port, Y => n22);
   U15 : INVX2 port map( A => state_0_port, Y => n15);
   U16 : NOR2X1 port map( A => state_1_port, B => state_2_port, Y => n10);
   U17 : NAND3X1 port map( A => state_3_port, B => n15, C => n10, Y => n11);
   U18 : INVX2 port map( A => n11, Y => BS_ERROR_port);
   U19 : NAND2X1 port map( A => n6, B => n15, Y => n50);
   U22 : NOR2X1 port map( A => state_3_port, B => n50, Y => BITSTUFF);
   U23 : INVX2 port map( A => n50, Y => n42);
   U24 : OR2X2 port map( A => EOP, B => state_3_port, Y => n37);
   U26 : INVX2 port map( A => n37, Y => n41);
   U27 : INVX2 port map( A => DP1_RX, Y => n12);
   U28 : XOR2X1 port map( A => n12, B => DP_hold2, Y => n33);
   U29 : INVX2 port map( A => n33, Y => n24);
   U30 : NOR2X1 port map( A => state_0_port, B => n24, Y => n13);
   U31 : MUX2X1 port map( B => n13, A => n24, S => n6, Y => n14);
   U32 : MUX2X1 port map( B => n15, A => n14, S => SHIFT_ENABLE, Y => n16);
   U33 : AND2X2 port map( A => n41, B => n16, Y => N29);
   U34 : INVX2 port map( A => state_2_port, Y => n18);
   U35 : NAND3X1 port map( A => state_1_port, B => n33, C => n18, Y => n35);
   U36 : INVX2 port map( A => n35, Y => n23);
   U37 : INVX2 port map( A => state_1_port, Y => n32_port);
   U38 : NAND2X1 port map( A => n33, B => n32_port, Y => n20);
   U39 : AOI21X1 port map( A => SHIFT_ENABLE, B => n20, C => n18, Y => n21);
   U40 : AOI21X1 port map( A => n23, B => n22, C => n21, Y => n25);
   U41 : NAND2X1 port map( A => n24, B => n42, Y => n29_port);
   U42 : AOI21X1 port map( A => n25, B => n29_port, C => n37, Y => N31);
   U43 : NAND3X1 port map( A => n33, B => n42, C => SHIFT_ENABLE, Y => n28);
   U44 : INVX2 port map( A => EOP, Y => n26);
   U45 : NAND2X1 port map( A => BS_ERROR_port, B => n26, Y => n27);
   U46 : OAI21X1 port map( A => n37, B => n28, C => n27, Y => N32);
   U47 : INVX2 port map( A => n29_port, Y => n30_port);
   U48 : AOI21X1 port map( A => state_1_port, B => n31_port, C => n30_port, Y 
                           => n39);
   U49 : NAND3X1 port map( A => SHIFT_ENABLE, B => n33, C => n32_port, Y => n34
                           );
   U50 : MUX2X1 port map( B => n35, A => n34, S => state_0_port, Y => n36);
   U51 : INVX2 port map( A => n36, Y => n38);
   U52 : AOI21X1 port map( A => n39, B => n38, C => n37, Y => N30);
   U53 : NAND2X1 port map( A => n41, B => n40, Y => n48);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_accumulator_0 is

   port( CLK, RST : in std_logic;  RCV_DATA : in std_logic_vector (7 downto 0);
         W_ENABLE : in std_logic;  rx_CHECK_CRC : out std_logic_vector (15 
         downto 0));

end rx_accumulator_0;

architecture SYN_Behavioral of rx_accumulator_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, rx_CHECK_CRC_13_port, 
      rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, rx_CHECK_CRC_10_port, 
      rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, rx_CHECK_CRC_7_port, 
      rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, rx_CHECK_CRC_4_port, 
      rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, rx_CHECK_CRC_1_port, 
      rx_CHECK_CRC_0_port, n1, n2, n5, n8, n11, n14, n17, n20, n23, n56, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108 : std_logic;

begin
   rx_CHECK_CRC <= ( rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, 
      rx_CHECK_CRC_13_port, rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, 
      rx_CHECK_CRC_10_port, rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, 
      rx_CHECK_CRC_7_port, rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, 
      rx_CHECK_CRC_4_port, rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, 
      rx_CHECK_CRC_1_port, rx_CHECK_CRC_0_port );
   
   present_CHECK_CRC_reg_7_inst : DFFSR port map( D => n61, CLK => CLK, R => n5
                           , S => n62, Q => rx_CHECK_CRC_7_port);
   present_CHECK_CRC_reg_15_inst : DFFSR port map( D => n63, CLK => CLK, R => 
                           n5, S => n64, Q => rx_CHECK_CRC_15_port);
   present_CHECK_CRC_reg_6_inst : DFFSR port map( D => n65, CLK => CLK, R => n5
                           , S => n66, Q => rx_CHECK_CRC_6_port);
   present_CHECK_CRC_reg_14_inst : DFFSR port map( D => n67, CLK => CLK, R => 
                           n5, S => n68, Q => rx_CHECK_CRC_14_port);
   present_CHECK_CRC_reg_5_inst : DFFSR port map( D => n69, CLK => CLK, R => n5
                           , S => n70, Q => rx_CHECK_CRC_5_port);
   present_CHECK_CRC_reg_13_inst : DFFSR port map( D => n71, CLK => CLK, R => 
                           n5, S => n72, Q => rx_CHECK_CRC_13_port);
   present_CHECK_CRC_reg_4_inst : DFFSR port map( D => n73, CLK => CLK, R => n5
                           , S => n74, Q => rx_CHECK_CRC_4_port);
   present_CHECK_CRC_reg_12_inst : DFFSR port map( D => n75, CLK => CLK, R => 
                           n5, S => n76, Q => rx_CHECK_CRC_12_port);
   present_CHECK_CRC_reg_3_inst : DFFSR port map( D => n77, CLK => CLK, R => n5
                           , S => n78, Q => rx_CHECK_CRC_3_port);
   present_CHECK_CRC_reg_11_inst : DFFSR port map( D => n79, CLK => CLK, R => 
                           n5, S => n80, Q => rx_CHECK_CRC_11_port);
   present_CHECK_CRC_reg_2_inst : DFFSR port map( D => n81, CLK => CLK, R => n5
                           , S => n82, Q => rx_CHECK_CRC_2_port);
   present_CHECK_CRC_reg_10_inst : DFFSR port map( D => n83, CLK => CLK, R => 
                           n5, S => n84, Q => rx_CHECK_CRC_10_port);
   present_CHECK_CRC_reg_1_inst : DFFSR port map( D => n85, CLK => CLK, R => n5
                           , S => n86, Q => rx_CHECK_CRC_1_port);
   present_CHECK_CRC_reg_9_inst : DFFSR port map( D => n87, CLK => CLK, R => n5
                           , S => n88, Q => rx_CHECK_CRC_9_port);
   present_CHECK_CRC_reg_0_inst : DFFSR port map( D => n89, CLK => CLK, R => n5
                           , S => n90, Q => rx_CHECK_CRC_0_port);
   present_CHECK_CRC_reg_8_inst : DFFSR port map( D => n91, CLK => CLK, R => n5
                           , S => n92, Q => rx_CHECK_CRC_8_port);
   U2 : OAI21X1 port map( A => n8, B => n60, C => n108, Y => n91);
   U3 : NAND2X1 port map( A => rx_CHECK_CRC_8_port, B => n8, Y => n108);
   U4 : OAI21X1 port map( A => n2, B => n60, C => n107, Y => n89);
   U5 : NAND2X1 port map( A => RCV_DATA(0), B => n2, Y => n107);
   U7 : OAI21X1 port map( A => n8, B => n59, C => n106, Y => n87);
   U8 : NAND2X1 port map( A => rx_CHECK_CRC_9_port, B => n8, Y => n106);
   U9 : OAI21X1 port map( A => n2, B => n59, C => n105, Y => n85);
   U10 : NAND2X1 port map( A => RCV_DATA(1), B => n2, Y => n105);
   U12 : OAI21X1 port map( A => n8, B => n56, C => n104, Y => n83);
   U13 : NAND2X1 port map( A => rx_CHECK_CRC_10_port, B => n8, Y => n104);
   U14 : OAI21X1 port map( A => n2, B => n56, C => n103, Y => n81);
   U15 : NAND2X1 port map( A => RCV_DATA(2), B => n2, Y => n103);
   U17 : OAI21X1 port map( A => n8, B => n23, C => n102, Y => n79);
   U18 : NAND2X1 port map( A => rx_CHECK_CRC_11_port, B => n8, Y => n102);
   U19 : OAI21X1 port map( A => n2, B => n23, C => n101, Y => n77);
   U20 : NAND2X1 port map( A => RCV_DATA(3), B => n2, Y => n101);
   U22 : OAI21X1 port map( A => n8, B => n20, C => n100, Y => n75);
   U23 : NAND2X1 port map( A => rx_CHECK_CRC_12_port, B => n8, Y => n100);
   U24 : OAI21X1 port map( A => n2, B => n20, C => n99, Y => n73);
   U25 : NAND2X1 port map( A => RCV_DATA(4), B => n2, Y => n99);
   U27 : OAI21X1 port map( A => n8, B => n17, C => n98, Y => n71);
   U28 : NAND2X1 port map( A => rx_CHECK_CRC_13_port, B => n8, Y => n98);
   U29 : OAI21X1 port map( A => n2, B => n17, C => n97, Y => n69);
   U30 : NAND2X1 port map( A => RCV_DATA(5), B => n2, Y => n97);
   U32 : OAI21X1 port map( A => n8, B => n14, C => n96, Y => n67);
   U33 : NAND2X1 port map( A => rx_CHECK_CRC_14_port, B => n8, Y => n96);
   U34 : OAI21X1 port map( A => n2, B => n14, C => n95, Y => n65);
   U35 : NAND2X1 port map( A => RCV_DATA(6), B => n2, Y => n95);
   U37 : OAI21X1 port map( A => n8, B => n11, C => n94, Y => n63);
   U38 : NAND2X1 port map( A => rx_CHECK_CRC_15_port, B => n8, Y => n94);
   U41 : OAI21X1 port map( A => n2, B => n11, C => n93, Y => n61);
   U42 : NAND2X1 port map( A => RCV_DATA(7), B => n2, Y => n93);
   n92 <= '1';
   n90 <= '1';
   n88 <= '1';
   n86 <= '1';
   n84 <= '1';
   n82 <= '1';
   n80 <= '1';
   n78 <= '1';
   n76 <= '1';
   n74 <= '1';
   n72 <= '1';
   n70 <= '1';
   n68 <= '1';
   n66 <= '1';
   n64 <= '1';
   n62 <= '1';
   U6 : INVX4 port map( A => n2, Y => n8);
   U11 : INVX4 port map( A => n1, Y => n2);
   U16 : INVX1 port map( A => W_ENABLE, Y => n1);
   U21 : INVX2 port map( A => RST, Y => n5);
   U26 : INVX2 port map( A => rx_CHECK_CRC_7_port, Y => n11);
   U31 : INVX2 port map( A => rx_CHECK_CRC_6_port, Y => n14);
   U36 : INVX2 port map( A => rx_CHECK_CRC_5_port, Y => n17);
   U39 : INVX2 port map( A => rx_CHECK_CRC_4_port, Y => n20);
   U40 : INVX2 port map( A => rx_CHECK_CRC_3_port, Y => n23);
   U43 : INVX2 port map( A => rx_CHECK_CRC_2_port, Y => n56);
   U60 : INVX2 port map( A => rx_CHECK_CRC_1_port, Y => n59);
   U61 : INVX2 port map( A => rx_CHECK_CRC_0_port, Y => n60);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_CRC_CALC_0 is

   port( CLK, RST, W_ENABLE : in std_logic;  OPCODE : in std_logic_vector (1 
         downto 0);  RCV_DATA : in std_logic_vector (7 downto 0);  RX_CRC : out
         std_logic_vector (15 downto 0));

end rx_CRC_CALC_0;

architecture SYN_moore of rx_CRC_CALC_0 is

   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port, current_crc_15_port, 
      current_crc_14_port, current_crc_13_port, current_crc_12_port, 
      current_crc_11_port, current_crc_10_port, current_crc_9_port, 
      current_crc_8_port, current_crc_7_port, current_crc_6_port, 
      current_crc_5_port, current_crc_4_port, current_crc_3_port, 
      current_crc_2_port, current_crc_1_port, current_crc_0_port, 
      cache_1_15_port, cache_1_14_port, cache_1_13_port, cache_1_12_port, 
      cache_1_11_port, cache_1_10_port, cache_1_9_port, cache_1_8_port, 
      cache_1_7_port, cache_1_6_port, cache_1_5_port, cache_1_4_port, 
      cache_1_3_port, cache_1_2_port, cache_1_1_port, cache_1_0_port, n1, n2, 
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n100, n102, n104, n106, n108, n110, n112, 
      n114, n116, n118, n120, n122, n124, n126, n128, n130, n131, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n_1021, n_1022, n_1023 : 
      std_logic;

begin
   RX_CRC <= ( RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port );
   
   cache_1_reg_0_inst : DFFPOSX1 port map( D => n186, CLK => CLK, Q => 
                           cache_1_0_port);
   cache_1_reg_8_inst : DFFPOSX1 port map( D => n187, CLK => CLK, Q => 
                           cache_1_8_port);
   cache_1_reg_15_inst : DFFPOSX1 port map( D => n188, CLK => CLK, Q => 
                           cache_1_15_port);
   cache_1_reg_1_inst : DFFPOSX1 port map( D => n189, CLK => CLK, Q => 
                           cache_1_1_port);
   cache_1_reg_9_inst : DFFPOSX1 port map( D => n190, CLK => CLK, Q => 
                           cache_1_9_port);
   cache_1_reg_2_inst : DFFPOSX1 port map( D => n191, CLK => CLK, Q => 
                           cache_1_2_port);
   cache_1_reg_10_inst : DFFPOSX1 port map( D => n192, CLK => CLK, Q => 
                           cache_1_10_port);
   cache_1_reg_3_inst : DFFPOSX1 port map( D => n193, CLK => CLK, Q => 
                           cache_1_3_port);
   cache_1_reg_11_inst : DFFPOSX1 port map( D => n194, CLK => CLK, Q => 
                           cache_1_11_port);
   cache_1_reg_4_inst : DFFPOSX1 port map( D => n195, CLK => CLK, Q => 
                           cache_1_4_port);
   cache_1_reg_12_inst : DFFPOSX1 port map( D => n196, CLK => CLK, Q => 
                           cache_1_12_port);
   cache_1_reg_5_inst : DFFPOSX1 port map( D => n197, CLK => CLK, Q => 
                           cache_1_5_port);
   cache_1_reg_13_inst : DFFPOSX1 port map( D => n198, CLK => CLK, Q => 
                           cache_1_13_port);
   cache_1_reg_6_inst : DFFPOSX1 port map( D => n199, CLK => CLK, Q => 
                           cache_1_6_port);
   cache_1_reg_14_inst : DFFPOSX1 port map( D => n200, CLK => CLK, Q => 
                           cache_1_14_port);
   cache_1_reg_7_inst : DFFPOSX1 port map( D => n201, CLK => CLK, Q => 
                           cache_1_7_port);
   cache_2_reg_15_inst : DFFPOSX1 port map( D => n202, CLK => CLK, Q => 
                           RX_CRC_15_port);
   cache_2_reg_14_inst : DFFPOSX1 port map( D => n203, CLK => CLK, Q => 
                           RX_CRC_14_port);
   cache_2_reg_13_inst : DFFPOSX1 port map( D => n204, CLK => CLK, Q => 
                           RX_CRC_13_port);
   cache_2_reg_12_inst : DFFPOSX1 port map( D => n205, CLK => CLK, Q => 
                           RX_CRC_12_port);
   cache_2_reg_11_inst : DFFPOSX1 port map( D => n206, CLK => CLK, Q => 
                           RX_CRC_11_port);
   cache_2_reg_10_inst : DFFPOSX1 port map( D => n207, CLK => CLK, Q => 
                           RX_CRC_10_port);
   cache_2_reg_9_inst : DFFPOSX1 port map( D => n208, CLK => CLK, Q => 
                           RX_CRC_9_port);
   cache_2_reg_8_inst : DFFPOSX1 port map( D => n209, CLK => CLK, Q => 
                           RX_CRC_8_port);
   cache_2_reg_7_inst : DFFPOSX1 port map( D => n210, CLK => CLK, Q => 
                           RX_CRC_7_port);
   cache_2_reg_6_inst : DFFPOSX1 port map( D => n211, CLK => CLK, Q => 
                           RX_CRC_6_port);
   cache_2_reg_5_inst : DFFPOSX1 port map( D => n212, CLK => CLK, Q => 
                           RX_CRC_5_port);
   cache_2_reg_4_inst : DFFPOSX1 port map( D => n213, CLK => CLK, Q => 
                           RX_CRC_4_port);
   cache_2_reg_3_inst : DFFPOSX1 port map( D => n214, CLK => CLK, Q => 
                           RX_CRC_3_port);
   cache_2_reg_2_inst : DFFPOSX1 port map( D => n215, CLK => CLK, Q => 
                           RX_CRC_2_port);
   cache_2_reg_1_inst : DFFPOSX1 port map( D => n216, CLK => CLK, Q => 
                           RX_CRC_1_port);
   cache_2_reg_0_inst : DFFPOSX1 port map( D => n217, CLK => CLK, Q => 
                           RX_CRC_0_port);
   current_crc_reg_5_inst : DFFSR port map( D => n175, CLK => CLK, R => n30, S 
                           => n16, Q => current_crc_5_port);
   current_crc_reg_3_inst : DFFSR port map( D => n173, CLK => CLK, R => n30, S 
                           => n15, Q => current_crc_3_port);
   current_crc_reg_15_inst : DFFSR port map( D => n185, CLK => CLK, R => n30, S
                           => n14, Q => current_crc_15_port);
   current_crc_reg_14_inst : DFFSR port map( D => n184, CLK => CLK, R => n30, S
                           => n13, Q => current_crc_14_port);
   current_crc_reg_13_inst : DFFSR port map( D => n183, CLK => CLK, R => n30, S
                           => n12, Q => current_crc_13_port);
   current_crc_reg_10_inst : DFFSR port map( D => n180, CLK => CLK, R => n30, S
                           => n11, Q => current_crc_10_port);
   current_crc_reg_9_inst : DFFSR port map( D => n179, CLK => CLK, R => n30, S 
                           => n10, Q => current_crc_9_port);
   current_crc_reg_4_inst : DFFSR port map( D => n174, CLK => CLK, R => n30, S 
                           => n9, Q => current_crc_4_port);
   current_crc_reg_0_inst : DFFSR port map( D => n170, CLK => CLK, R => n30, S 
                           => n8, Q => current_crc_0_port);
   current_crc_reg_12_inst : DFFSR port map( D => n182, CLK => CLK, R => n30, S
                           => n7, Q => current_crc_12_port);
   current_crc_reg_11_inst : DFFSR port map( D => n181, CLK => CLK, R => n30, S
                           => n6, Q => current_crc_11_port);
   current_crc_reg_8_inst : DFFSR port map( D => n178, CLK => CLK, R => n30, S 
                           => n5, Q => current_crc_8_port);
   current_crc_reg_6_inst : DFFSR port map( D => n176, CLK => CLK, R => n30, S 
                           => n4, Q => current_crc_6_port);
   current_crc_reg_2_inst : DFFSR port map( D => n172, CLK => CLK, R => n30, S 
                           => n3, Q => current_crc_2_port);
   current_crc_reg_1_inst : DFFSR port map( D => n171, CLK => CLK, R => n30, S 
                           => n2, Q => current_crc_1_port);
   current_crc_reg_7_inst : DFFSR port map( D => n177, CLK => CLK, R => n30, S 
                           => n1, Q => current_crc_7_port);
   U3 : INVX2 port map( A => n79, Y => n167);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   U20 : INVX8 port map( A => n29, Y => n26);
   U21 : INVX4 port map( A => n160, Y => n29);
   U22 : AND2X2 port map( A => W_ENABLE, B => OPCODE(0), Y => n17);
   U23 : INVX8 port map( A => n29, Y => n27);
   U24 : INVX1 port map( A => OPCODE(1), Y => n51);
   U25 : INVX2 port map( A => n18, Y => n24);
   U26 : INVX2 port map( A => n18, Y => n25);
   U27 : INVX2 port map( A => n29, Y => n28);
   U28 : AND2X2 port map( A => n52, B => n79, Y => n18);
   U29 : INVX2 port map( A => RST, Y => n30);
   U30 : XNOR2X1 port map( A => n58, B => n23, Y => n59);
   U31 : XNOR2X1 port map( A => RCV_DATA(6), B => current_crc_14_port, Y => 
                           n156);
   U32 : XNOR2X1 port map( A => RCV_DATA(7), B => current_crc_15_port, Y => 
                           n124);
   U33 : XOR2X1 port map( A => RCV_DATA(0), B => current_crc_8_port, Y => n19);
   U34 : XNOR2X1 port map( A => RCV_DATA(5), B => current_crc_13_port, Y => n58
                           );
   U35 : XOR2X1 port map( A => RCV_DATA(1), B => current_crc_9_port, Y => n20);
   U36 : XOR2X1 port map( A => RCV_DATA(3), B => current_crc_11_port, Y => n21)
                           ;
   U37 : XOR2X1 port map( A => RCV_DATA(2), B => current_crc_10_port, Y => n22)
                           ;
   U38 : XOR2X1 port map( A => RCV_DATA(4), B => current_crc_12_port, Y => n23)
                           ;
   U39 : INVX2 port map( A => RX_CRC_0_port, Y => n33);
   U40 : INVX2 port map( A => cache_1_0_port, Y => n161);
   U41 : NOR2X1 port map( A => RST, B => OPCODE(1), Y => n31);
   U42 : NAND2X1 port map( A => n31, B => n17, Y => n32);
   U43 : INVX2 port map( A => n32, Y => n160);
   U44 : MUX2X1 port map( B => n33, A => n161, S => n26, Y => n217);
   U45 : INVX2 port map( A => RX_CRC_1_port, Y => n34);
   U46 : INVX2 port map( A => cache_1_1_port, Y => n116);
   U47 : MUX2X1 port map( B => n34, A => n116, S => n26, Y => n216);
   U48 : INVX2 port map( A => RX_CRC_2_port, Y => n35);
   U49 : INVX2 port map( A => cache_1_2_port, Y => n100);
   U50 : MUX2X1 port map( B => n35, A => n100, S => n26, Y => n215);
   U51 : INVX2 port map( A => RX_CRC_3_port, Y => n36);
   U52 : INVX2 port map( A => cache_1_3_port, Y => n77);
   U53 : MUX2X1 port map( B => n36, A => n77, S => n26, Y => n214);
   U54 : INVX2 port map( A => RX_CRC_4_port, Y => n37);
   U55 : INVX2 port map( A => cache_1_4_port, Y => n70);
   U56 : MUX2X1 port map( B => n37, A => n70, S => n26, Y => n213);
   U57 : INVX2 port map( A => RX_CRC_5_port, Y => n38);
   U58 : INVX2 port map( A => cache_1_5_port, Y => n65);
   U59 : MUX2X1 port map( B => n38, A => n65, S => n26, Y => n212);
   U60 : INVX2 port map( A => RX_CRC_6_port, Y => n39);
   U61 : INVX2 port map( A => cache_1_6_port, Y => n57);
   U62 : MUX2X1 port map( B => n39, A => n57, S => n26, Y => n211);
   U63 : INVX2 port map( A => RX_CRC_7_port, Y => n40);
   U64 : INVX2 port map( A => cache_1_7_port, Y => n49);
   U65 : MUX2X1 port map( B => n40, A => n49, S => n26, Y => n210);
   U66 : INVX2 port map( A => RX_CRC_8_port, Y => n41);
   U67 : INVX2 port map( A => cache_1_8_port, Y => n155);
   U68 : MUX2X1 port map( B => n41, A => n155, S => n26, Y => n209);
   U69 : INVX2 port map( A => RX_CRC_9_port, Y => n42);
   U70 : INVX2 port map( A => cache_1_9_port, Y => n108);
   U71 : MUX2X1 port map( B => n42, A => n108, S => n26, Y => n208);
   U72 : INVX2 port map( A => RX_CRC_10_port, Y => n43);
   U73 : INVX2 port map( A => cache_1_10_port, Y => n80);
   U74 : MUX2X1 port map( B => n43, A => n80, S => n26, Y => n207);
   U75 : INVX2 port map( A => RX_CRC_11_port, Y => n44);
   U76 : INVX2 port map( A => cache_1_11_port, Y => n74);
   U77 : MUX2X1 port map( B => n44, A => n74, S => n26, Y => n206);
   U78 : INVX2 port map( A => RX_CRC_12_port, Y => n45);
   U79 : INVX2 port map( A => cache_1_12_port, Y => n67);
   U80 : MUX2X1 port map( B => n45, A => n67, S => n26, Y => n205);
   U81 : INVX2 port map( A => RX_CRC_13_port, Y => n46);
   U82 : INVX2 port map( A => cache_1_13_port, Y => n62);
   U83 : MUX2X1 port map( B => n46, A => n62, S => n27, Y => n204);
   U84 : INVX2 port map( A => RX_CRC_14_port, Y => n47);
   U85 : INVX2 port map( A => cache_1_14_port, Y => n54);
   U86 : MUX2X1 port map( B => n47, A => n54, S => n27, Y => n203);
   U87 : INVX2 port map( A => RX_CRC_15_port, Y => n48);
   U88 : INVX2 port map( A => cache_1_15_port, Y => n148);
   U89 : MUX2X1 port map( B => n48, A => n148, S => n27, Y => n202);
   U90 : INVX2 port map( A => current_crc_7_port, Y => n53);
   U91 : MUX2X1 port map( B => n49, A => n53, S => n27, Y => n201);
   U92 : INVX2 port map( A => n156, Y => n50);
   U93 : XOR2X1 port map( A => n58, B => n50, Y => n164);
   U94 : NAND2X1 port map( A => n17, B => n51, Y => n79);
   U95 : NAND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n52);
   U96 : OAI22X1 port map( A => n164, B => n79, C => n24, D => n53, Y => n177);
   U97 : INVX2 port map( A => current_crc_14_port, Y => n56);
   U98 : MUX2X1 port map( B => n54, A => n56, S => n27, Y => n200);
   U99 : NAND2X1 port map( A => current_crc_6_port, B => n167, Y => n55);
   U100 : OAI21X1 port map( A => n25, B => n56, C => n55, Y => n184);
   U101 : INVX2 port map( A => current_crc_6_port, Y => n61);
   U102 : MUX2X1 port map( B => n57, A => n61, S => n27, Y => n199);
   U103 : NAND2X1 port map( A => n167, B => n59, Y => n60);
   U104 : OAI21X1 port map( A => n24, B => n61, C => n60, Y => n176);
   U105 : INVX2 port map( A => current_crc_13_port, Y => n64);
   U106 : MUX2X1 port map( B => n62, A => n64, S => n27, Y => n198);
   U107 : NAND2X1 port map( A => current_crc_5_port, B => n167, Y => n63);
   U108 : OAI21X1 port map( A => n25, B => n64, C => n63, Y => n183);
   U109 : INVX2 port map( A => current_crc_5_port, Y => n66);
   U110 : MUX2X1 port map( B => n65, A => n66, S => n27, Y => n197);
   U111 : XNOR2X1 port map( A => n23, B => n21, Y => n118);
   U112 : OAI22X1 port map( A => n118, B => n79, C => n25, D => n66, Y => n175)
                           ;
   U113 : INVX2 port map( A => current_crc_12_port, Y => n69);
   U114 : MUX2X1 port map( B => n67, A => n69, S => n27, Y => n196);
   U115 : NAND2X1 port map( A => current_crc_4_port, B => n167, Y => n68);
   U116 : OAI21X1 port map( A => n24, B => n69, C => n68, Y => n182);
   U117 : INVX2 port map( A => current_crc_4_port, Y => n73);
   U118 : MUX2X1 port map( B => n70, A => n73, S => n27, Y => n195);
   U119 : XOR2X1 port map( A => n21, B => n22, Y => n71);
   U120 : NAND2X1 port map( A => n167, B => n71, Y => n72);
   U121 : OAI21X1 port map( A => n25, B => n73, C => n72, Y => n174);
   U122 : INVX2 port map( A => current_crc_11_port, Y => n76);
   U123 : MUX2X1 port map( B => n74, A => n76, S => n27, Y => n194);
   U124 : NAND2X1 port map( A => current_crc_3_port, B => n167, Y => n75);
   U125 : OAI21X1 port map( A => n24, B => n76, C => n75, Y => n181);
   U126 : INVX2 port map( A => current_crc_3_port, Y => n78);
   U127 : MUX2X1 port map( B => n77, A => n78, S => n27, Y => n193);
   U128 : XNOR2X1 port map( A => n22, B => n20, Y => n122);
   U129 : OAI22X1 port map( A => n122, B => n79, C => n24, D => n78, Y => n173)
                           ;
   U130 : INVX2 port map( A => current_crc_10_port, Y => n82);
   U131 : MUX2X1 port map( B => n80, A => n82, S => n27, Y => n192);
   U132 : NAND2X1 port map( A => current_crc_2_port, B => n167, Y => n81);
   U133 : OAI21X1 port map( A => n25, B => n82, C => n81, Y => n180);
   U134 : INVX2 port map( A => current_crc_2_port, Y => n106);
   U135 : MUX2X1 port map( B => n100, A => n106, S => n28, Y => n191);
   U136 : XOR2X1 port map( A => n19, B => n20, Y => n102);
   U137 : NAND2X1 port map( A => n167, B => n102, Y => n104);
   U138 : OAI21X1 port map( A => n24, B => n106, C => n104, Y => n172);
   U139 : INVX2 port map( A => current_crc_9_port, Y => n114);
   U140 : MUX2X1 port map( B => n108, A => n114, S => n28, Y => n190);
   U141 : INVX2 port map( A => n124, Y => n162);
   U142 : INVX2 port map( A => current_crc_1_port, Y => n131);
   U143 : XNOR2X1 port map( A => n162, B => n131, Y => n110);
   U144 : NAND2X1 port map( A => n167, B => n110, Y => n112);
   U145 : OAI21X1 port map( A => n25, B => n114, C => n112, Y => n179);
   U146 : MUX2X1 port map( B => n116, A => n131, S => n28, Y => n189);
   U147 : INVX2 port map( A => n118, Y => n120);
   U148 : XOR2X1 port map( A => n122, B => n120, Y => n163);
   U149 : INVX2 port map( A => n163, Y => n151);
   U150 : XNOR2X1 port map( A => n164, B => n124, Y => n126);
   U151 : XNOR2X1 port map( A => n151, B => n126, Y => n128);
   U152 : NAND2X1 port map( A => n167, B => n128, Y => n130);
   U153 : OAI21X1 port map( A => n24, B => n131, C => n130, Y => n171);
   U154 : INVX2 port map( A => current_crc_15_port, Y => n154);
   U155 : MUX2X1 port map( B => n148, A => n154, S => n28, Y => n188);
   U156 : FAX1 port map( A => current_crc_7_port, B => n19, C => n162, YC => 
                           n_1021, YS => n149);
   U157 : XNOR2X1 port map( A => n149, B => n164, Y => n150);
   U158 : XOR2X1 port map( A => n151, B => n150, Y => n152);
   U159 : NAND2X1 port map( A => n167, B => n152, Y => n153);
   U160 : OAI21X1 port map( A => n25, B => n154, C => n153, Y => n185);
   U161 : INVX2 port map( A => current_crc_8_port, Y => n159);
   U162 : MUX2X1 port map( B => n155, A => n159, S => n28, Y => n187);
   U163 : INVX2 port map( A => current_crc_0_port, Y => n169);
   U164 : FAX1 port map( A => n162, B => n169, C => n156, YC => n_1022, YS => 
                           n157);
   U165 : NAND2X1 port map( A => n167, B => n157, Y => n158);
   U166 : OAI21X1 port map( A => n24, B => n159, C => n158, Y => n178);
   U167 : MUX2X1 port map( B => n161, A => n169, S => n28, Y => n186);
   U168 : XOR2X1 port map( A => n19, B => n162, Y => n165);
   U169 : FAX1 port map( A => n165, B => n164, C => n163, YC => n_1023, YS => 
                           n166);
   U170 : NAND2X1 port map( A => n167, B => n166, Y => n168);
   U171 : OAI21X1 port map( A => n25, B => n169, C => n168, Y => n170);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RFIFO_0 is

   port( CLK, RST, W_ENABLE, R_ENABLE : in std_logic;  RCV_DATA : in 
         std_logic_vector (7 downto 0);  RCV_OPCODE : in std_logic_vector (1 
         downto 0);  DATA : out std_logic_vector (7 downto 0);  OUT_OPCODE : 
         out std_logic_vector (1 downto 0);  BYTE_COUNT : out std_logic_vector 
         (4 downto 0);  EMPTY, FULL : out std_logic);

end RFIFO_0;

architecture SYN_BRFIFO of RFIFO_0 is

   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, 
      DATA_3_port, DATA_2_port, DATA_1_port, DATA_0_port, OUT_OPCODE_1_port, 
      OUT_OPCODE_0_port, EMPTY_port, FULL_port, readptr_4_port, readptr_3_port,
      readptr_2_port, readptr_1_port, readptr_0_port, writeptr_4_port, 
      writeptr_3_port, writeptr_2_port, writeptr_1_port, writeptr_0_port, state
      , opcode_0_1_port, opcode_0_0_port, opcode_1_1_port, opcode_1_0_port, 
      opcode_2_1_port, opcode_2_0_port, opcode_3_1_port, opcode_3_0_port, 
      opcode_4_1_port, opcode_4_0_port, opcode_5_1_port, opcode_5_0_port, 
      opcode_6_1_port, opcode_6_0_port, opcode_7_1_port, opcode_7_0_port, 
      opcode_8_1_port, opcode_8_0_port, opcode_9_1_port, opcode_9_0_port, 
      opcode_10_1_port, opcode_10_0_port, opcode_11_1_port, opcode_11_0_port, 
      opcode_12_1_port, opcode_12_0_port, opcode_13_1_port, opcode_13_0_port, 
      opcode_14_1_port, opcode_14_0_port, opcode_15_1_port, opcode_15_0_port, 
      opcode_16_1_port, opcode_16_0_port, opcode_17_1_port, opcode_17_0_port, 
      opcode_18_1_port, opcode_18_0_port, opcode_19_1_port, opcode_19_0_port, 
      opcode_20_1_port, opcode_20_0_port, opcode_21_1_port, opcode_21_0_port, 
      opcode_22_1_port, opcode_22_0_port, opcode_23_1_port, opcode_23_0_port, 
      opcode_24_1_port, opcode_24_0_port, opcode_25_1_port, opcode_25_0_port, 
      opcode_26_1_port, opcode_26_0_port, opcode_27_1_port, opcode_27_0_port, 
      opcode_28_1_port, opcode_28_0_port, opcode_29_1_port, opcode_29_0_port, 
      opcode_30_1_port, opcode_30_0_port, opcode_31_1_port, opcode_31_0_port, 
      memory_0_7_port, memory_0_6_port, memory_0_5_port, memory_0_4_port, 
      memory_0_3_port, memory_0_2_port, memory_0_1_port, memory_0_0_port, 
      memory_1_7_port, memory_1_6_port, memory_1_5_port, memory_1_4_port, 
      memory_1_3_port, memory_1_2_port, memory_1_1_port, memory_1_0_port, 
      memory_2_7_port, memory_2_6_port, memory_2_5_port, memory_2_4_port, 
      memory_2_3_port, memory_2_2_port, memory_2_1_port, memory_2_0_port, 
      memory_3_7_port, memory_3_6_port, memory_3_5_port, memory_3_4_port, 
      memory_3_3_port, memory_3_2_port, memory_3_1_port, memory_3_0_port, 
      memory_4_7_port, memory_4_6_port, memory_4_5_port, memory_4_4_port, 
      memory_4_3_port, memory_4_2_port, memory_4_1_port, memory_4_0_port, 
      memory_5_7_port, memory_5_6_port, memory_5_5_port, memory_5_4_port, 
      memory_5_3_port, memory_5_2_port, memory_5_1_port, memory_5_0_port, 
      memory_6_7_port, memory_6_6_port, memory_6_5_port, memory_6_4_port, 
      memory_6_3_port, memory_6_2_port, memory_6_1_port, memory_6_0_port, 
      memory_7_7_port, memory_7_6_port, memory_7_5_port, memory_7_4_port, 
      memory_7_3_port, memory_7_2_port, memory_7_1_port, memory_7_0_port, 
      memory_8_7_port, memory_8_6_port, memory_8_5_port, memory_8_4_port, 
      memory_8_3_port, memory_8_2_port, memory_8_1_port, memory_8_0_port, 
      memory_9_7_port, memory_9_6_port, memory_9_5_port, memory_9_4_port, 
      memory_9_3_port, memory_9_2_port, memory_9_1_port, memory_9_0_port, 
      memory_10_7_port, memory_10_6_port, memory_10_5_port, memory_10_4_port, 
      memory_10_3_port, memory_10_2_port, memory_10_1_port, memory_10_0_port, 
      memory_11_7_port, memory_11_6_port, memory_11_5_port, memory_11_4_port, 
      memory_11_3_port, memory_11_2_port, memory_11_1_port, memory_11_0_port, 
      memory_12_7_port, memory_12_6_port, memory_12_5_port, memory_12_4_port, 
      memory_12_3_port, memory_12_2_port, memory_12_1_port, memory_12_0_port, 
      memory_13_7_port, memory_13_6_port, memory_13_5_port, memory_13_4_port, 
      memory_13_3_port, memory_13_2_port, memory_13_1_port, memory_13_0_port, 
      memory_14_7_port, memory_14_6_port, memory_14_5_port, memory_14_4_port, 
      memory_14_3_port, memory_14_2_port, memory_14_1_port, memory_14_0_port, 
      memory_15_7_port, memory_15_6_port, memory_15_5_port, memory_15_4_port, 
      memory_15_3_port, memory_15_2_port, memory_15_1_port, memory_15_0_port, 
      memory_16_7_port, memory_16_6_port, memory_16_5_port, memory_16_4_port, 
      memory_16_3_port, memory_16_2_port, memory_16_1_port, memory_16_0_port, 
      memory_17_7_port, memory_17_6_port, memory_17_5_port, memory_17_4_port, 
      memory_17_3_port, memory_17_2_port, memory_17_1_port, memory_17_0_port, 
      memory_18_7_port, memory_18_6_port, memory_18_5_port, memory_18_4_port, 
      memory_18_3_port, memory_18_2_port, memory_18_1_port, memory_18_0_port, 
      memory_19_7_port, memory_19_6_port, memory_19_5_port, memory_19_4_port, 
      memory_19_3_port, memory_19_2_port, memory_19_1_port, memory_19_0_port, 
      memory_20_7_port, memory_20_6_port, memory_20_5_port, memory_20_4_port, 
      memory_20_3_port, memory_20_2_port, memory_20_1_port, memory_20_0_port, 
      memory_21_7_port, memory_21_6_port, memory_21_5_port, memory_21_4_port, 
      memory_21_3_port, memory_21_2_port, memory_21_1_port, memory_21_0_port, 
      memory_22_7_port, memory_22_6_port, memory_22_5_port, memory_22_4_port, 
      memory_22_3_port, memory_22_2_port, memory_22_1_port, memory_22_0_port, 
      memory_23_7_port, memory_23_6_port, memory_23_5_port, memory_23_4_port, 
      memory_23_3_port, memory_23_2_port, memory_23_1_port, memory_23_0_port, 
      memory_24_7_port, memory_24_6_port, memory_24_5_port, memory_24_4_port, 
      memory_24_3_port, memory_24_2_port, memory_24_1_port, memory_24_0_port, 
      memory_25_7_port, memory_25_6_port, memory_25_5_port, memory_25_4_port, 
      memory_25_3_port, memory_25_2_port, memory_25_1_port, memory_25_0_port, 
      memory_26_7_port, memory_26_6_port, memory_26_5_port, memory_26_4_port, 
      memory_26_3_port, memory_26_2_port, memory_26_1_port, memory_26_0_port, 
      memory_27_7_port, memory_27_6_port, memory_27_5_port, memory_27_4_port, 
      memory_27_3_port, memory_27_2_port, memory_27_1_port, memory_27_0_port, 
      memory_28_7_port, memory_28_6_port, memory_28_5_port, memory_28_4_port, 
      memory_28_3_port, memory_28_2_port, memory_28_1_port, memory_28_0_port, 
      memory_29_7_port, memory_29_6_port, memory_29_5_port, memory_29_4_port, 
      memory_29_3_port, memory_29_2_port, memory_29_1_port, memory_29_0_port, 
      memory_30_7_port, memory_30_6_port, memory_30_5_port, memory_30_4_port, 
      memory_30_3_port, memory_30_2_port, memory_30_1_port, memory_30_0_port, 
      memory_31_7_port, memory_31_6_port, memory_31_5_port, memory_31_4_port, 
      memory_31_3_port, memory_31_2_port, memory_31_1_port, memory_31_0_port, 
      N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338_port, n339_port, n340_port, n341_port, 
      n342_port, n343_port, n344_port, n345_port, n346_port, n347_port, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
      n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, 
      n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, 
      n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n852, n861, n863, n865, n909, n910, 
      n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, 
      n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, 
      n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, 
      n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, 
      n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, 
      n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, 
      n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, 
      n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, 
      n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, 
      n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, 
      n1026, n1027, n1028, n1029, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, 
      n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, 
      n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, 
      n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, 
      n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
      n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, 
      n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
      n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, 
      n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, 
      n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, 
      n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, 
      n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620 : std_logic;

begin
   DATA <= ( DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, 
      DATA_2_port, DATA_1_port, DATA_0_port );
   OUT_OPCODE <= ( OUT_OPCODE_1_port, OUT_OPCODE_0_port );
   EMPTY <= EMPTY_port;
   FULL <= FULL_port;
   
   X_Logic1_port <= '1';
   state_reg : DFFSR port map( D => X_Logic1_port, CLK => CLK, R => n163, S => 
                           n1603, Q => state);
   readptr_reg_0_inst : DFFSR port map( D => N343, CLK => CLK, R => n163, S => 
                           n1604, Q => readptr_0_port);
   readptr_reg_1_inst : DFFSR port map( D => N344, CLK => CLK, R => n163, S => 
                           n1605, Q => readptr_1_port);
   readptr_reg_3_inst : DFFSR port map( D => N346, CLK => CLK, R => n163, S => 
                           n1606, Q => readptr_3_port);
   writeptr_reg_3_inst : DFFSR port map( D => n1608, CLK => CLK, R => n163, S 
                           => n1609, Q => writeptr_3_port);
   writeptr_reg_0_inst : DFFSR port map( D => n1610, CLK => CLK, R => n163, S 
                           => n1611, Q => writeptr_0_port);
   writeptr_reg_1_inst : DFFSR port map( D => n1612, CLK => CLK, R => n163, S 
                           => n1613, Q => writeptr_1_port);
   writeptr_reg_2_inst : DFFSR port map( D => n1614, CLK => CLK, R => n163, S 
                           => n1615, Q => writeptr_2_port);
   FULL_reg : DFFPOSX1 port map( D => n1431, CLK => CLK, Q => FULL_port);
   BYTE_COUNT_reg_4_inst : DFFSR port map( D => N342, CLK => CLK, R => n163, S 
                           => n1616, Q => BYTE_COUNT(4));
   BYTE_COUNT_reg_3_inst : DFFSR port map( D => N341, CLK => CLK, R => n163, S 
                           => n1617, Q => BYTE_COUNT(3));
   BYTE_COUNT_reg_2_inst : DFFSR port map( D => N340, CLK => CLK, R => n163, S 
                           => n1618, Q => BYTE_COUNT(2));
   BYTE_COUNT_reg_1_inst : DFFSR port map( D => N339, CLK => CLK, R => n163, S 
                           => n1619, Q => BYTE_COUNT(1));
   BYTE_COUNT_reg_0_inst : DFFSR port map( D => N338, CLK => CLK, R => n163, S 
                           => n1620, Q => BYTE_COUNT(0));
   memory_reg_0_7_inst : DFFPOSX1 port map( D => n1406, CLK => CLK, Q => 
                           memory_0_7_port);
   memory_reg_0_6_inst : DFFPOSX1 port map( D => n1405, CLK => CLK, Q => 
                           memory_0_6_port);
   memory_reg_0_5_inst : DFFPOSX1 port map( D => n1404, CLK => CLK, Q => 
                           memory_0_5_port);
   memory_reg_0_4_inst : DFFPOSX1 port map( D => n1403, CLK => CLK, Q => 
                           memory_0_4_port);
   memory_reg_0_3_inst : DFFPOSX1 port map( D => n1402, CLK => CLK, Q => 
                           memory_0_3_port);
   memory_reg_0_2_inst : DFFPOSX1 port map( D => n1401, CLK => CLK, Q => 
                           memory_0_2_port);
   memory_reg_0_1_inst : DFFPOSX1 port map( D => n1400, CLK => CLK, Q => 
                           memory_0_1_port);
   memory_reg_0_0_inst : DFFPOSX1 port map( D => n1399, CLK => CLK, Q => 
                           memory_0_0_port);
   memory_reg_1_7_inst : DFFPOSX1 port map( D => n1414, CLK => CLK, Q => 
                           memory_1_7_port);
   memory_reg_1_6_inst : DFFPOSX1 port map( D => n1413, CLK => CLK, Q => 
                           memory_1_6_port);
   memory_reg_1_5_inst : DFFPOSX1 port map( D => n1412, CLK => CLK, Q => 
                           memory_1_5_port);
   memory_reg_1_4_inst : DFFPOSX1 port map( D => n1411, CLK => CLK, Q => 
                           memory_1_4_port);
   memory_reg_1_3_inst : DFFPOSX1 port map( D => n1410, CLK => CLK, Q => 
                           memory_1_3_port);
   memory_reg_1_2_inst : DFFPOSX1 port map( D => n1409, CLK => CLK, Q => 
                           memory_1_2_port);
   memory_reg_1_1_inst : DFFPOSX1 port map( D => n1408, CLK => CLK, Q => 
                           memory_1_1_port);
   memory_reg_1_0_inst : DFFPOSX1 port map( D => n1407, CLK => CLK, Q => 
                           memory_1_0_port);
   memory_reg_2_7_inst : DFFPOSX1 port map( D => n1422, CLK => CLK, Q => 
                           memory_2_7_port);
   memory_reg_2_6_inst : DFFPOSX1 port map( D => n1421, CLK => CLK, Q => 
                           memory_2_6_port);
   memory_reg_2_5_inst : DFFPOSX1 port map( D => n1420, CLK => CLK, Q => 
                           memory_2_5_port);
   memory_reg_2_4_inst : DFFPOSX1 port map( D => n1419, CLK => CLK, Q => 
                           memory_2_4_port);
   memory_reg_2_3_inst : DFFPOSX1 port map( D => n1418, CLK => CLK, Q => 
                           memory_2_3_port);
   memory_reg_2_2_inst : DFFPOSX1 port map( D => n1417, CLK => CLK, Q => 
                           memory_2_2_port);
   memory_reg_2_1_inst : DFFPOSX1 port map( D => n1416, CLK => CLK, Q => 
                           memory_2_1_port);
   memory_reg_2_0_inst : DFFPOSX1 port map( D => n1415, CLK => CLK, Q => 
                           memory_2_0_port);
   memory_reg_3_7_inst : DFFPOSX1 port map( D => n1430, CLK => CLK, Q => 
                           memory_3_7_port);
   memory_reg_3_6_inst : DFFPOSX1 port map( D => n1429, CLK => CLK, Q => 
                           memory_3_6_port);
   memory_reg_3_5_inst : DFFPOSX1 port map( D => n1428, CLK => CLK, Q => 
                           memory_3_5_port);
   memory_reg_3_4_inst : DFFPOSX1 port map( D => n1427, CLK => CLK, Q => 
                           memory_3_4_port);
   memory_reg_3_3_inst : DFFPOSX1 port map( D => n1426, CLK => CLK, Q => 
                           memory_3_3_port);
   memory_reg_3_2_inst : DFFPOSX1 port map( D => n1425, CLK => CLK, Q => 
                           memory_3_2_port);
   memory_reg_3_1_inst : DFFPOSX1 port map( D => n1424, CLK => CLK, Q => 
                           memory_3_1_port);
   memory_reg_3_0_inst : DFFPOSX1 port map( D => n1423, CLK => CLK, Q => 
                           memory_3_0_port);
   memory_reg_4_7_inst : DFFPOSX1 port map( D => n1602, CLK => CLK, Q => 
                           memory_4_7_port);
   memory_reg_4_6_inst : DFFPOSX1 port map( D => n1601, CLK => CLK, Q => 
                           memory_4_6_port);
   memory_reg_4_5_inst : DFFPOSX1 port map( D => n1600, CLK => CLK, Q => 
                           memory_4_5_port);
   memory_reg_4_4_inst : DFFPOSX1 port map( D => n1599, CLK => CLK, Q => 
                           memory_4_4_port);
   memory_reg_4_3_inst : DFFPOSX1 port map( D => n1598, CLK => CLK, Q => 
                           memory_4_3_port);
   memory_reg_4_2_inst : DFFPOSX1 port map( D => n1597, CLK => CLK, Q => 
                           memory_4_2_port);
   memory_reg_4_1_inst : DFFPOSX1 port map( D => n1596, CLK => CLK, Q => 
                           memory_4_1_port);
   memory_reg_4_0_inst : DFFPOSX1 port map( D => n1595, CLK => CLK, Q => 
                           memory_4_0_port);
   memory_reg_5_7_inst : DFFPOSX1 port map( D => n1592, CLK => CLK, Q => 
                           memory_5_7_port);
   memory_reg_5_6_inst : DFFPOSX1 port map( D => n1591, CLK => CLK, Q => 
                           memory_5_6_port);
   memory_reg_5_5_inst : DFFPOSX1 port map( D => n1590, CLK => CLK, Q => 
                           memory_5_5_port);
   memory_reg_5_4_inst : DFFPOSX1 port map( D => n1589, CLK => CLK, Q => 
                           memory_5_4_port);
   memory_reg_5_3_inst : DFFPOSX1 port map( D => n1588, CLK => CLK, Q => 
                           memory_5_3_port);
   memory_reg_5_2_inst : DFFPOSX1 port map( D => n1587, CLK => CLK, Q => 
                           memory_5_2_port);
   memory_reg_5_1_inst : DFFPOSX1 port map( D => n1586, CLK => CLK, Q => 
                           memory_5_1_port);
   memory_reg_5_0_inst : DFFPOSX1 port map( D => n1585, CLK => CLK, Q => 
                           memory_5_0_port);
   memory_reg_6_7_inst : DFFPOSX1 port map( D => n1582, CLK => CLK, Q => 
                           memory_6_7_port);
   memory_reg_6_6_inst : DFFPOSX1 port map( D => n1581, CLK => CLK, Q => 
                           memory_6_6_port);
   memory_reg_6_5_inst : DFFPOSX1 port map( D => n1580, CLK => CLK, Q => 
                           memory_6_5_port);
   memory_reg_6_4_inst : DFFPOSX1 port map( D => n1579, CLK => CLK, Q => 
                           memory_6_4_port);
   memory_reg_6_3_inst : DFFPOSX1 port map( D => n1578, CLK => CLK, Q => 
                           memory_6_3_port);
   memory_reg_6_2_inst : DFFPOSX1 port map( D => n1577, CLK => CLK, Q => 
                           memory_6_2_port);
   memory_reg_6_1_inst : DFFPOSX1 port map( D => n1576, CLK => CLK, Q => 
                           memory_6_1_port);
   memory_reg_6_0_inst : DFFPOSX1 port map( D => n1575, CLK => CLK, Q => 
                           memory_6_0_port);
   memory_reg_7_7_inst : DFFPOSX1 port map( D => n1572, CLK => CLK, Q => 
                           memory_7_7_port);
   memory_reg_7_6_inst : DFFPOSX1 port map( D => n1571, CLK => CLK, Q => 
                           memory_7_6_port);
   memory_reg_7_5_inst : DFFPOSX1 port map( D => n1570, CLK => CLK, Q => 
                           memory_7_5_port);
   memory_reg_7_4_inst : DFFPOSX1 port map( D => n1569, CLK => CLK, Q => 
                           memory_7_4_port);
   memory_reg_7_3_inst : DFFPOSX1 port map( D => n1568, CLK => CLK, Q => 
                           memory_7_3_port);
   memory_reg_7_2_inst : DFFPOSX1 port map( D => n1567, CLK => CLK, Q => 
                           memory_7_2_port);
   memory_reg_7_1_inst : DFFPOSX1 port map( D => n1566, CLK => CLK, Q => 
                           memory_7_1_port);
   memory_reg_7_0_inst : DFFPOSX1 port map( D => n1565, CLK => CLK, Q => 
                           memory_7_0_port);
   memory_reg_8_7_inst : DFFPOSX1 port map( D => n1433, CLK => CLK, Q => 
                           memory_8_7_port);
   memory_reg_8_6_inst : DFFPOSX1 port map( D => n1434, CLK => CLK, Q => 
                           memory_8_6_port);
   memory_reg_8_5_inst : DFFPOSX1 port map( D => n1435, CLK => CLK, Q => 
                           memory_8_5_port);
   memory_reg_8_4_inst : DFFPOSX1 port map( D => n1436, CLK => CLK, Q => 
                           memory_8_4_port);
   memory_reg_8_3_inst : DFFPOSX1 port map( D => n1437, CLK => CLK, Q => 
                           memory_8_3_port);
   memory_reg_8_2_inst : DFFPOSX1 port map( D => n1438, CLK => CLK, Q => 
                           memory_8_2_port);
   memory_reg_8_1_inst : DFFPOSX1 port map( D => n1439, CLK => CLK, Q => 
                           memory_8_1_port);
   memory_reg_8_0_inst : DFFPOSX1 port map( D => n1440, CLK => CLK, Q => 
                           memory_8_0_port);
   memory_reg_9_7_inst : DFFPOSX1 port map( D => n1441, CLK => CLK, Q => 
                           memory_9_7_port);
   memory_reg_9_6_inst : DFFPOSX1 port map( D => n1442, CLK => CLK, Q => 
                           memory_9_6_port);
   memory_reg_9_5_inst : DFFPOSX1 port map( D => n1443, CLK => CLK, Q => 
                           memory_9_5_port);
   memory_reg_9_4_inst : DFFPOSX1 port map( D => n1444, CLK => CLK, Q => 
                           memory_9_4_port);
   memory_reg_9_3_inst : DFFPOSX1 port map( D => n1445, CLK => CLK, Q => 
                           memory_9_3_port);
   memory_reg_9_2_inst : DFFPOSX1 port map( D => n1446, CLK => CLK, Q => 
                           memory_9_2_port);
   memory_reg_9_1_inst : DFFPOSX1 port map( D => n1447, CLK => CLK, Q => 
                           memory_9_1_port);
   memory_reg_9_0_inst : DFFPOSX1 port map( D => n1448, CLK => CLK, Q => 
                           memory_9_0_port);
   memory_reg_10_7_inst : DFFPOSX1 port map( D => n1449, CLK => CLK, Q => 
                           memory_10_7_port);
   memory_reg_10_6_inst : DFFPOSX1 port map( D => n1450, CLK => CLK, Q => 
                           memory_10_6_port);
   memory_reg_10_5_inst : DFFPOSX1 port map( D => n1451, CLK => CLK, Q => 
                           memory_10_5_port);
   memory_reg_10_4_inst : DFFPOSX1 port map( D => n1452, CLK => CLK, Q => 
                           memory_10_4_port);
   memory_reg_10_3_inst : DFFPOSX1 port map( D => n1453, CLK => CLK, Q => 
                           memory_10_3_port);
   memory_reg_10_2_inst : DFFPOSX1 port map( D => n1454, CLK => CLK, Q => 
                           memory_10_2_port);
   memory_reg_10_1_inst : DFFPOSX1 port map( D => n1455, CLK => CLK, Q => 
                           memory_10_1_port);
   memory_reg_10_0_inst : DFFPOSX1 port map( D => n1456, CLK => CLK, Q => 
                           memory_10_0_port);
   memory_reg_11_7_inst : DFFPOSX1 port map( D => n1457, CLK => CLK, Q => 
                           memory_11_7_port);
   memory_reg_11_6_inst : DFFPOSX1 port map( D => n1458, CLK => CLK, Q => 
                           memory_11_6_port);
   memory_reg_11_5_inst : DFFPOSX1 port map( D => n1459, CLK => CLK, Q => 
                           memory_11_5_port);
   memory_reg_11_4_inst : DFFPOSX1 port map( D => n1460, CLK => CLK, Q => 
                           memory_11_4_port);
   memory_reg_11_3_inst : DFFPOSX1 port map( D => n1461, CLK => CLK, Q => 
                           memory_11_3_port);
   memory_reg_11_2_inst : DFFPOSX1 port map( D => n1462, CLK => CLK, Q => 
                           memory_11_2_port);
   memory_reg_11_1_inst : DFFPOSX1 port map( D => n1463, CLK => CLK, Q => 
                           memory_11_1_port);
   memory_reg_11_0_inst : DFFPOSX1 port map( D => n1464, CLK => CLK, Q => 
                           memory_11_0_port);
   memory_reg_12_7_inst : DFFPOSX1 port map( D => n1391, CLK => CLK, Q => 
                           memory_12_7_port);
   memory_reg_12_6_inst : DFFPOSX1 port map( D => n1392, CLK => CLK, Q => 
                           memory_12_6_port);
   memory_reg_12_5_inst : DFFPOSX1 port map( D => n1393, CLK => CLK, Q => 
                           memory_12_5_port);
   memory_reg_12_4_inst : DFFPOSX1 port map( D => n1394, CLK => CLK, Q => 
                           memory_12_4_port);
   memory_reg_12_3_inst : DFFPOSX1 port map( D => n1395, CLK => CLK, Q => 
                           memory_12_3_port);
   memory_reg_12_2_inst : DFFPOSX1 port map( D => n1396, CLK => CLK, Q => 
                           memory_12_2_port);
   memory_reg_12_1_inst : DFFPOSX1 port map( D => n1397, CLK => CLK, Q => 
                           memory_12_1_port);
   memory_reg_12_0_inst : DFFPOSX1 port map( D => n1398, CLK => CLK, Q => 
                           memory_12_0_port);
   memory_reg_13_7_inst : DFFPOSX1 port map( D => n1383, CLK => CLK, Q => 
                           memory_13_7_port);
   memory_reg_13_6_inst : DFFPOSX1 port map( D => n1384, CLK => CLK, Q => 
                           memory_13_6_port);
   memory_reg_13_5_inst : DFFPOSX1 port map( D => n1385, CLK => CLK, Q => 
                           memory_13_5_port);
   memory_reg_13_4_inst : DFFPOSX1 port map( D => n1386, CLK => CLK, Q => 
                           memory_13_4_port);
   memory_reg_13_3_inst : DFFPOSX1 port map( D => n1387, CLK => CLK, Q => 
                           memory_13_3_port);
   memory_reg_13_2_inst : DFFPOSX1 port map( D => n1388, CLK => CLK, Q => 
                           memory_13_2_port);
   memory_reg_13_1_inst : DFFPOSX1 port map( D => n1389, CLK => CLK, Q => 
                           memory_13_1_port);
   memory_reg_13_0_inst : DFFPOSX1 port map( D => n1390, CLK => CLK, Q => 
                           memory_13_0_port);
   memory_reg_14_7_inst : DFFPOSX1 port map( D => n1375, CLK => CLK, Q => 
                           memory_14_7_port);
   memory_reg_14_6_inst : DFFPOSX1 port map( D => n1376, CLK => CLK, Q => 
                           memory_14_6_port);
   memory_reg_14_5_inst : DFFPOSX1 port map( D => n1377, CLK => CLK, Q => 
                           memory_14_5_port);
   memory_reg_14_4_inst : DFFPOSX1 port map( D => n1378, CLK => CLK, Q => 
                           memory_14_4_port);
   memory_reg_14_3_inst : DFFPOSX1 port map( D => n1379, CLK => CLK, Q => 
                           memory_14_3_port);
   memory_reg_14_2_inst : DFFPOSX1 port map( D => n1380, CLK => CLK, Q => 
                           memory_14_2_port);
   memory_reg_14_1_inst : DFFPOSX1 port map( D => n1381, CLK => CLK, Q => 
                           memory_14_1_port);
   memory_reg_14_0_inst : DFFPOSX1 port map( D => n1382, CLK => CLK, Q => 
                           memory_14_0_port);
   memory_reg_15_7_inst : DFFPOSX1 port map( D => n1367, CLK => CLK, Q => 
                           memory_15_7_port);
   memory_reg_15_6_inst : DFFPOSX1 port map( D => n1368, CLK => CLK, Q => 
                           memory_15_6_port);
   memory_reg_15_5_inst : DFFPOSX1 port map( D => n1369, CLK => CLK, Q => 
                           memory_15_5_port);
   memory_reg_15_4_inst : DFFPOSX1 port map( D => n1370, CLK => CLK, Q => 
                           memory_15_4_port);
   memory_reg_15_3_inst : DFFPOSX1 port map( D => n1371, CLK => CLK, Q => 
                           memory_15_3_port);
   memory_reg_15_2_inst : DFFPOSX1 port map( D => n1372, CLK => CLK, Q => 
                           memory_15_2_port);
   memory_reg_15_1_inst : DFFPOSX1 port map( D => n1373, CLK => CLK, Q => 
                           memory_15_1_port);
   memory_reg_15_0_inst : DFFPOSX1 port map( D => n1374, CLK => CLK, Q => 
                           memory_15_0_port);
   memory_reg_16_7_inst : DFFPOSX1 port map( D => n1465, CLK => CLK, Q => 
                           memory_16_7_port);
   memory_reg_16_6_inst : DFFPOSX1 port map( D => n1466, CLK => CLK, Q => 
                           memory_16_6_port);
   memory_reg_16_5_inst : DFFPOSX1 port map( D => n1467, CLK => CLK, Q => 
                           memory_16_5_port);
   memory_reg_16_4_inst : DFFPOSX1 port map( D => n1468, CLK => CLK, Q => 
                           memory_16_4_port);
   memory_reg_16_3_inst : DFFPOSX1 port map( D => n1469, CLK => CLK, Q => 
                           memory_16_3_port);
   memory_reg_16_2_inst : DFFPOSX1 port map( D => n1470, CLK => CLK, Q => 
                           memory_16_2_port);
   memory_reg_16_1_inst : DFFPOSX1 port map( D => n1471, CLK => CLK, Q => 
                           memory_16_1_port);
   memory_reg_16_0_inst : DFFPOSX1 port map( D => n1472, CLK => CLK, Q => 
                           memory_16_0_port);
   memory_reg_17_7_inst : DFFPOSX1 port map( D => n1473, CLK => CLK, Q => 
                           memory_17_7_port);
   memory_reg_17_6_inst : DFFPOSX1 port map( D => n1474, CLK => CLK, Q => 
                           memory_17_6_port);
   memory_reg_17_5_inst : DFFPOSX1 port map( D => n1475, CLK => CLK, Q => 
                           memory_17_5_port);
   memory_reg_17_4_inst : DFFPOSX1 port map( D => n1476, CLK => CLK, Q => 
                           memory_17_4_port);
   memory_reg_17_3_inst : DFFPOSX1 port map( D => n1477, CLK => CLK, Q => 
                           memory_17_3_port);
   memory_reg_17_2_inst : DFFPOSX1 port map( D => n1478, CLK => CLK, Q => 
                           memory_17_2_port);
   memory_reg_17_1_inst : DFFPOSX1 port map( D => n1479, CLK => CLK, Q => 
                           memory_17_1_port);
   memory_reg_17_0_inst : DFFPOSX1 port map( D => n1480, CLK => CLK, Q => 
                           memory_17_0_port);
   memory_reg_18_7_inst : DFFPOSX1 port map( D => n1481, CLK => CLK, Q => 
                           memory_18_7_port);
   memory_reg_18_6_inst : DFFPOSX1 port map( D => n1482, CLK => CLK, Q => 
                           memory_18_6_port);
   memory_reg_18_5_inst : DFFPOSX1 port map( D => n1483, CLK => CLK, Q => 
                           memory_18_5_port);
   memory_reg_18_4_inst : DFFPOSX1 port map( D => n1484, CLK => CLK, Q => 
                           memory_18_4_port);
   memory_reg_18_3_inst : DFFPOSX1 port map( D => n1485, CLK => CLK, Q => 
                           memory_18_3_port);
   memory_reg_18_2_inst : DFFPOSX1 port map( D => n1486, CLK => CLK, Q => 
                           memory_18_2_port);
   memory_reg_18_1_inst : DFFPOSX1 port map( D => n1487, CLK => CLK, Q => 
                           memory_18_1_port);
   memory_reg_18_0_inst : DFFPOSX1 port map( D => n1488, CLK => CLK, Q => 
                           memory_18_0_port);
   memory_reg_19_7_inst : DFFPOSX1 port map( D => n1489, CLK => CLK, Q => 
                           memory_19_7_port);
   memory_reg_19_6_inst : DFFPOSX1 port map( D => n1490, CLK => CLK, Q => 
                           memory_19_6_port);
   memory_reg_19_5_inst : DFFPOSX1 port map( D => n1491, CLK => CLK, Q => 
                           memory_19_5_port);
   memory_reg_19_4_inst : DFFPOSX1 port map( D => n1492, CLK => CLK, Q => 
                           memory_19_4_port);
   memory_reg_19_3_inst : DFFPOSX1 port map( D => n1493, CLK => CLK, Q => 
                           memory_19_3_port);
   memory_reg_19_2_inst : DFFPOSX1 port map( D => n1494, CLK => CLK, Q => 
                           memory_19_2_port);
   memory_reg_19_1_inst : DFFPOSX1 port map( D => n1495, CLK => CLK, Q => 
                           memory_19_1_port);
   memory_reg_19_0_inst : DFFPOSX1 port map( D => n1496, CLK => CLK, Q => 
                           memory_19_0_port);
   memory_reg_20_7_inst : DFFPOSX1 port map( D => n1359, CLK => CLK, Q => 
                           memory_20_7_port);
   memory_reg_20_6_inst : DFFPOSX1 port map( D => n1360, CLK => CLK, Q => 
                           memory_20_6_port);
   memory_reg_20_5_inst : DFFPOSX1 port map( D => n1361, CLK => CLK, Q => 
                           memory_20_5_port);
   memory_reg_20_4_inst : DFFPOSX1 port map( D => n1362, CLK => CLK, Q => 
                           memory_20_4_port);
   memory_reg_20_3_inst : DFFPOSX1 port map( D => n1363, CLK => CLK, Q => 
                           memory_20_3_port);
   memory_reg_20_2_inst : DFFPOSX1 port map( D => n1364, CLK => CLK, Q => 
                           memory_20_2_port);
   memory_reg_20_1_inst : DFFPOSX1 port map( D => n1365, CLK => CLK, Q => 
                           memory_20_1_port);
   memory_reg_20_0_inst : DFFPOSX1 port map( D => n1366, CLK => CLK, Q => 
                           memory_20_0_port);
   memory_reg_21_7_inst : DFFPOSX1 port map( D => n1351, CLK => CLK, Q => 
                           memory_21_7_port);
   memory_reg_21_6_inst : DFFPOSX1 port map( D => n1352, CLK => CLK, Q => 
                           memory_21_6_port);
   memory_reg_21_5_inst : DFFPOSX1 port map( D => n1353, CLK => CLK, Q => 
                           memory_21_5_port);
   memory_reg_21_4_inst : DFFPOSX1 port map( D => n1354, CLK => CLK, Q => 
                           memory_21_4_port);
   memory_reg_21_3_inst : DFFPOSX1 port map( D => n1355, CLK => CLK, Q => 
                           memory_21_3_port);
   memory_reg_21_2_inst : DFFPOSX1 port map( D => n1356, CLK => CLK, Q => 
                           memory_21_2_port);
   memory_reg_21_1_inst : DFFPOSX1 port map( D => n1357, CLK => CLK, Q => 
                           memory_21_1_port);
   memory_reg_21_0_inst : DFFPOSX1 port map( D => n1358, CLK => CLK, Q => 
                           memory_21_0_port);
   memory_reg_22_7_inst : DFFPOSX1 port map( D => n1343, CLK => CLK, Q => 
                           memory_22_7_port);
   memory_reg_22_6_inst : DFFPOSX1 port map( D => n1344, CLK => CLK, Q => 
                           memory_22_6_port);
   memory_reg_22_5_inst : DFFPOSX1 port map( D => n1345, CLK => CLK, Q => 
                           memory_22_5_port);
   memory_reg_22_4_inst : DFFPOSX1 port map( D => n1346, CLK => CLK, Q => 
                           memory_22_4_port);
   memory_reg_22_3_inst : DFFPOSX1 port map( D => n1347, CLK => CLK, Q => 
                           memory_22_3_port);
   memory_reg_22_2_inst : DFFPOSX1 port map( D => n1348, CLK => CLK, Q => 
                           memory_22_2_port);
   memory_reg_22_1_inst : DFFPOSX1 port map( D => n1349, CLK => CLK, Q => 
                           memory_22_1_port);
   memory_reg_22_0_inst : DFFPOSX1 port map( D => n1350, CLK => CLK, Q => 
                           memory_22_0_port);
   memory_reg_23_7_inst : DFFPOSX1 port map( D => n1335, CLK => CLK, Q => 
                           memory_23_7_port);
   memory_reg_23_6_inst : DFFPOSX1 port map( D => n1336, CLK => CLK, Q => 
                           memory_23_6_port);
   memory_reg_23_5_inst : DFFPOSX1 port map( D => n1337, CLK => CLK, Q => 
                           memory_23_5_port);
   memory_reg_23_4_inst : DFFPOSX1 port map( D => n1338, CLK => CLK, Q => 
                           memory_23_4_port);
   memory_reg_23_3_inst : DFFPOSX1 port map( D => n1339, CLK => CLK, Q => 
                           memory_23_3_port);
   memory_reg_23_2_inst : DFFPOSX1 port map( D => n1340, CLK => CLK, Q => 
                           memory_23_2_port);
   memory_reg_23_1_inst : DFFPOSX1 port map( D => n1341, CLK => CLK, Q => 
                           memory_23_1_port);
   memory_reg_23_0_inst : DFFPOSX1 port map( D => n1342, CLK => CLK, Q => 
                           memory_23_0_port);
   memory_reg_24_7_inst : DFFPOSX1 port map( D => n1327, CLK => CLK, Q => 
                           memory_24_7_port);
   memory_reg_24_6_inst : DFFPOSX1 port map( D => n1328, CLK => CLK, Q => 
                           memory_24_6_port);
   memory_reg_24_5_inst : DFFPOSX1 port map( D => n1329, CLK => CLK, Q => 
                           memory_24_5_port);
   memory_reg_24_4_inst : DFFPOSX1 port map( D => n1330, CLK => CLK, Q => 
                           memory_24_4_port);
   memory_reg_24_3_inst : DFFPOSX1 port map( D => n1331, CLK => CLK, Q => 
                           memory_24_3_port);
   memory_reg_24_2_inst : DFFPOSX1 port map( D => n1332, CLK => CLK, Q => 
                           memory_24_2_port);
   memory_reg_24_1_inst : DFFPOSX1 port map( D => n1333, CLK => CLK, Q => 
                           memory_24_1_port);
   memory_reg_24_0_inst : DFFPOSX1 port map( D => n1334, CLK => CLK, Q => 
                           memory_24_0_port);
   memory_reg_25_7_inst : DFFPOSX1 port map( D => n1319, CLK => CLK, Q => 
                           memory_25_7_port);
   memory_reg_25_6_inst : DFFPOSX1 port map( D => n1320, CLK => CLK, Q => 
                           memory_25_6_port);
   memory_reg_25_5_inst : DFFPOSX1 port map( D => n1321, CLK => CLK, Q => 
                           memory_25_5_port);
   memory_reg_25_4_inst : DFFPOSX1 port map( D => n1322, CLK => CLK, Q => 
                           memory_25_4_port);
   memory_reg_25_3_inst : DFFPOSX1 port map( D => n1323, CLK => CLK, Q => 
                           memory_25_3_port);
   memory_reg_25_2_inst : DFFPOSX1 port map( D => n1324, CLK => CLK, Q => 
                           memory_25_2_port);
   memory_reg_25_1_inst : DFFPOSX1 port map( D => n1325, CLK => CLK, Q => 
                           memory_25_1_port);
   memory_reg_25_0_inst : DFFPOSX1 port map( D => n1326, CLK => CLK, Q => 
                           memory_25_0_port);
   memory_reg_26_7_inst : DFFPOSX1 port map( D => n1311, CLK => CLK, Q => 
                           memory_26_7_port);
   memory_reg_26_6_inst : DFFPOSX1 port map( D => n1312, CLK => CLK, Q => 
                           memory_26_6_port);
   memory_reg_26_5_inst : DFFPOSX1 port map( D => n1313, CLK => CLK, Q => 
                           memory_26_5_port);
   memory_reg_26_4_inst : DFFPOSX1 port map( D => n1314, CLK => CLK, Q => 
                           memory_26_4_port);
   memory_reg_26_3_inst : DFFPOSX1 port map( D => n1315, CLK => CLK, Q => 
                           memory_26_3_port);
   memory_reg_26_2_inst : DFFPOSX1 port map( D => n1316, CLK => CLK, Q => 
                           memory_26_2_port);
   memory_reg_26_1_inst : DFFPOSX1 port map( D => n1317, CLK => CLK, Q => 
                           memory_26_1_port);
   memory_reg_26_0_inst : DFFPOSX1 port map( D => n1318, CLK => CLK, Q => 
                           memory_26_0_port);
   memory_reg_27_7_inst : DFFPOSX1 port map( D => n1303, CLK => CLK, Q => 
                           memory_27_7_port);
   memory_reg_27_6_inst : DFFPOSX1 port map( D => n1304, CLK => CLK, Q => 
                           memory_27_6_port);
   memory_reg_27_5_inst : DFFPOSX1 port map( D => n1305, CLK => CLK, Q => 
                           memory_27_5_port);
   memory_reg_27_4_inst : DFFPOSX1 port map( D => n1306, CLK => CLK, Q => 
                           memory_27_4_port);
   memory_reg_27_3_inst : DFFPOSX1 port map( D => n1307, CLK => CLK, Q => 
                           memory_27_3_port);
   memory_reg_27_2_inst : DFFPOSX1 port map( D => n1308, CLK => CLK, Q => 
                           memory_27_2_port);
   memory_reg_27_1_inst : DFFPOSX1 port map( D => n1309, CLK => CLK, Q => 
                           memory_27_1_port);
   memory_reg_27_0_inst : DFFPOSX1 port map( D => n1310, CLK => CLK, Q => 
                           memory_27_0_port);
   memory_reg_28_7_inst : DFFPOSX1 port map( D => n1497, CLK => CLK, Q => 
                           memory_28_7_port);
   memory_reg_28_6_inst : DFFPOSX1 port map( D => n1498, CLK => CLK, Q => 
                           memory_28_6_port);
   memory_reg_28_5_inst : DFFPOSX1 port map( D => n1499, CLK => CLK, Q => 
                           memory_28_5_port);
   memory_reg_28_4_inst : DFFPOSX1 port map( D => n1500, CLK => CLK, Q => 
                           memory_28_4_port);
   memory_reg_28_3_inst : DFFPOSX1 port map( D => n1501, CLK => CLK, Q => 
                           memory_28_3_port);
   memory_reg_28_2_inst : DFFPOSX1 port map( D => n1502, CLK => CLK, Q => 
                           memory_28_2_port);
   memory_reg_28_1_inst : DFFPOSX1 port map( D => n1503, CLK => CLK, Q => 
                           memory_28_1_port);
   memory_reg_28_0_inst : DFFPOSX1 port map( D => n1504, CLK => CLK, Q => 
                           memory_28_0_port);
   memory_reg_29_7_inst : DFFPOSX1 port map( D => n1505, CLK => CLK, Q => 
                           memory_29_7_port);
   memory_reg_29_6_inst : DFFPOSX1 port map( D => n1506, CLK => CLK, Q => 
                           memory_29_6_port);
   memory_reg_29_5_inst : DFFPOSX1 port map( D => n1507, CLK => CLK, Q => 
                           memory_29_5_port);
   memory_reg_29_4_inst : DFFPOSX1 port map( D => n1508, CLK => CLK, Q => 
                           memory_29_4_port);
   memory_reg_29_3_inst : DFFPOSX1 port map( D => n1509, CLK => CLK, Q => 
                           memory_29_3_port);
   memory_reg_29_2_inst : DFFPOSX1 port map( D => n1510, CLK => CLK, Q => 
                           memory_29_2_port);
   memory_reg_29_1_inst : DFFPOSX1 port map( D => n1511, CLK => CLK, Q => 
                           memory_29_1_port);
   memory_reg_29_0_inst : DFFPOSX1 port map( D => n1512, CLK => CLK, Q => 
                           memory_29_0_port);
   memory_reg_30_7_inst : DFFPOSX1 port map( D => n1513, CLK => CLK, Q => 
                           memory_30_7_port);
   memory_reg_30_6_inst : DFFPOSX1 port map( D => n1514, CLK => CLK, Q => 
                           memory_30_6_port);
   memory_reg_30_5_inst : DFFPOSX1 port map( D => n1515, CLK => CLK, Q => 
                           memory_30_5_port);
   memory_reg_30_4_inst : DFFPOSX1 port map( D => n1516, CLK => CLK, Q => 
                           memory_30_4_port);
   memory_reg_30_3_inst : DFFPOSX1 port map( D => n1517, CLK => CLK, Q => 
                           memory_30_3_port);
   memory_reg_30_2_inst : DFFPOSX1 port map( D => n1518, CLK => CLK, Q => 
                           memory_30_2_port);
   memory_reg_30_1_inst : DFFPOSX1 port map( D => n1519, CLK => CLK, Q => 
                           memory_30_1_port);
   memory_reg_30_0_inst : DFFPOSX1 port map( D => n1520, CLK => CLK, Q => 
                           memory_30_0_port);
   memory_reg_31_7_inst : DFFPOSX1 port map( D => n1521, CLK => CLK, Q => 
                           memory_31_7_port);
   memory_reg_31_6_inst : DFFPOSX1 port map( D => n1522, CLK => CLK, Q => 
                           memory_31_6_port);
   memory_reg_31_5_inst : DFFPOSX1 port map( D => n1523, CLK => CLK, Q => 
                           memory_31_5_port);
   memory_reg_31_4_inst : DFFPOSX1 port map( D => n1524, CLK => CLK, Q => 
                           memory_31_4_port);
   memory_reg_31_3_inst : DFFPOSX1 port map( D => n1525, CLK => CLK, Q => 
                           memory_31_3_port);
   memory_reg_31_2_inst : DFFPOSX1 port map( D => n1526, CLK => CLK, Q => 
                           memory_31_2_port);
   memory_reg_31_1_inst : DFFPOSX1 port map( D => n1527, CLK => CLK, Q => 
                           memory_31_1_port);
   memory_reg_31_0_inst : DFFPOSX1 port map( D => n1528, CLK => CLK, Q => 
                           memory_31_0_port);
   opcode_reg_0_1_inst : DFFPOSX1 port map( D => n1296, CLK => CLK, Q => 
                           opcode_0_1_port);
   opcode_reg_0_0_inst : DFFPOSX1 port map( D => n1295, CLK => CLK, Q => 
                           opcode_0_0_port);
   opcode_reg_1_1_inst : DFFPOSX1 port map( D => n1298, CLK => CLK, Q => 
                           opcode_1_1_port);
   opcode_reg_1_0_inst : DFFPOSX1 port map( D => n1297, CLK => CLK, Q => 
                           opcode_1_0_port);
   opcode_reg_2_1_inst : DFFPOSX1 port map( D => n1300, CLK => CLK, Q => 
                           opcode_2_1_port);
   opcode_reg_2_0_inst : DFFPOSX1 port map( D => n1299, CLK => CLK, Q => 
                           opcode_2_0_port);
   opcode_reg_3_1_inst : DFFPOSX1 port map( D => n1302, CLK => CLK, Q => 
                           opcode_3_1_port);
   opcode_reg_3_0_inst : DFFPOSX1 port map( D => n1301, CLK => CLK, Q => 
                           opcode_3_0_port);
   opcode_reg_4_1_inst : DFFPOSX1 port map( D => n1594, CLK => CLK, Q => 
                           opcode_4_1_port);
   opcode_reg_4_0_inst : DFFPOSX1 port map( D => n1593, CLK => CLK, Q => 
                           opcode_4_0_port);
   opcode_reg_5_1_inst : DFFPOSX1 port map( D => n1584, CLK => CLK, Q => 
                           opcode_5_1_port);
   opcode_reg_5_0_inst : DFFPOSX1 port map( D => n1583, CLK => CLK, Q => 
                           opcode_5_0_port);
   opcode_reg_6_1_inst : DFFPOSX1 port map( D => n1574, CLK => CLK, Q => 
                           opcode_6_1_port);
   opcode_reg_6_0_inst : DFFPOSX1 port map( D => n1573, CLK => CLK, Q => 
                           opcode_6_0_port);
   opcode_reg_7_1_inst : DFFPOSX1 port map( D => n1564, CLK => CLK, Q => 
                           opcode_7_1_port);
   opcode_reg_7_0_inst : DFFPOSX1 port map( D => n1563, CLK => CLK, Q => 
                           opcode_7_0_port);
   opcode_reg_8_1_inst : DFFPOSX1 port map( D => n1529, CLK => CLK, Q => 
                           opcode_8_1_port);
   opcode_reg_8_0_inst : DFFPOSX1 port map( D => n1530, CLK => CLK, Q => 
                           opcode_8_0_port);
   opcode_reg_9_1_inst : DFFPOSX1 port map( D => n1531, CLK => CLK, Q => 
                           opcode_9_1_port);
   opcode_reg_9_0_inst : DFFPOSX1 port map( D => n1532, CLK => CLK, Q => 
                           opcode_9_0_port);
   opcode_reg_10_1_inst : DFFPOSX1 port map( D => n1533, CLK => CLK, Q => 
                           opcode_10_1_port);
   opcode_reg_10_0_inst : DFFPOSX1 port map( D => n1534, CLK => CLK, Q => 
                           opcode_10_0_port);
   opcode_reg_11_1_inst : DFFPOSX1 port map( D => n1535, CLK => CLK, Q => 
                           opcode_11_1_port);
   opcode_reg_11_0_inst : DFFPOSX1 port map( D => n1536, CLK => CLK, Q => 
                           opcode_11_0_port);
   opcode_reg_12_1_inst : DFFPOSX1 port map( D => n1293, CLK => CLK, Q => 
                           opcode_12_1_port);
   opcode_reg_12_0_inst : DFFPOSX1 port map( D => n1294, CLK => CLK, Q => 
                           opcode_12_0_port);
   opcode_reg_13_1_inst : DFFPOSX1 port map( D => n1291, CLK => CLK, Q => 
                           opcode_13_1_port);
   opcode_reg_13_0_inst : DFFPOSX1 port map( D => n1292, CLK => CLK, Q => 
                           opcode_13_0_port);
   opcode_reg_14_1_inst : DFFPOSX1 port map( D => n1289, CLK => CLK, Q => 
                           opcode_14_1_port);
   opcode_reg_14_0_inst : DFFPOSX1 port map( D => n1290, CLK => CLK, Q => 
                           opcode_14_0_port);
   opcode_reg_15_1_inst : DFFPOSX1 port map( D => n1287, CLK => CLK, Q => 
                           opcode_15_1_port);
   opcode_reg_15_0_inst : DFFPOSX1 port map( D => n1288, CLK => CLK, Q => 
                           opcode_15_0_port);
   opcode_reg_16_1_inst : DFFPOSX1 port map( D => n1537, CLK => CLK, Q => 
                           opcode_16_1_port);
   opcode_reg_16_0_inst : DFFPOSX1 port map( D => n1538, CLK => CLK, Q => 
                           opcode_16_0_port);
   opcode_reg_17_1_inst : DFFPOSX1 port map( D => n1539, CLK => CLK, Q => 
                           opcode_17_1_port);
   opcode_reg_17_0_inst : DFFPOSX1 port map( D => n1540, CLK => CLK, Q => 
                           opcode_17_0_port);
   opcode_reg_18_1_inst : DFFPOSX1 port map( D => n1541, CLK => CLK, Q => 
                           opcode_18_1_port);
   opcode_reg_18_0_inst : DFFPOSX1 port map( D => n1542, CLK => CLK, Q => 
                           opcode_18_0_port);
   opcode_reg_19_1_inst : DFFPOSX1 port map( D => n1543, CLK => CLK, Q => 
                           opcode_19_1_port);
   opcode_reg_19_0_inst : DFFPOSX1 port map( D => n1544, CLK => CLK, Q => 
                           opcode_19_0_port);
   opcode_reg_20_1_inst : DFFPOSX1 port map( D => n1285, CLK => CLK, Q => 
                           opcode_20_1_port);
   opcode_reg_20_0_inst : DFFPOSX1 port map( D => n1286, CLK => CLK, Q => 
                           opcode_20_0_port);
   opcode_reg_21_1_inst : DFFPOSX1 port map( D => n1283, CLK => CLK, Q => 
                           opcode_21_1_port);
   opcode_reg_21_0_inst : DFFPOSX1 port map( D => n1284, CLK => CLK, Q => 
                           opcode_21_0_port);
   opcode_reg_22_1_inst : DFFPOSX1 port map( D => n1281, CLK => CLK, Q => 
                           opcode_22_1_port);
   opcode_reg_22_0_inst : DFFPOSX1 port map( D => n1282, CLK => CLK, Q => 
                           opcode_22_0_port);
   opcode_reg_23_1_inst : DFFPOSX1 port map( D => n1279, CLK => CLK, Q => 
                           opcode_23_1_port);
   opcode_reg_23_0_inst : DFFPOSX1 port map( D => n1280, CLK => CLK, Q => 
                           opcode_23_0_port);
   opcode_reg_24_1_inst : DFFPOSX1 port map( D => n1277, CLK => CLK, Q => 
                           opcode_24_1_port);
   opcode_reg_24_0_inst : DFFPOSX1 port map( D => n1278, CLK => CLK, Q => 
                           opcode_24_0_port);
   opcode_reg_25_1_inst : DFFPOSX1 port map( D => n1275, CLK => CLK, Q => 
                           opcode_25_1_port);
   opcode_reg_25_0_inst : DFFPOSX1 port map( D => n1276, CLK => CLK, Q => 
                           opcode_25_0_port);
   opcode_reg_26_1_inst : DFFPOSX1 port map( D => n1273, CLK => CLK, Q => 
                           opcode_26_1_port);
   opcode_reg_26_0_inst : DFFPOSX1 port map( D => n1274, CLK => CLK, Q => 
                           opcode_26_0_port);
   opcode_reg_27_1_inst : DFFPOSX1 port map( D => n1271, CLK => CLK, Q => 
                           opcode_27_1_port);
   opcode_reg_27_0_inst : DFFPOSX1 port map( D => n1272, CLK => CLK, Q => 
                           opcode_27_0_port);
   opcode_reg_28_1_inst : DFFPOSX1 port map( D => n1545, CLK => CLK, Q => 
                           opcode_28_1_port);
   opcode_reg_28_0_inst : DFFPOSX1 port map( D => n1546, CLK => CLK, Q => 
                           opcode_28_0_port);
   opcode_reg_29_1_inst : DFFPOSX1 port map( D => n1547, CLK => CLK, Q => 
                           opcode_29_1_port);
   opcode_reg_29_0_inst : DFFPOSX1 port map( D => n1548, CLK => CLK, Q => 
                           opcode_29_0_port);
   opcode_reg_30_1_inst : DFFPOSX1 port map( D => n1549, CLK => CLK, Q => 
                           opcode_30_1_port);
   opcode_reg_30_0_inst : DFFPOSX1 port map( D => n1550, CLK => CLK, Q => 
                           opcode_30_0_port);
   opcode_reg_31_1_inst : DFFPOSX1 port map( D => n1551, CLK => CLK, Q => 
                           opcode_31_1_port);
   opcode_reg_31_0_inst : DFFPOSX1 port map( D => n1552, CLK => CLK, Q => 
                           opcode_31_0_port);
   DATA_reg_7_inst : DFFPOSX1 port map( D => n1553, CLK => CLK, Q => 
                           DATA_7_port);
   DATA_reg_6_inst : DFFPOSX1 port map( D => n1554, CLK => CLK, Q => 
                           DATA_6_port);
   DATA_reg_5_inst : DFFPOSX1 port map( D => n1555, CLK => CLK, Q => 
                           DATA_5_port);
   DATA_reg_4_inst : DFFPOSX1 port map( D => n1556, CLK => CLK, Q => 
                           DATA_4_port);
   DATA_reg_3_inst : DFFPOSX1 port map( D => n1557, CLK => CLK, Q => 
                           DATA_3_port);
   DATA_reg_2_inst : DFFPOSX1 port map( D => n1558, CLK => CLK, Q => 
                           DATA_2_port);
   DATA_reg_1_inst : DFFPOSX1 port map( D => n1559, CLK => CLK, Q => 
                           DATA_1_port);
   DATA_reg_0_inst : DFFPOSX1 port map( D => n1560, CLK => CLK, Q => 
                           DATA_0_port);
   OUT_OPCODE_reg_1_inst : DFFPOSX1 port map( D => n1561, CLK => CLK, Q => 
                           OUT_OPCODE_1_port);
   OUT_OPCODE_reg_0_inst : DFFPOSX1 port map( D => n1562, CLK => CLK, Q => 
                           OUT_OPCODE_0_port);
   EMPTY_reg : DFFPOSX1 port map( D => n1432, CLK => CLK, Q => EMPTY_port);
   n1620 <= '1';
   n1619 <= '1';
   n1618 <= '1';
   n1617 <= '1';
   n1616 <= '1';
   n1615 <= '1';
   n1613 <= '1';
   n1611 <= '1';
   n1609 <= '1';
   n1606 <= '1';
   n1605 <= '1';
   n1604 <= '1';
   n1603 <= '1';
   readptr_reg_2_inst : DFFSR port map( D => N345, CLK => CLK, R => n163, S => 
                           n21, Q => readptr_2_port);
   readptr_reg_4_inst : DFFSR port map( D => N347, CLK => CLK, R => n163, S => 
                           n20, Q => readptr_4_port);
   writeptr_reg_4_inst : DFFSR port map( D => n1607, CLK => CLK, R => n163, S 
                           => n19, Q => writeptr_4_port);
   U3 : INVX2 port map( A => n17, Y => n127);
   U4 : INVX2 port map( A => writeptr_0_port, Y => n132);
   U5 : INVX1 port map( A => n88, Y => n40);
   U6 : XOR2X1 port map( A => n46, B => n134, Y => n575);
   U7 : INVX2 port map( A => n46, Y => n131);
   U8 : XNOR2X1 port map( A => n101, B => n135, Y => n82);
   U9 : INVX4 port map( A => n135, Y => n136);
   U10 : INVX2 port map( A => n534, Y => n542);
   U11 : NAND2X1 port map( A => RCV_OPCODE(1), B => RCV_OPCODE(0), Y => n1);
   U12 : NAND2X1 port map( A => RCV_OPCODE(1), B => RCV_OPCODE(0), Y => n2);
   U13 : INVX2 port map( A => n1, Y => n3);
   U14 : NAND2X1 port map( A => n2, B => n230, Y => n4);
   U15 : NAND2X1 port map( A => n1, B => n241, Y => n5);
   U16 : AND2X2 port map( A => n209, B => n218, Y => n6);
   U17 : INVX1 port map( A => n331, Y => n115);
   U18 : AND2X2 port map( A => n1237, B => n1247, Y => n7);
   U19 : AND2X2 port map( A => n1267, B => n1237, Y => n8);
   U20 : AND2X1 port map( A => n1258, B => n1237, Y => n9);
   U21 : AND2X2 port map( A => n1267, B => n86, Y => n10);
   U22 : AND2X1 port map( A => n1237, B => n1248, Y => n11);
   U23 : AND2X1 port map( A => n1238, B => n1237, Y => n12);
   U24 : AND2X1 port map( A => n1238, B => n86, Y => n13);
   U25 : AND2X1 port map( A => n1248, B => n86, Y => n14);
   U26 : AND2X1 port map( A => n1259, B => n86, Y => n15);
   U27 : AND2X2 port map( A => n1259, B => n1237, Y => n16);
   U28 : AND2X2 port map( A => n1268, B => n1237, Y => n17);
   U29 : AND2X2 port map( A => n1268, B => n86, Y => n18);
   U30 : INVX1 port map( A => RCV_DATA(5), Y => n540);
   U31 : INVX1 port map( A => RCV_DATA(0), Y => n535);
   U32 : INVX1 port map( A => RCV_DATA(2), Y => n537);
   U33 : INVX1 port map( A => RCV_DATA(3), Y => n538);
   U34 : INVX1 port map( A => RCV_DATA(4), Y => n539);
   n19 <= '1';
   n20 <= '1';
   n21 <= '1';
   U38 : NAND2X1 port map( A => n227, B => n161, Y => n22);
   U39 : NAND2X1 port map( A => n251, B => n161, Y => n23);
   U40 : NAND3X1 port map( A => n66, B => n64, C => n191, Y => n24);
   U41 : INVX1 port map( A => RCV_DATA(1), Y => n536);
   U42 : NAND2X1 port map( A => readptr_0_port, B => n219, Y => n25);
   U43 : INVX2 port map( A => n134, Y => n219);
   U44 : NAND2X1 port map( A => n293, B => n161, Y => n26);
   U45 : INVX2 port map( A => n247, Y => n249);
   U46 : NAND2X1 port map( A => n276, B => n160, Y => n27);
   U47 : INVX1 port map( A => RCV_DATA(6), Y => n541);
   U48 : INVX1 port map( A => n575, Y => n576);
   U49 : OR2X1 port map( A => n132, B => n129, Y => n28);
   U50 : XNOR2X1 port map( A => n569, B => n51, Y => n64);
   U51 : INVX2 port map( A => n618, Y => n51);
   U52 : BUFX2 port map( A => n67, Y => n29);
   U53 : NAND2X1 port map( A => n261, B => n160, Y => n30);
   U54 : NAND3X1 port map( A => n70, B => n134, C => n130, Y => n31);
   U55 : INVX2 port map( A => n322, Y => n323);
   U56 : NAND2X1 port map( A => n160, B => n296, Y => n32);
   U57 : NAND2X1 port map( A => n265, B => n161, Y => n33);
   U58 : NOR2X1 port map( A => n614, B => n57, Y => n34);
   U59 : INVX1 port map( A => n34, Y => n612);
   U60 : NAND2X1 port map( A => n193, B => n160, Y => n35);
   U61 : NAND2X1 port map( A => n160, B => n220, Y => n36);
   U62 : NAND2X1 port map( A => n161, B => n210, Y => n37);
   U63 : NAND2X1 port map( A => n160, B => n246, Y => n38);
   U64 : NAND2X1 port map( A => n161, B => n254, Y => n39);
   U65 : INVX8 port map( A => n128, Y => n70);
   U66 : INVX2 port map( A => n297, Y => n298);
   U67 : AND2X2 port map( A => n40, B => n41, Y => n166);
   U68 : INVX1 port map( A => n41, Y => n543);
   U69 : INVX2 port map( A => n266, Y => n268);
   U70 : MUX2X1 port map( B => n116, A => n321, S => n3, Y => n287);
   U71 : INVX4 port map( A => n480, Y => n481);
   U72 : INVX4 port map( A => n448, Y => n456);
   U73 : AND2X2 port map( A => n545, B => n164, Y => n41);
   U74 : NAND2X1 port map( A => n83, B => W_ENABLE, Y => n42);
   U75 : INVX8 port map( A => n162, Y => n161);
   U76 : BUFX4 port map( A => readptr_2_port, Y => n43);
   U77 : INVX1 port map( A => n189, Y => n44);
   U78 : INVX2 port map( A => n44, Y => n45);
   U79 : INVX4 port map( A => n488, Y => n496);
   U80 : INVX4 port map( A => n528, Y => n529);
   U81 : INVX4 port map( A => n518, Y => n526);
   U82 : INVX4 port map( A => n530, Y => n531);
   U83 : INVX1 port map( A => writeptr_1_port, Y => n46);
   U84 : INVX8 port map( A => n132, Y => n134);
   U85 : INVX4 port map( A => n508, Y => n516);
   U86 : INVX4 port map( A => n532, Y => n533);
   U87 : INVX1 port map( A => RCV_OPCODE(1), Y => n341_port);
   U88 : AND2X2 port map( A => n49, B => n618, Y => n86);
   U89 : AND2X2 port map( A => n49, B => n43, Y => n87);
   U90 : OR2X2 port map( A => n68, B => n42, Y => n47);
   U91 : BUFX2 port map( A => n592, Y => n48);
   U92 : BUFX4 port map( A => readptr_1_port, Y => n49);
   U93 : INVX4 port map( A => n57, Y => n50);
   U94 : INVX2 port map( A => readptr_0_port, Y => n57);
   U95 : INVX2 port map( A => n115, Y => n116);
   U96 : INVX4 port map( A => n568, Y => n162);
   U97 : BUFX2 port map( A => writeptr_4_port, Y => n52);
   U98 : INVX1 port map( A => n31, Y => n117);
   U99 : INVX2 port map( A => n620, Y => n53);
   U100 : INVX2 port map( A => readptr_4_port, Y => n620);
   U101 : NAND2X1 port map( A => n116, B => n45, Y => n54);
   U102 : NAND2X1 port map( A => W_ENABLE, B => n83, Y => n55);
   U103 : BUFX2 port map( A => n29, Y => n56);
   U104 : INVX1 port map( A => readptr_0_port, Y => n617);
   U105 : INVX2 port map( A => n226, Y => n58);
   U106 : INVX4 port map( A => n58, Y => n59);
   U107 : INVX2 port map( A => n260, Y => n60);
   U108 : INVX4 port map( A => n60, Y => n61);
   U109 : AND2X2 port map( A => n52, B => n264, Y => n89);
   U110 : AND2X2 port map( A => n52, B => n73, Y => n90);
   U111 : INVX1 port map( A => writeptr_4_port, Y => n591);
   U112 : INVX4 port map( A => n498, Y => n506);
   U113 : NAND2X1 port map( A => n160, B => n290, Y => n62);
   U114 : NOR2X1 port map( A => n129, B => n132, Y => n63);
   U115 : INVX2 port map( A => writeptr_1_port, Y => n129);
   U116 : INVX1 port map( A => n64, Y => n561);
   U117 : NAND2X1 port map( A => n161, B => n281, Y => n65);
   U118 : BUFX4 port map( A => n305, Y => n91);
   U119 : BUFX4 port map( A => n305, Y => n92);
   U120 : BUFX4 port map( A => n236, Y => n94);
   U121 : BUFX4 port map( A => n336, Y => n96);
   U122 : BUFX4 port map( A => n271, Y => n98);
   U123 : INVX4 port map( A => n32, Y => n487);
   U124 : INVX1 port map( A => n67, Y => n579);
   U125 : INVX4 port map( A => n30, Y => n437);
   U126 : INVX4 port map( A => n23, Y => n431);
   U127 : INVX4 port map( A => n390, Y => n398);
   U128 : INVX4 port map( A => n22, Y => n389);
   U129 : NOR2X1 port map( A => n41, B => n190, Y => n66);
   U130 : INVX4 port map( A => n382, Y => n383);
   U131 : INVX4 port map( A => n70, Y => n218);
   U132 : INVX4 port map( A => n35, Y => n350);
   U133 : INVX4 port map( A => n38, Y => n428);
   U134 : INVX4 port map( A => n37, Y => n380);
   U135 : INVX4 port map( A => n39, Y => n433);
   U136 : INVX4 port map( A => n36, Y => n385);
   U137 : INVX4 port map( A => n434, Y => n435);
   U138 : INVX4 port map( A => n386, Y => n387);
   U139 : INVX4 port map( A => n410, Y => n418);
   U140 : INVX4 port map( A => n362, Y => n370);
   U141 : INVX4 port map( A => n400, Y => n408);
   U142 : INVX4 port map( A => n352, Y => n360);
   U143 : INVX4 port map( A => n65, Y => n476);
   U144 : INVX2 port map( A => n24, Y => n68);
   U145 : INVX4 port map( A => n27, Y => n466);
   U146 : INVX4 port map( A => n26, Y => n485);
   U147 : INVX4 port map( A => n62, Y => n483);
   U148 : INVX4 port map( A => n33, Y => n446);
   U149 : AND2X2 port map( A => n24, B => W_ENABLE, Y => n67);
   U150 : OR2X1 port map( A => n316, B => n55, Y => n69);
   U151 : OR2X2 port map( A => n68, B => n71, Y => n478);
   U152 : NAND2X1 port map( A => n83, B => W_ENABLE, Y => n71);
   U153 : INVX1 port map( A => n478, Y => n479);
   U154 : INVX8 port map( A => n162, Y => n160);
   U155 : INVX2 port map( A => n14, Y => n105);
   U156 : INVX2 port map( A => n341_port, Y => n143);
   U157 : INVX2 port map( A => n11, Y => n123);
   U158 : INVX2 port map( A => n9, Y => n124);
   U159 : INVX1 port map( A => n802, Y => n106);
   U160 : INVX2 port map( A => n13, Y => n102);
   U161 : INVX2 port map( A => n15, Y => n108);
   U162 : INVX2 port map( A => n139, Y => n137);
   U163 : INVX2 port map( A => n139, Y => n138);
   U164 : INVX2 port map( A => n339_port, Y => n139);
   U165 : INVX2 port map( A => n143, Y => n140);
   U166 : INVX2 port map( A => n143, Y => n141);
   U167 : BUFX2 port map( A => n336, Y => n95);
   U168 : INVX2 port map( A => n143, Y => n142);
   U169 : AND2X2 port map( A => RCV_OPCODE(0), B => RCV_OPCODE(1), Y => n72);
   U170 : BUFX2 port map( A => n271, Y => n97);
   U171 : BUFX2 port map( A => n236, Y => n93);
   U172 : INVX2 port map( A => n6, Y => n118);
   U173 : NOR2X1 port map( A => RST, B => n100, Y => n73);
   U174 : INVX2 port map( A => RST, Y => n163);
   U175 : AND2X2 port map( A => n1268, B => n87, Y => n74);
   U176 : AND2X2 port map( A => n1238, B => n87, Y => n75);
   U177 : AND2X2 port map( A => n1259, B => n87, Y => n76);
   U178 : AND2X2 port map( A => n1248, B => n87, Y => n77);
   U179 : AND2X2 port map( A => n1267, B => n87, Y => n78);
   U180 : AND2X2 port map( A => n1236, B => n87, Y => n79);
   U181 : AND2X2 port map( A => n1247, B => n87, Y => n80);
   U182 : AND2X2 port map( A => n1258, B => n87, Y => n81);
   U183 : XOR2X1 port map( A => n586, B => n82, Y => n562);
   U184 : XNOR2X1 port map( A => n592, B => n558, Y => n563);
   U185 : INVX1 port map( A => n219, Y => n133);
   U186 : INVX2 port map( A => n7, Y => n122);
   U187 : INVX4 port map( A => n8, Y => n126);
   U188 : INVX2 port map( A => n119, Y => n120);
   U189 : INVX1 port map( A => n793, Y => n119);
   U190 : INVX4 port map( A => n16, Y => n125);
   U191 : INVX2 port map( A => n12, Y => n121);
   U192 : INVX4 port map( A => n10, Y => n112);
   U193 : INVX2 port map( A => n103, Y => n104);
   U194 : INVX1 port map( A => n794, Y => n103);
   U195 : INVX2 port map( A => n106, Y => n107);
   U196 : INVX2 port map( A => n109, Y => n110);
   U197 : INVX1 port map( A => n812, Y => n109);
   U198 : INVX4 port map( A => n18, Y => n111);
   U199 : INVX4 port map( A => n129, Y => n130);
   U200 : AND2X2 port map( A => n264, B => n591, Y => n83);
   U201 : AND2X2 port map( A => n73, B => n591, Y => n84);
   U202 : INVX2 port map( A => n85, Y => n113);
   U203 : INVX2 port map( A => n85, Y => n114);
   U204 : INVX2 port map( A => n145, Y => n144);
   U205 : INVX2 port map( A => n147, Y => n146);
   U206 : INVX2 port map( A => n149, Y => n148);
   U207 : INVX2 port map( A => n151, Y => n150);
   U208 : INVX2 port map( A => n153, Y => n152);
   U209 : INVX2 port map( A => n157, Y => n156);
   U210 : INVX2 port map( A => RCV_DATA(7), Y => n158);
   U211 : INVX2 port map( A => RCV_DATA(7), Y => n159);
   U212 : INVX2 port map( A => n155, Y => n154);
   U213 : OR2X2 port map( A => n614, B => n168, Y => n85);
   U214 : XOR2X1 port map( A => n130, B => n49, Y => n88);
   U215 : INVX2 port map( A => readptr_3_port, Y => n135);
   U216 : INVX2 port map( A => n538, Y => n151);
   U217 : INVX2 port map( A => n540, Y => n155);
   U218 : INVX2 port map( A => n535, Y => n145);
   U219 : INVX2 port map( A => n536, Y => n147);
   U220 : INVX2 port map( A => n537, Y => n149);
   U221 : INVX2 port map( A => n539, Y => n153);
   U222 : INVX2 port map( A => n541, Y => n157);
   U223 : INVX2 port map( A => writeptr_3_port, Y => n99);
   U224 : INVX2 port map( A => n99, Y => n100);
   U225 : INVX2 port map( A => n99, Y => n101);
   U226 : INVX1 port map( A => n100, Y => n587);
   U227 : INVX2 port map( A => writeptr_2_port, Y => n128);
   U228 : AND2X2 port map( A => n1238, B => n1239, Y => n796);
   U229 : AND2X2 port map( A => n1236, B => n1239, Y => n795);
   U230 : AND2X2 port map( A => n1239, B => n1248, Y => n804);
   U231 : AND2X2 port map( A => n1239, B => n1247, Y => n803);
   U232 : AND2X2 port map( A => n1259, B => n1239, Y => n814);
   U233 : AND2X2 port map( A => n1258, B => n1239, Y => n813);
   U234 : AND2X2 port map( A => n1268, B => n1239, Y => n821);
   U235 : AND2X2 port map( A => n1267, B => n1239, Y => n820);
   U236 : INVX2 port map( A => memory_16_7_port, Y => n735);
   U237 : INVX2 port map( A => memory_17_7_port, Y => n743);
   U238 : INVX2 port map( A => memory_18_7_port, Y => n751);
   U239 : INVX2 port map( A => readptr_2_port, Y => n618);
   U240 : INVX2 port map( A => memory_19_7_port, Y => n759);
   U241 : NAND2X1 port map( A => n1236, B => n86, Y => n794);
   U242 : INVX2 port map( A => memory_24_7_port, Y => n661);
   U243 : INVX2 port map( A => memory_25_7_port, Y => n653);
   U244 : INVX2 port map( A => memory_26_7_port, Y => n645);
   U245 : INVX2 port map( A => memory_27_7_port, Y => n637);
   U246 : NAND2X1 port map( A => n1247, B => n86, Y => n802);
   U247 : INVX2 port map( A => memory_3_7_port, Y => n700);
   U248 : INVX2 port map( A => memory_2_7_port, Y => n692);
   U249 : NAND2X1 port map( A => n1258, B => n86, Y => n812);
   U250 : INVX2 port map( A => memory_1_7_port, Y => n684);
   U251 : INVX2 port map( A => memory_0_7_port, Y => n676);
   U252 : INVX2 port map( A => memory_8_7_port, Y => n703);
   U253 : INVX2 port map( A => memory_9_7_port, Y => n711);
   U254 : INVX2 port map( A => memory_10_7_port, Y => n719);
   U255 : INVX2 port map( A => memory_11_7_port, Y => n727);
   U256 : INVX2 port map( A => memory_16_6_port, Y => n736);
   U257 : INVX2 port map( A => memory_17_6_port, Y => n744);
   U258 : INVX2 port map( A => memory_18_6_port, Y => n752);
   U259 : INVX2 port map( A => memory_19_6_port, Y => n760);
   U260 : INVX2 port map( A => memory_24_6_port, Y => n662);
   U261 : INVX2 port map( A => memory_25_6_port, Y => n654);
   U262 : INVX2 port map( A => memory_26_6_port, Y => n646);
   U263 : INVX2 port map( A => memory_27_6_port, Y => n638);
   U264 : INVX2 port map( A => memory_3_6_port, Y => n699);
   U265 : INVX2 port map( A => memory_2_6_port, Y => n691);
   U266 : INVX2 port map( A => memory_1_6_port, Y => n683);
   U267 : INVX2 port map( A => memory_0_6_port, Y => n675);
   U268 : INVX2 port map( A => memory_8_6_port, Y => n704);
   U269 : INVX2 port map( A => memory_9_6_port, Y => n712);
   U270 : INVX2 port map( A => memory_10_6_port, Y => n720);
   U271 : INVX2 port map( A => memory_11_6_port, Y => n728);
   U272 : INVX2 port map( A => memory_16_5_port, Y => n737);
   U273 : INVX2 port map( A => memory_17_5_port, Y => n745);
   U274 : INVX2 port map( A => memory_18_5_port, Y => n753);
   U275 : INVX2 port map( A => memory_19_5_port, Y => n761);
   U276 : INVX2 port map( A => memory_24_5_port, Y => n663);
   U277 : INVX2 port map( A => memory_25_5_port, Y => n655);
   U278 : INVX2 port map( A => memory_26_5_port, Y => n647);
   U279 : INVX2 port map( A => memory_27_5_port, Y => n639);
   U280 : INVX2 port map( A => memory_3_5_port, Y => n698);
   U281 : INVX2 port map( A => memory_2_5_port, Y => n690);
   U282 : INVX2 port map( A => memory_1_5_port, Y => n682);
   U283 : INVX2 port map( A => memory_0_5_port, Y => n674);
   U284 : INVX2 port map( A => memory_8_5_port, Y => n705);
   U285 : INVX2 port map( A => memory_9_5_port, Y => n713);
   U286 : INVX2 port map( A => memory_10_5_port, Y => n721);
   U287 : INVX2 port map( A => memory_11_5_port, Y => n729);
   U288 : INVX2 port map( A => memory_16_4_port, Y => n738);
   U289 : INVX2 port map( A => memory_17_4_port, Y => n746);
   U290 : INVX2 port map( A => memory_18_4_port, Y => n754);
   U291 : INVX2 port map( A => memory_19_4_port, Y => n762);
   U292 : INVX2 port map( A => memory_24_4_port, Y => n664);
   U293 : INVX2 port map( A => memory_25_4_port, Y => n656);
   U294 : INVX2 port map( A => memory_26_4_port, Y => n648);
   U295 : INVX2 port map( A => memory_27_4_port, Y => n640);
   U296 : INVX2 port map( A => memory_3_4_port, Y => n697);
   U297 : INVX2 port map( A => memory_2_4_port, Y => n689);
   U298 : INVX2 port map( A => memory_1_4_port, Y => n681);
   U299 : INVX2 port map( A => memory_0_4_port, Y => n673);
   U300 : INVX2 port map( A => memory_8_4_port, Y => n706);
   U301 : INVX2 port map( A => memory_9_4_port, Y => n714);
   U302 : INVX2 port map( A => memory_10_4_port, Y => n722);
   U303 : INVX2 port map( A => memory_11_4_port, Y => n730);
   U304 : INVX2 port map( A => memory_16_3_port, Y => n739);
   U305 : INVX2 port map( A => memory_17_3_port, Y => n747);
   U306 : INVX2 port map( A => memory_18_3_port, Y => n755);
   U307 : INVX2 port map( A => memory_19_3_port, Y => n763);
   U308 : INVX2 port map( A => memory_24_3_port, Y => n665);
   U309 : INVX2 port map( A => memory_25_3_port, Y => n657);
   U310 : INVX2 port map( A => memory_26_3_port, Y => n649);
   U311 : INVX2 port map( A => memory_27_3_port, Y => n641);
   U312 : INVX2 port map( A => memory_3_3_port, Y => n696);
   U313 : INVX2 port map( A => memory_2_3_port, Y => n688);
   U314 : INVX2 port map( A => memory_1_3_port, Y => n680);
   U315 : INVX2 port map( A => memory_0_3_port, Y => n672);
   U316 : INVX2 port map( A => memory_8_3_port, Y => n707);
   U317 : INVX2 port map( A => memory_9_3_port, Y => n715);
   U318 : INVX2 port map( A => memory_10_3_port, Y => n723);
   U319 : INVX2 port map( A => memory_11_3_port, Y => n731);
   U320 : INVX2 port map( A => memory_16_2_port, Y => n740);
   U321 : INVX2 port map( A => memory_17_2_port, Y => n748);
   U322 : INVX2 port map( A => memory_18_2_port, Y => n756);
   U323 : INVX2 port map( A => memory_19_2_port, Y => n764);
   U324 : INVX2 port map( A => memory_24_2_port, Y => n666);
   U325 : INVX2 port map( A => memory_25_2_port, Y => n658);
   U326 : INVX2 port map( A => memory_26_2_port, Y => n650);
   U327 : INVX2 port map( A => memory_27_2_port, Y => n642);
   U328 : INVX2 port map( A => memory_3_2_port, Y => n695);
   U329 : INVX2 port map( A => memory_2_2_port, Y => n687);
   U330 : INVX2 port map( A => memory_1_2_port, Y => n679);
   U331 : INVX2 port map( A => memory_0_2_port, Y => n671);
   U332 : INVX2 port map( A => memory_8_2_port, Y => n708);
   U333 : INVX2 port map( A => memory_9_2_port, Y => n716);
   U334 : INVX2 port map( A => memory_10_2_port, Y => n724);
   U335 : INVX2 port map( A => memory_11_2_port, Y => n732);
   U336 : INVX2 port map( A => memory_16_1_port, Y => n741);
   U337 : INVX2 port map( A => memory_17_1_port, Y => n749);
   U338 : INVX2 port map( A => memory_18_1_port, Y => n757);
   U339 : INVX2 port map( A => memory_19_1_port, Y => n765);
   U340 : INVX2 port map( A => memory_24_1_port, Y => n667);
   U341 : INVX2 port map( A => memory_25_1_port, Y => n659);
   U342 : INVX2 port map( A => memory_26_1_port, Y => n651);
   U343 : INVX2 port map( A => memory_27_1_port, Y => n643);
   U344 : INVX2 port map( A => memory_3_1_port, Y => n694);
   U345 : INVX2 port map( A => memory_2_1_port, Y => n686);
   U346 : INVX2 port map( A => memory_1_1_port, Y => n678);
   U347 : INVX2 port map( A => memory_0_1_port, Y => n670);
   U348 : INVX2 port map( A => memory_8_1_port, Y => n709);
   U349 : INVX2 port map( A => memory_9_1_port, Y => n717);
   U350 : INVX2 port map( A => memory_10_1_port, Y => n725);
   U351 : INVX2 port map( A => memory_11_1_port, Y => n733);
   U352 : INVX2 port map( A => memory_16_0_port, Y => n742);
   U353 : INVX2 port map( A => memory_17_0_port, Y => n750);
   U354 : INVX2 port map( A => memory_18_0_port, Y => n758);
   U355 : INVX2 port map( A => memory_19_0_port, Y => n766);
   U356 : INVX2 port map( A => memory_24_0_port, Y => n668);
   U357 : INVX2 port map( A => memory_25_0_port, Y => n660);
   U358 : INVX2 port map( A => memory_26_0_port, Y => n652);
   U359 : INVX2 port map( A => memory_27_0_port, Y => n644);
   U360 : INVX2 port map( A => memory_3_0_port, Y => n693);
   U361 : INVX2 port map( A => memory_2_0_port, Y => n685);
   U362 : INVX2 port map( A => memory_1_0_port, Y => n677);
   U363 : INVX2 port map( A => memory_0_0_port, Y => n669);
   U364 : INVX2 port map( A => memory_8_0_port, Y => n710);
   U365 : INVX2 port map( A => memory_9_0_port, Y => n718);
   U366 : INVX2 port map( A => memory_10_0_port, Y => n726);
   U367 : INVX2 port map( A => memory_11_0_port, Y => n734);
   U368 : INVX2 port map( A => opcode_16_1_port, Y => n775);
   U369 : INVX2 port map( A => opcode_17_1_port, Y => n777);
   U370 : INVX2 port map( A => opcode_18_1_port, Y => n779);
   U371 : INVX2 port map( A => opcode_19_1_port, Y => n781);
   U372 : INVX2 port map( A => opcode_24_1_port, Y => n627);
   U373 : INVX2 port map( A => opcode_25_1_port, Y => n625);
   U374 : INVX2 port map( A => opcode_26_1_port, Y => n623);
   U375 : INVX2 port map( A => opcode_27_1_port, Y => n621);
   U376 : INVX2 port map( A => opcode_3_1_port, Y => n636);
   U377 : INVX2 port map( A => opcode_2_1_port, Y => n634);
   U378 : INVX2 port map( A => opcode_1_1_port, Y => n632);
   U379 : INVX2 port map( A => opcode_0_1_port, Y => n630);
   U380 : INVX2 port map( A => opcode_8_1_port, Y => n767);
   U381 : INVX2 port map( A => opcode_9_1_port, Y => n769);
   U382 : INVX2 port map( A => opcode_10_1_port, Y => n771);
   U383 : INVX2 port map( A => opcode_11_1_port, Y => n773);
   U384 : INVX2 port map( A => opcode_16_0_port, Y => n776);
   U385 : INVX2 port map( A => opcode_17_0_port, Y => n778);
   U386 : INVX2 port map( A => opcode_18_0_port, Y => n780);
   U387 : INVX2 port map( A => opcode_19_0_port, Y => n782);
   U388 : INVX2 port map( A => n136, Y => n619);
   U389 : INVX2 port map( A => opcode_24_0_port, Y => n628);
   U390 : INVX2 port map( A => opcode_25_0_port, Y => n626);
   U391 : INVX2 port map( A => opcode_26_0_port, Y => n624);
   U392 : INVX2 port map( A => opcode_27_0_port, Y => n622);
   U393 : INVX2 port map( A => opcode_3_0_port, Y => n635);
   U394 : INVX2 port map( A => opcode_2_0_port, Y => n633);
   U395 : INVX2 port map( A => opcode_1_0_port, Y => n631);
   U396 : INVX2 port map( A => opcode_0_0_port, Y => n629);
   U397 : INVX2 port map( A => opcode_8_0_port, Y => n768);
   U398 : INVX2 port map( A => opcode_9_0_port, Y => n770);
   U399 : INVX2 port map( A => opcode_10_0_port, Y => n772);
   U400 : INVX2 port map( A => opcode_11_0_port, Y => n774);
   U401 : NAND2X1 port map( A => readptr_0_port, B => n219, Y => n545);
   U402 : NAND2X1 port map( A => n134, B => n617, Y => n164);
   U403 : XNOR2X1 port map( A => n70, B => n43, Y => n548);
   U404 : XNOR2X1 port map( A => n101, B => n136, Y => n553);
   U405 : XNOR2X1 port map( A => writeptr_4_port, B => readptr_4_port, Y => 
                           n558);
   U406 : AND2X2 port map( A => n553, B => n558, Y => n165);
   U407 : NAND3X1 port map( A => n166, B => n548, C => n165, Y => n167);
   U408 : MUX2X1 port map( B => n167, A => n702, S => RST, Y => n1432);
   U409 : INVX2 port map( A => OUT_OPCODE_0_port, Y => n170);
   U410 : INVX2 port map( A => n1226, Y => n169);
   U411 : NAND2X1 port map( A => R_ENABLE, B => n167, Y => n614);
   U412 : NAND2X1 port map( A => n163, B => state, Y => n168);
   U413 : MUX2X1 port map( B => n170, A => n169, S => n113, Y => n1562);
   U414 : INVX2 port map( A => OUT_OPCODE_1_port, Y => n172);
   U415 : INVX2 port map( A => n1199, Y => n171);
   U416 : MUX2X1 port map( B => n172, A => n171, S => n114, Y => n1561);
   U417 : INVX2 port map( A => DATA_0_port, Y => n174);
   U418 : INVX2 port map( A => n1172, Y => n173);
   U419 : MUX2X1 port map( B => n174, A => n173, S => n113, Y => n1560);
   U420 : INVX2 port map( A => DATA_1_port, Y => n176);
   U421 : INVX2 port map( A => n1015, Y => n175);
   U422 : MUX2X1 port map( B => n176, A => n175, S => n114, Y => n1559);
   U423 : INVX2 port map( A => DATA_2_port, Y => n178);
   U424 : INVX2 port map( A => n988, Y => n177);
   U425 : MUX2X1 port map( B => n178, A => n177, S => n113, Y => n1558);
   U426 : INVX2 port map( A => DATA_3_port, Y => n180);
   U427 : INVX2 port map( A => n961, Y => n179);
   U428 : MUX2X1 port map( B => n180, A => n179, S => n114, Y => n1557);
   U429 : INVX2 port map( A => DATA_4_port, Y => n182);
   U430 : INVX2 port map( A => n934, Y => n181);
   U431 : MUX2X1 port map( B => n182, A => n181, S => n113, Y => n1556);
   U432 : INVX2 port map( A => DATA_5_port, Y => n184);
   U433 : INVX2 port map( A => n863, Y => n183);
   U434 : MUX2X1 port map( B => n184, A => n183, S => n114, Y => n1555);
   U435 : INVX2 port map( A => DATA_6_port, Y => n186);
   U436 : INVX2 port map( A => n822, Y => n185);
   U437 : MUX2X1 port map( B => n186, A => n185, S => n113, Y => n1554);
   U438 : INVX2 port map( A => DATA_7_port, Y => n188);
   U439 : INVX2 port map( A => n783, Y => n187);
   U440 : MUX2X1 port map( B => n188, A => n187, S => n114, Y => n1553);
   U441 : INVX2 port map( A => RCV_OPCODE(0), Y => n339_port);
   U442 : INVX2 port map( A => opcode_31_0_port, Y => n195);
   U443 : INVX2 port map( A => n130, Y => n203);
   U444 : NAND3X1 port map( A => n134, B => n218, C => n203, Y => n328);
   U445 : NAND3X1 port map( A => n134, B => n218, C => n131, Y => n331);
   U446 : NAND2X1 port map( A => n70, B => n28, Y => n189);
   U447 : NAND2X1 port map( A => n331, B => n189, Y => n569);
   U448 : NAND3X1 port map( A => n70, B => n134, C => n130, Y => n586);
   U449 : INVX2 port map( A => n562, Y => n190);
   U450 : NOR2X1 port map( A => n41, B => n190, Y => n192);
   U451 : INVX2 port map( A => n49, Y => n611);
   U452 : XNOR2X1 port map( A => n575, B => n611, Y => n565);
   U453 : NAND3X1 port map( A => n100, B => n63, C => n70, Y => n592);
   U454 : AND2X2 port map( A => n565, B => n563, Y => n191);
   U455 : NAND3X1 port map( A => n192, B => n64, C => n191, Y => n299);
   U456 : NAND3X1 port map( A => n72, B => n67, C => n84, Y => n336);
   U457 : NAND2X1 port map( A => n100, B => n163, Y => n286);
   U458 : INVX2 port map( A => n286, Y => n264);
   U459 : NAND3X1 port map( A => n89, B => W_ENABLE, C => n299, Y => n226);
   U460 : NOR2X1 port map( A => n31, B => n59, Y => n193);
   U461 : NAND2X1 port map( A => RCV_OPCODE(1), B => RCV_OPCODE(0), Y => n568);
   U462 : NAND2X1 port map( A => n193, B => n160, Y => n342_port);
   U463 : OAI21X1 port map( A => n328, B => n95, C => n342_port, Y => n194);
   U464 : INVX2 port map( A => n194, Y => n196);
   U465 : MUX2X1 port map( B => n137, A => n195, S => n196, Y => n1552);
   U466 : INVX2 port map( A => opcode_31_1_port, Y => n197);
   U467 : MUX2X1 port map( B => n140, A => n197, S => n196, Y => n1551);
   U468 : INVX2 port map( A => opcode_30_0_port, Y => n200);
   U469 : OR2X2 port map( A => n130, B => n134, Y => n577);
   U470 : INVX2 port map( A => n577, Y => n209);
   U471 : NAND3X1 port map( A => n70, B => n130, C => n219, Y => n316);
   U472 : NOR2X1 port map( A => n316, B => n59, Y => n198);
   U473 : NAND2X1 port map( A => n161, B => n198, Y => n352);
   U474 : OAI21X1 port map( A => n118, B => n96, C => n352, Y => n199);
   U475 : INVX2 port map( A => n199, Y => n201);
   U476 : MUX2X1 port map( B => n138, A => n200, S => n201, Y => n1550);
   U477 : INVX2 port map( A => opcode_30_1_port, Y => n202);
   U478 : MUX2X1 port map( B => n142, A => n202, S => n201, Y => n1549);
   U479 : INVX2 port map( A => opcode_29_0_port, Y => n206);
   U480 : NAND3X1 port map( A => n72, B => n67, C => n89, Y => n236);
   U481 : NAND3X1 port map( A => n70, B => n134, C => n203, Y => n321);
   U482 : NOR2X1 port map( A => n321, B => n59, Y => n204);
   U483 : NAND2X1 port map( A => n1, B => n204, Y => n362);
   U484 : OAI21X1 port map( A => n31, B => n94, C => n362, Y => n205);
   U485 : INVX2 port map( A => n205, Y => n207);
   U486 : MUX2X1 port map( B => n339_port, A => n206, S => n207, Y => n1548);
   U487 : INVX2 port map( A => opcode_29_1_port, Y => n208);
   U488 : MUX2X1 port map( B => n142, A => n208, S => n207, Y => n1547);
   U489 : INVX2 port map( A => opcode_28_0_port, Y => n212);
   U490 : NAND2X1 port map( A => n209, B => n70, Y => n325);
   U491 : NOR2X1 port map( A => n325, B => n59, Y => n210);
   U492 : NAND2X1 port map( A => n161, B => n210, Y => n372);
   U493 : OAI21X1 port map( A => n316, B => n94, C => n372, Y => n211);
   U494 : INVX2 port map( A => n211, Y => n213);
   U495 : MUX2X1 port map( B => n339_port, A => n212, S => n213, Y => n1546);
   U496 : INVX2 port map( A => opcode_28_1_port, Y => n214);
   U497 : MUX2X1 port map( B => n142, A => n214, S => n213, Y => n1545);
   U498 : NOR2X1 port map( A => n116, B => n59, Y => n215);
   U499 : NAND2X1 port map( A => n215, B => n2, Y => n382);
   U500 : OAI21X1 port map( A => n321, B => n93, C => n382, Y => n216);
   U501 : INVX2 port map( A => n216, Y => n217);
   U502 : MUX2X1 port map( B => n339_port, A => n622, S => n217, Y => n1272);
   U503 : MUX2X1 port map( B => n142, A => n621, S => n217, Y => n1271);
   U504 : NAND3X1 port map( A => n131, B => n219, C => n218, Y => n337);
   U505 : NOR2X1 port map( A => n337, B => n59, Y => n220);
   U506 : NAND2X1 port map( A => n160, B => n220, Y => n384);
   U507 : OAI21X1 port map( A => n325, B => n93, C => n384, Y => n221);
   U508 : INVX2 port map( A => n221, Y => n222);
   U509 : MUX2X1 port map( B => n339_port, A => n624, S => n222, Y => n1274);
   U510 : MUX2X1 port map( B => n142, A => n623, S => n222, Y => n1273);
   U511 : NOR2X1 port map( A => n328, B => n59, Y => n223);
   U512 : NAND2X1 port map( A => n223, B => n160, Y => n386);
   U513 : OAI21X1 port map( A => n116, B => n94, C => n386, Y => n224);
   U514 : INVX2 port map( A => n224, Y => n225);
   U515 : MUX2X1 port map( B => n339_port, A => n626, S => n225, Y => n1276);
   U516 : MUX2X1 port map( B => n142, A => n625, S => n225, Y => n1275);
   U517 : NOR2X1 port map( A => n118, B => n59, Y => n227);
   U518 : NAND2X1 port map( A => n227, B => n160, Y => n388);
   U519 : OAI21X1 port map( A => n337, B => n94, C => n388, Y => n228);
   U520 : INVX2 port map( A => n228, Y => n229);
   U521 : MUX2X1 port map( B => n339_port, A => n628, S => n229, Y => n1278);
   U522 : MUX2X1 port map( B => n142, A => n627, S => n229, Y => n1277);
   U523 : INVX2 port map( A => opcode_23_0_port, Y => n232);
   U524 : NAND3X1 port map( A => n90, B => W_ENABLE, C => n299, Y => n260);
   U525 : NOR2X1 port map( A => n31, B => n61, Y => n230);
   U526 : NAND2X1 port map( A => n2, B => n230, Y => n390);
   U527 : OAI21X1 port map( A => n328, B => n93, C => n4, Y => n231);
   U528 : INVX2 port map( A => n231, Y => n233);
   U529 : MUX2X1 port map( B => n138, A => n232, S => n233, Y => n1280);
   U530 : INVX2 port map( A => opcode_23_1_port, Y => n234);
   U531 : MUX2X1 port map( B => n141, A => n234, S => n233, Y => n1279);
   U532 : INVX2 port map( A => opcode_22_0_port, Y => n238);
   U533 : NOR2X1 port map( A => n316, B => n61, Y => n235);
   U534 : NAND2X1 port map( A => n160, B => n235, Y => n400);
   U535 : OAI21X1 port map( A => n118, B => n94, C => n400, Y => n237);
   U536 : INVX2 port map( A => n237, Y => n239);
   U537 : MUX2X1 port map( B => n138, A => n238, S => n239, Y => n1282);
   U538 : INVX2 port map( A => opcode_22_1_port, Y => n240);
   U539 : MUX2X1 port map( B => n141, A => n240, S => n239, Y => n1281);
   U540 : INVX2 port map( A => opcode_21_0_port, Y => n243);
   U541 : NAND3X1 port map( A => n72, B => n67, C => n90, Y => n271);
   U542 : NOR2X1 port map( A => n321, B => n61, Y => n241);
   U543 : NAND2X1 port map( A => n161, B => n241, Y => n410);
   U544 : OAI21X1 port map( A => n31, B => n97, C => n5, Y => n242);
   U545 : INVX2 port map( A => n242, Y => n244);
   U546 : MUX2X1 port map( B => n138, A => n243, S => n244, Y => n1284);
   U547 : INVX2 port map( A => opcode_21_1_port, Y => n245);
   U548 : MUX2X1 port map( B => n141, A => n245, S => n244, Y => n1283);
   U549 : INVX2 port map( A => opcode_20_0_port, Y => n248);
   U550 : NOR2X1 port map( A => n325, B => n61, Y => n246);
   U551 : NAND2X1 port map( A => n160, B => n246, Y => n420);
   U552 : OAI21X1 port map( A => n316, B => n97, C => n420, Y => n247);
   U553 : MUX2X1 port map( B => n138, A => n248, S => n249, Y => n1286);
   U554 : INVX2 port map( A => opcode_20_1_port, Y => n250);
   U555 : MUX2X1 port map( B => n141, A => n250, S => n249, Y => n1285);
   U556 : NOR2X1 port map( A => n116, B => n61, Y => n251);
   U557 : NAND2X1 port map( A => n251, B => n161, Y => n430);
   U558 : OAI21X1 port map( A => n321, B => n97, C => n430, Y => n252);
   U559 : INVX2 port map( A => n252, Y => n253);
   U560 : MUX2X1 port map( B => n138, A => n782, S => n253, Y => n1544);
   U561 : MUX2X1 port map( B => n141, A => n781, S => n253, Y => n1543);
   U562 : NOR2X1 port map( A => n337, B => n61, Y => n254);
   U563 : NAND2X1 port map( A => n160, B => n254, Y => n432);
   U564 : OAI21X1 port map( A => n325, B => n98, C => n432, Y => n255);
   U565 : INVX2 port map( A => n255, Y => n256);
   U566 : MUX2X1 port map( B => n138, A => n780, S => n256, Y => n1542);
   U567 : MUX2X1 port map( B => n141, A => n779, S => n256, Y => n1541);
   U568 : NOR2X1 port map( A => n328, B => n61, Y => n257);
   U569 : NAND2X1 port map( A => n161, B => n257, Y => n434);
   U570 : OAI21X1 port map( A => n116, B => n98, C => n434, Y => n258);
   U571 : INVX2 port map( A => n258, Y => n259);
   U572 : MUX2X1 port map( B => n138, A => n778, S => n259, Y => n1540);
   U573 : MUX2X1 port map( B => n141, A => n777, S => n259, Y => n1539);
   U574 : NOR2X1 port map( A => n118, B => n61, Y => n261);
   U575 : NAND2X1 port map( A => n261, B => n160, Y => n436);
   U576 : OAI21X1 port map( A => n337, B => n98, C => n436, Y => n262);
   U577 : INVX2 port map( A => n262, Y => n263);
   U578 : MUX2X1 port map( B => n138, A => n776, S => n263, Y => n1538);
   U579 : MUX2X1 port map( B => n141, A => n775, S => n263, Y => n1537);
   U580 : INVX2 port map( A => opcode_15_0_port, Y => n267);
   U581 : NOR2X1 port map( A => n31, B => n478, Y => n265);
   U582 : NAND2X1 port map( A => n161, B => n265, Y => n438);
   U583 : OAI21X1 port map( A => n328, B => n98, C => n438, Y => n266);
   U584 : MUX2X1 port map( B => n138, A => n267, S => n268, Y => n1288);
   U585 : INVX2 port map( A => opcode_15_1_port, Y => n269);
   U586 : MUX2X1 port map( B => n141, A => n269, S => n268, Y => n1287);
   U587 : INVX2 port map( A => opcode_14_0_port, Y => n273);
   U588 : NOR2X1 port map( A => n68, B => n69, Y => n270);
   U589 : NAND2X1 port map( A => n270, B => n161, Y => n448);
   U590 : OAI21X1 port map( A => n118, B => n98, C => n448, Y => n272);
   U591 : INVX2 port map( A => n272, Y => n274);
   U592 : MUX2X1 port map( B => n138, A => n273, S => n274, Y => n1290);
   U593 : INVX2 port map( A => opcode_14_1_port, Y => n275);
   U594 : MUX2X1 port map( B => n141, A => n275, S => n274, Y => n1289);
   U595 : INVX2 port map( A => opcode_13_0_port, Y => n278);
   U596 : NAND3X1 port map( A => n72, B => n67, C => n83, Y => n305);
   U597 : NOR2X1 port map( A => n321, B => n47, Y => n276);
   U598 : NAND2X1 port map( A => n276, B => n161, Y => n458);
   U599 : OAI21X1 port map( A => n31, B => n92, C => n458, Y => n277);
   U600 : INVX2 port map( A => n277, Y => n279);
   U601 : MUX2X1 port map( B => n138, A => n278, S => n279, Y => n1292);
   U602 : INVX2 port map( A => opcode_13_1_port, Y => n280);
   U603 : MUX2X1 port map( B => n141, A => n280, S => n279, Y => n1291);
   U604 : INVX2 port map( A => opcode_12_0_port, Y => n283);
   U605 : NOR2X1 port map( A => n325, B => n47, Y => n281);
   U606 : NAND2X1 port map( A => n281, B => n161, Y => n468);
   U607 : OAI21X1 port map( A => n316, B => n91, C => n468, Y => n282);
   U608 : INVX2 port map( A => n282, Y => n284);
   U609 : MUX2X1 port map( B => n137, A => n283, S => n284, Y => n1294);
   U610 : INVX2 port map( A => opcode_12_1_port, Y => n285);
   U611 : MUX2X1 port map( B => n140, A => n285, S => n284, Y => n1293);
   U612 : NOR3X1 port map( A => n52, B => n579, C => n286, Y => n288);
   U613 : AND2X2 port map( A => n288, B => n287, Y => n289);
   U614 : MUX2X1 port map( B => n774, A => n137, S => n289, Y => n1536);
   U615 : MUX2X1 port map( B => n773, A => n142, S => n289, Y => n1535);
   U616 : NOR2X1 port map( A => n337, B => n478, Y => n290);
   U617 : NAND2X1 port map( A => n290, B => n161, Y => n482);
   U618 : OAI21X1 port map( A => n325, B => n92, C => n482, Y => n291);
   U619 : INVX2 port map( A => n291, Y => n292);
   U620 : MUX2X1 port map( B => n137, A => n772, S => n292, Y => n1534);
   U621 : MUX2X1 port map( B => n140, A => n771, S => n292, Y => n1533);
   U622 : NOR2X1 port map( A => n328, B => n47, Y => n293);
   U623 : NAND2X1 port map( A => n293, B => n160, Y => n484);
   U624 : OAI21X1 port map( A => n116, B => n92, C => n484, Y => n294);
   U625 : INVX2 port map( A => n294, Y => n295);
   U626 : MUX2X1 port map( B => n137, A => n770, S => n295, Y => n1532);
   U627 : MUX2X1 port map( B => n140, A => n769, S => n295, Y => n1531);
   U628 : NOR2X1 port map( A => n478, B => n118, Y => n296);
   U629 : NAND2X1 port map( A => n161, B => n296, Y => n486);
   U630 : OAI21X1 port map( A => n337, B => n91, C => n486, Y => n297);
   U631 : MUX2X1 port map( B => n137, A => n768, S => n298, Y => n1530);
   U632 : MUX2X1 port map( B => n140, A => n767, S => n298, Y => n1529);
   U633 : INVX2 port map( A => opcode_7_0_port, Y => n301);
   U634 : NAND3X1 port map( A => n84, B => n24, C => W_ENABLE, Y => n334);
   U635 : INVX2 port map( A => n334, Y => n329);
   U636 : NAND3X1 port map( A => n117, B => n329, C => n2, Y => n488);
   U637 : OAI21X1 port map( A => n328, B => n91, C => n488, Y => n300);
   U638 : INVX2 port map( A => n300, Y => n302);
   U639 : MUX2X1 port map( B => n137, A => n301, S => n302, Y => n1563);
   U640 : INVX2 port map( A => opcode_7_1_port, Y => n303);
   U641 : MUX2X1 port map( B => n140, A => n303, S => n302, Y => n1564);
   U642 : INVX2 port map( A => opcode_6_0_port, Y => n307);
   U643 : INVX2 port map( A => n316, Y => n304);
   U644 : NAND3X1 port map( A => n304, B => n329, C => n2, Y => n498);
   U645 : OAI21X1 port map( A => n118, B => n92, C => n498, Y => n306);
   U646 : INVX2 port map( A => n306, Y => n308);
   U647 : MUX2X1 port map( B => n137, A => n307, S => n308, Y => n1573);
   U648 : INVX2 port map( A => opcode_6_1_port, Y => n309);
   U649 : MUX2X1 port map( B => n140, A => n309, S => n308, Y => n1574);
   U650 : INVX2 port map( A => opcode_5_0_port, Y => n312);
   U651 : INVX2 port map( A => n321, Y => n310);
   U652 : NAND3X1 port map( A => n310, B => n329, C => n2, Y => n508);
   U653 : OAI21X1 port map( A => n31, B => n95, C => n508, Y => n311);
   U654 : INVX2 port map( A => n311, Y => n313);
   U655 : MUX2X1 port map( B => n137, A => n312, S => n313, Y => n1583);
   U656 : INVX2 port map( A => opcode_5_1_port, Y => n314);
   U657 : MUX2X1 port map( B => n140, A => n314, S => n313, Y => n1584);
   U658 : INVX2 port map( A => opcode_4_0_port, Y => n318);
   U659 : INVX2 port map( A => n325, Y => n315);
   U660 : NAND3X1 port map( A => n315, B => n329, C => n2, Y => n518);
   U661 : OAI21X1 port map( A => n316, B => n95, C => n518, Y => n317);
   U662 : INVX2 port map( A => n317, Y => n319);
   U663 : MUX2X1 port map( B => n137, A => n318, S => n319, Y => n1593);
   U664 : INVX2 port map( A => opcode_4_1_port, Y => n320);
   U665 : MUX2X1 port map( B => n140, A => n320, S => n319, Y => n1594);
   U666 : NAND3X1 port map( A => n115, B => n329, C => n2, Y => n528);
   U667 : OAI21X1 port map( A => n321, B => n96, C => n528, Y => n322);
   U668 : MUX2X1 port map( B => n137, A => n635, S => n323, Y => n1301);
   U669 : MUX2X1 port map( B => n140, A => n636, S => n323, Y => n1302);
   U670 : INVX2 port map( A => n337, Y => n324);
   U671 : NAND3X1 port map( A => n324, B => n329, C => n2, Y => n530);
   U672 : OAI21X1 port map( A => n325, B => n96, C => n530, Y => n326);
   U673 : INVX2 port map( A => n326, Y => n327);
   U674 : MUX2X1 port map( B => n137, A => n633, S => n327, Y => n1299);
   U675 : MUX2X1 port map( B => n140, A => n634, S => n327, Y => n1300);
   U676 : INVX2 port map( A => n328, Y => n330);
   U677 : NAND3X1 port map( A => n330, B => n329, C => n160, Y => n532);
   U678 : OAI21X1 port map( A => n116, B => n96, C => n532, Y => n332);
   U679 : INVX2 port map( A => n332, Y => n333);
   U680 : MUX2X1 port map( B => n137, A => n631, S => n333, Y => n1297);
   U681 : MUX2X1 port map( B => n140, A => n632, S => n333, Y => n1298);
   U682 : NOR2X1 port map( A => n118, B => n334, Y => n335);
   U683 : NAND2X1 port map( A => n335, B => n2, Y => n534);
   U684 : OAI21X1 port map( A => n337, B => n96, C => n534, Y => n338_port);
   U685 : INVX2 port map( A => n338_port, Y => n340_port);
   U686 : MUX2X1 port map( B => n138, A => n629, S => n340_port, Y => n1295);
   U687 : MUX2X1 port map( B => n141, A => n630, S => n340_port, Y => n1296);
   U688 : INVX2 port map( A => memory_31_0_port, Y => n343_port);
   U689 : MUX2X1 port map( B => n343_port, A => n144, S => n350, Y => n1528);
   U690 : INVX2 port map( A => memory_31_1_port, Y => n344_port);
   U691 : MUX2X1 port map( B => n344_port, A => n146, S => n350, Y => n1527);
   U692 : INVX2 port map( A => memory_31_2_port, Y => n345_port);
   U693 : MUX2X1 port map( B => n345_port, A => n148, S => n350, Y => n1526);
   U694 : INVX2 port map( A => memory_31_3_port, Y => n346_port);
   U695 : MUX2X1 port map( B => n346_port, A => n150, S => n350, Y => n1525);
   U696 : INVX2 port map( A => memory_31_4_port, Y => n347_port);
   U697 : MUX2X1 port map( B => n347_port, A => n152, S => n350, Y => n1524);
   U698 : INVX2 port map( A => memory_31_5_port, Y => n348);
   U699 : MUX2X1 port map( B => n348, A => n154, S => n350, Y => n1523);
   U700 : INVX2 port map( A => memory_31_6_port, Y => n349);
   U701 : MUX2X1 port map( B => n349, A => n156, S => n350, Y => n1522);
   U702 : INVX2 port map( A => memory_31_7_port, Y => n351);
   U703 : MUX2X1 port map( B => n351, A => n158, S => n350, Y => n1521);
   U704 : INVX2 port map( A => memory_30_0_port, Y => n353);
   U705 : MUX2X1 port map( B => n353, A => n144, S => n360, Y => n1520);
   U706 : INVX2 port map( A => memory_30_1_port, Y => n354);
   U707 : MUX2X1 port map( B => n354, A => n146, S => n360, Y => n1519);
   U708 : INVX2 port map( A => memory_30_2_port, Y => n355);
   U709 : MUX2X1 port map( B => n355, A => n148, S => n360, Y => n1518);
   U710 : INVX2 port map( A => memory_30_3_port, Y => n356);
   U711 : MUX2X1 port map( B => n356, A => n150, S => n360, Y => n1517);
   U712 : INVX2 port map( A => memory_30_4_port, Y => n357);
   U713 : MUX2X1 port map( B => n357, A => n152, S => n360, Y => n1516);
   U714 : INVX2 port map( A => memory_30_5_port, Y => n358);
   U715 : MUX2X1 port map( B => n358, A => n154, S => n360, Y => n1515);
   U716 : INVX2 port map( A => memory_30_6_port, Y => n359);
   U717 : MUX2X1 port map( B => n359, A => n156, S => n360, Y => n1514);
   U718 : INVX2 port map( A => memory_30_7_port, Y => n361);
   U719 : MUX2X1 port map( B => n361, A => n158, S => n360, Y => n1513);
   U720 : INVX2 port map( A => memory_29_0_port, Y => n363);
   U721 : MUX2X1 port map( B => n363, A => n144, S => n370, Y => n1512);
   U722 : INVX2 port map( A => memory_29_1_port, Y => n364);
   U723 : MUX2X1 port map( B => n364, A => n146, S => n370, Y => n1511);
   U724 : INVX2 port map( A => memory_29_2_port, Y => n365);
   U725 : MUX2X1 port map( B => n365, A => n148, S => n370, Y => n1510);
   U726 : INVX2 port map( A => memory_29_3_port, Y => n366);
   U727 : MUX2X1 port map( B => n366, A => n150, S => n370, Y => n1509);
   U728 : INVX2 port map( A => memory_29_4_port, Y => n367);
   U729 : MUX2X1 port map( B => n367, A => n152, S => n370, Y => n1508);
   U730 : INVX2 port map( A => memory_29_5_port, Y => n368);
   U731 : MUX2X1 port map( B => n368, A => n154, S => n370, Y => n1507);
   U732 : INVX2 port map( A => memory_29_6_port, Y => n369);
   U733 : MUX2X1 port map( B => n369, A => n156, S => n370, Y => n1506);
   U734 : INVX2 port map( A => memory_29_7_port, Y => n371);
   U735 : MUX2X1 port map( B => n371, A => n158, S => n370, Y => n1505);
   U736 : INVX2 port map( A => memory_28_0_port, Y => n373);
   U737 : MUX2X1 port map( B => n373, A => n144, S => n380, Y => n1504);
   U738 : INVX2 port map( A => memory_28_1_port, Y => n374);
   U739 : MUX2X1 port map( B => n374, A => n146, S => n380, Y => n1503);
   U740 : INVX2 port map( A => memory_28_2_port, Y => n375);
   U741 : MUX2X1 port map( B => n375, A => n148, S => n380, Y => n1502);
   U742 : INVX2 port map( A => memory_28_3_port, Y => n376);
   U743 : MUX2X1 port map( B => n376, A => n150, S => n380, Y => n1501);
   U744 : INVX2 port map( A => memory_28_4_port, Y => n377);
   U745 : MUX2X1 port map( B => n377, A => n152, S => n380, Y => n1500);
   U746 : INVX2 port map( A => memory_28_5_port, Y => n378);
   U747 : MUX2X1 port map( B => n378, A => n154, S => n380, Y => n1499);
   U748 : INVX2 port map( A => memory_28_6_port, Y => n379);
   U749 : MUX2X1 port map( B => n379, A => n156, S => n380, Y => n1498);
   U750 : INVX2 port map( A => memory_28_7_port, Y => n381);
   U751 : MUX2X1 port map( B => n381, A => n158, S => n380, Y => n1497);
   U752 : MUX2X1 port map( B => n644, A => n144, S => n383, Y => n1310);
   U753 : MUX2X1 port map( B => n643, A => n146, S => n383, Y => n1309);
   U754 : MUX2X1 port map( B => n642, A => n148, S => n383, Y => n1308);
   U755 : MUX2X1 port map( B => n641, A => n150, S => n383, Y => n1307);
   U756 : MUX2X1 port map( B => n640, A => n152, S => n383, Y => n1306);
   U757 : MUX2X1 port map( B => n639, A => n154, S => n383, Y => n1305);
   U758 : MUX2X1 port map( B => n638, A => n156, S => n383, Y => n1304);
   U759 : MUX2X1 port map( B => n637, A => n158, S => n383, Y => n1303);
   U760 : MUX2X1 port map( B => n652, A => n144, S => n385, Y => n1318);
   U761 : MUX2X1 port map( B => n651, A => n146, S => n385, Y => n1317);
   U762 : MUX2X1 port map( B => n650, A => n148, S => n385, Y => n1316);
   U763 : MUX2X1 port map( B => n649, A => n150, S => n385, Y => n1315);
   U764 : MUX2X1 port map( B => n648, A => n152, S => n385, Y => n1314);
   U765 : MUX2X1 port map( B => n647, A => n154, S => n385, Y => n1313);
   U766 : MUX2X1 port map( B => n646, A => n156, S => n385, Y => n1312);
   U767 : MUX2X1 port map( B => n645, A => n158, S => n385, Y => n1311);
   U768 : MUX2X1 port map( B => n660, A => n144, S => n387, Y => n1326);
   U769 : MUX2X1 port map( B => n659, A => n146, S => n387, Y => n1325);
   U770 : MUX2X1 port map( B => n658, A => n148, S => n387, Y => n1324);
   U771 : MUX2X1 port map( B => n657, A => n150, S => n387, Y => n1323);
   U772 : MUX2X1 port map( B => n656, A => n152, S => n387, Y => n1322);
   U773 : MUX2X1 port map( B => n655, A => n154, S => n387, Y => n1321);
   U774 : MUX2X1 port map( B => n654, A => n156, S => n387, Y => n1320);
   U775 : MUX2X1 port map( B => n653, A => n158, S => n387, Y => n1319);
   U776 : MUX2X1 port map( B => n668, A => n144, S => n389, Y => n1334);
   U777 : MUX2X1 port map( B => n667, A => n146, S => n389, Y => n1333);
   U778 : MUX2X1 port map( B => n666, A => n148, S => n389, Y => n1332);
   U779 : MUX2X1 port map( B => n665, A => n150, S => n389, Y => n1331);
   U780 : MUX2X1 port map( B => n664, A => n152, S => n389, Y => n1330);
   U781 : MUX2X1 port map( B => n663, A => n540, S => n389, Y => n1329);
   U782 : MUX2X1 port map( B => n662, A => n156, S => n389, Y => n1328);
   U783 : MUX2X1 port map( B => n661, A => n158, S => n389, Y => n1327);
   U784 : INVX2 port map( A => memory_23_0_port, Y => n391);
   U785 : MUX2X1 port map( B => n391, A => n144, S => n398, Y => n1342);
   U786 : INVX2 port map( A => memory_23_1_port, Y => n392);
   U787 : MUX2X1 port map( B => n392, A => n146, S => n398, Y => n1341);
   U788 : INVX2 port map( A => memory_23_2_port, Y => n393);
   U789 : MUX2X1 port map( B => n393, A => n148, S => n398, Y => n1340);
   U790 : INVX2 port map( A => memory_23_3_port, Y => n394);
   U791 : MUX2X1 port map( B => n394, A => n150, S => n398, Y => n1339);
   U792 : INVX2 port map( A => memory_23_4_port, Y => n395);
   U793 : MUX2X1 port map( B => n395, A => n152, S => n398, Y => n1338);
   U794 : INVX2 port map( A => memory_23_5_port, Y => n396);
   U795 : MUX2X1 port map( B => n396, A => n540, S => n398, Y => n1337);
   U796 : INVX2 port map( A => memory_23_6_port, Y => n397);
   U797 : MUX2X1 port map( B => n397, A => n156, S => n398, Y => n1336);
   U798 : INVX2 port map( A => memory_23_7_port, Y => n399);
   U799 : MUX2X1 port map( B => n399, A => n158, S => n398, Y => n1335);
   U800 : INVX2 port map( A => memory_22_0_port, Y => n401);
   U801 : MUX2X1 port map( B => n401, A => n144, S => n408, Y => n1350);
   U802 : INVX2 port map( A => memory_22_1_port, Y => n402);
   U803 : MUX2X1 port map( B => n402, A => n146, S => n408, Y => n1349);
   U804 : INVX2 port map( A => memory_22_2_port, Y => n403);
   U805 : MUX2X1 port map( B => n403, A => n148, S => n408, Y => n1348);
   U806 : INVX2 port map( A => memory_22_3_port, Y => n404);
   U807 : MUX2X1 port map( B => n404, A => n150, S => n408, Y => n1347);
   U808 : INVX2 port map( A => memory_22_4_port, Y => n405);
   U809 : MUX2X1 port map( B => n405, A => n152, S => n408, Y => n1346);
   U810 : INVX2 port map( A => memory_22_5_port, Y => n406);
   U811 : MUX2X1 port map( B => n406, A => n540, S => n408, Y => n1345);
   U812 : INVX2 port map( A => memory_22_6_port, Y => n407);
   U813 : MUX2X1 port map( B => n407, A => n156, S => n408, Y => n1344);
   U814 : INVX2 port map( A => memory_22_7_port, Y => n409);
   U815 : MUX2X1 port map( B => n409, A => n158, S => n408, Y => n1343);
   U816 : INVX2 port map( A => memory_21_0_port, Y => n411);
   U817 : MUX2X1 port map( B => n411, A => n144, S => n418, Y => n1358);
   U818 : INVX2 port map( A => memory_21_1_port, Y => n412);
   U819 : MUX2X1 port map( B => n412, A => n146, S => n418, Y => n1357);
   U820 : INVX2 port map( A => memory_21_2_port, Y => n413);
   U821 : MUX2X1 port map( B => n413, A => n148, S => n418, Y => n1356);
   U822 : INVX2 port map( A => memory_21_3_port, Y => n414);
   U823 : MUX2X1 port map( B => n414, A => n150, S => n418, Y => n1355);
   U824 : INVX2 port map( A => memory_21_4_port, Y => n415);
   U825 : MUX2X1 port map( B => n415, A => n152, S => n418, Y => n1354);
   U826 : INVX2 port map( A => memory_21_5_port, Y => n416);
   U827 : MUX2X1 port map( B => n416, A => n540, S => n418, Y => n1353);
   U828 : INVX2 port map( A => memory_21_6_port, Y => n417);
   U829 : MUX2X1 port map( B => n417, A => n156, S => n418, Y => n1352);
   U830 : INVX2 port map( A => memory_21_7_port, Y => n419);
   U831 : MUX2X1 port map( B => n419, A => n158, S => n418, Y => n1351);
   U832 : INVX2 port map( A => memory_20_0_port, Y => n421);
   U833 : MUX2X1 port map( B => n421, A => n144, S => n428, Y => n1366);
   U834 : INVX2 port map( A => memory_20_1_port, Y => n422);
   U835 : MUX2X1 port map( B => n422, A => n146, S => n428, Y => n1365);
   U836 : INVX2 port map( A => memory_20_2_port, Y => n423);
   U837 : MUX2X1 port map( B => n423, A => n148, S => n428, Y => n1364);
   U838 : INVX2 port map( A => memory_20_3_port, Y => n424);
   U839 : MUX2X1 port map( B => n424, A => n150, S => n428, Y => n1363);
   U840 : INVX2 port map( A => memory_20_4_port, Y => n425);
   U841 : MUX2X1 port map( B => n425, A => n152, S => n428, Y => n1362);
   U842 : INVX2 port map( A => memory_20_5_port, Y => n426);
   U843 : MUX2X1 port map( B => n426, A => n154, S => n428, Y => n1361);
   U844 : INVX2 port map( A => memory_20_6_port, Y => n427);
   U845 : MUX2X1 port map( B => n427, A => n156, S => n428, Y => n1360);
   U846 : INVX2 port map( A => memory_20_7_port, Y => n429);
   U847 : MUX2X1 port map( B => n429, A => n158, S => n428, Y => n1359);
   U848 : MUX2X1 port map( B => n766, A => n144, S => n431, Y => n1496);
   U849 : MUX2X1 port map( B => n765, A => n146, S => n431, Y => n1495);
   U850 : MUX2X1 port map( B => n764, A => n148, S => n431, Y => n1494);
   U851 : MUX2X1 port map( B => n763, A => n150, S => n431, Y => n1493);
   U852 : MUX2X1 port map( B => n762, A => n152, S => n431, Y => n1492);
   U853 : MUX2X1 port map( B => n761, A => n540, S => n431, Y => n1491);
   U854 : MUX2X1 port map( B => n760, A => n156, S => n431, Y => n1490);
   U855 : MUX2X1 port map( B => n759, A => n159, S => n431, Y => n1489);
   U856 : MUX2X1 port map( B => n758, A => n144, S => n433, Y => n1488);
   U857 : MUX2X1 port map( B => n757, A => n146, S => n433, Y => n1487);
   U858 : MUX2X1 port map( B => n756, A => n148, S => n433, Y => n1486);
   U859 : MUX2X1 port map( B => n755, A => n150, S => n433, Y => n1485);
   U860 : MUX2X1 port map( B => n754, A => n152, S => n433, Y => n1484);
   U861 : MUX2X1 port map( B => n753, A => n540, S => n433, Y => n1483);
   U862 : MUX2X1 port map( B => n752, A => n156, S => n433, Y => n1482);
   U863 : MUX2X1 port map( B => n751, A => n159, S => n433, Y => n1481);
   U864 : MUX2X1 port map( B => n750, A => n144, S => n435, Y => n1480);
   U865 : MUX2X1 port map( B => n749, A => n146, S => n435, Y => n1479);
   U866 : MUX2X1 port map( B => n748, A => n148, S => n435, Y => n1478);
   U867 : MUX2X1 port map( B => n747, A => n150, S => n435, Y => n1477);
   U868 : MUX2X1 port map( B => n746, A => n152, S => n435, Y => n1476);
   U869 : MUX2X1 port map( B => n745, A => n540, S => n435, Y => n1475);
   U870 : MUX2X1 port map( B => n744, A => n156, S => n435, Y => n1474);
   U871 : MUX2X1 port map( B => n743, A => n159, S => n435, Y => n1473);
   U872 : MUX2X1 port map( B => n742, A => n144, S => n437, Y => n1472);
   U873 : MUX2X1 port map( B => n741, A => n146, S => n437, Y => n1471);
   U874 : MUX2X1 port map( B => n740, A => n148, S => n437, Y => n1470);
   U875 : MUX2X1 port map( B => n739, A => n150, S => n437, Y => n1469);
   U876 : MUX2X1 port map( B => n738, A => n152, S => n437, Y => n1468);
   U877 : MUX2X1 port map( B => n737, A => n540, S => n437, Y => n1467);
   U878 : MUX2X1 port map( B => n736, A => n156, S => n437, Y => n1466);
   U879 : MUX2X1 port map( B => n735, A => n159, S => n437, Y => n1465);
   U880 : INVX2 port map( A => memory_15_0_port, Y => n439);
   U881 : MUX2X1 port map( B => n439, A => n144, S => n446, Y => n1374);
   U882 : INVX2 port map( A => memory_15_1_port, Y => n440);
   U883 : MUX2X1 port map( B => n440, A => n146, S => n446, Y => n1373);
   U884 : INVX2 port map( A => memory_15_2_port, Y => n441);
   U885 : MUX2X1 port map( B => n441, A => n148, S => n446, Y => n1372);
   U886 : INVX2 port map( A => memory_15_3_port, Y => n442);
   U887 : MUX2X1 port map( B => n442, A => n150, S => n446, Y => n1371);
   U888 : INVX2 port map( A => memory_15_4_port, Y => n443);
   U889 : MUX2X1 port map( B => n443, A => n152, S => n446, Y => n1370);
   U890 : INVX2 port map( A => memory_15_5_port, Y => n444);
   U891 : MUX2X1 port map( B => n444, A => n540, S => n446, Y => n1369);
   U892 : INVX2 port map( A => memory_15_6_port, Y => n445);
   U893 : MUX2X1 port map( B => n445, A => n156, S => n446, Y => n1368);
   U894 : INVX2 port map( A => memory_15_7_port, Y => n447);
   U895 : MUX2X1 port map( B => n447, A => n159, S => n446, Y => n1367);
   U896 : INVX2 port map( A => memory_14_0_port, Y => n449);
   U897 : MUX2X1 port map( B => n449, A => n144, S => n456, Y => n1382);
   U898 : INVX2 port map( A => memory_14_1_port, Y => n450);
   U899 : MUX2X1 port map( B => n450, A => n536, S => n456, Y => n1381);
   U900 : INVX2 port map( A => memory_14_2_port, Y => n451);
   U901 : MUX2X1 port map( B => n451, A => n148, S => n456, Y => n1380);
   U902 : INVX2 port map( A => memory_14_3_port, Y => n452);
   U903 : MUX2X1 port map( B => n452, A => n150, S => n456, Y => n1379);
   U904 : INVX2 port map( A => memory_14_4_port, Y => n453);
   U905 : MUX2X1 port map( B => n453, A => n152, S => n456, Y => n1378);
   U906 : INVX2 port map( A => memory_14_5_port, Y => n454);
   U907 : MUX2X1 port map( B => n454, A => n540, S => n456, Y => n1377);
   U908 : INVX2 port map( A => memory_14_6_port, Y => n455);
   U909 : MUX2X1 port map( B => n455, A => n541, S => n456, Y => n1376);
   U910 : INVX2 port map( A => memory_14_7_port, Y => n457);
   U911 : MUX2X1 port map( B => n457, A => n159, S => n456, Y => n1375);
   U912 : INVX2 port map( A => memory_13_0_port, Y => n459);
   U913 : MUX2X1 port map( B => n459, A => n144, S => n466, Y => n1390);
   U914 : INVX2 port map( A => memory_13_1_port, Y => n460);
   U915 : MUX2X1 port map( B => n460, A => n536, S => n466, Y => n1389);
   U916 : INVX2 port map( A => memory_13_2_port, Y => n461);
   U917 : MUX2X1 port map( B => n461, A => n148, S => n466, Y => n1388);
   U918 : INVX2 port map( A => memory_13_3_port, Y => n462);
   U919 : MUX2X1 port map( B => n462, A => n150, S => n466, Y => n1387);
   U920 : INVX2 port map( A => memory_13_4_port, Y => n463);
   U921 : MUX2X1 port map( B => n463, A => n152, S => n466, Y => n1386);
   U922 : INVX2 port map( A => memory_13_5_port, Y => n464);
   U923 : MUX2X1 port map( B => n464, A => n540, S => n466, Y => n1385);
   U924 : INVX2 port map( A => memory_13_6_port, Y => n465);
   U925 : MUX2X1 port map( B => n465, A => n541, S => n466, Y => n1384);
   U926 : INVX2 port map( A => memory_13_7_port, Y => n467);
   U927 : MUX2X1 port map( B => n467, A => n159, S => n466, Y => n1383);
   U928 : INVX2 port map( A => memory_12_0_port, Y => n469);
   U929 : MUX2X1 port map( B => n469, A => n535, S => n476, Y => n1398);
   U930 : INVX2 port map( A => memory_12_1_port, Y => n470);
   U931 : MUX2X1 port map( B => n470, A => n536, S => n476, Y => n1397);
   U932 : INVX2 port map( A => memory_12_2_port, Y => n471);
   U933 : MUX2X1 port map( B => n471, A => n537, S => n476, Y => n1396);
   U934 : INVX2 port map( A => memory_12_3_port, Y => n472);
   U935 : MUX2X1 port map( B => n472, A => n538, S => n476, Y => n1395);
   U936 : INVX2 port map( A => memory_12_4_port, Y => n473);
   U937 : MUX2X1 port map( B => n473, A => n539, S => n476, Y => n1394);
   U938 : INVX2 port map( A => memory_12_5_port, Y => n474);
   U939 : MUX2X1 port map( B => n474, A => n154, S => n476, Y => n1393);
   U940 : INVX2 port map( A => memory_12_6_port, Y => n475);
   U941 : MUX2X1 port map( B => n475, A => n541, S => n476, Y => n1392);
   U942 : INVX2 port map( A => memory_12_7_port, Y => n477);
   U943 : MUX2X1 port map( B => n477, A => n159, S => n476, Y => n1391);
   U944 : NAND3X1 port map( A => n115, B => n160, C => n479, Y => n480);
   U945 : MUX2X1 port map( B => n734, A => n535, S => n481, Y => n1464);
   U946 : MUX2X1 port map( B => n733, A => n536, S => n481, Y => n1463);
   U947 : MUX2X1 port map( B => n732, A => n537, S => n481, Y => n1462);
   U948 : MUX2X1 port map( B => n731, A => n538, S => n481, Y => n1461);
   U949 : MUX2X1 port map( B => n730, A => n539, S => n481, Y => n1460);
   U950 : MUX2X1 port map( B => n729, A => n154, S => n481, Y => n1459);
   U951 : MUX2X1 port map( B => n728, A => n541, S => n481, Y => n1458);
   U952 : MUX2X1 port map( B => n727, A => n159, S => n481, Y => n1457);
   U953 : MUX2X1 port map( B => n726, A => n535, S => n483, Y => n1456);
   U954 : MUX2X1 port map( B => n725, A => n536, S => n483, Y => n1455);
   U955 : MUX2X1 port map( B => n724, A => n537, S => n483, Y => n1454);
   U956 : MUX2X1 port map( B => n723, A => n538, S => n483, Y => n1453);
   U957 : MUX2X1 port map( B => n722, A => n539, S => n483, Y => n1452);
   U958 : MUX2X1 port map( B => n721, A => n154, S => n483, Y => n1451);
   U959 : MUX2X1 port map( B => n720, A => n541, S => n483, Y => n1450);
   U960 : MUX2X1 port map( B => n719, A => n159, S => n483, Y => n1449);
   U961 : MUX2X1 port map( B => n718, A => n144, S => n485, Y => n1448);
   U962 : MUX2X1 port map( B => n717, A => n536, S => n485, Y => n1447);
   U963 : MUX2X1 port map( B => n716, A => n148, S => n485, Y => n1446);
   U964 : MUX2X1 port map( B => n715, A => n150, S => n485, Y => n1445);
   U965 : MUX2X1 port map( B => n714, A => n152, S => n485, Y => n1444);
   U966 : MUX2X1 port map( B => n713, A => n154, S => n485, Y => n1443);
   U967 : MUX2X1 port map( B => n712, A => n541, S => n485, Y => n1442);
   U968 : MUX2X1 port map( B => n711, A => n159, S => n485, Y => n1441);
   U969 : MUX2X1 port map( B => n710, A => n144, S => n487, Y => n1440);
   U970 : MUX2X1 port map( B => n709, A => n536, S => n487, Y => n1439);
   U971 : MUX2X1 port map( B => n708, A => n148, S => n487, Y => n1438);
   U972 : MUX2X1 port map( B => n707, A => n150, S => n487, Y => n1437);
   U973 : MUX2X1 port map( B => n706, A => n152, S => n487, Y => n1436);
   U974 : MUX2X1 port map( B => n705, A => n154, S => n487, Y => n1435);
   U975 : MUX2X1 port map( B => n704, A => n541, S => n487, Y => n1434);
   U976 : MUX2X1 port map( B => n703, A => n159, S => n487, Y => n1433);
   U977 : INVX2 port map( A => memory_7_0_port, Y => n489);
   U978 : MUX2X1 port map( B => n489, A => n535, S => n496, Y => n1565);
   U979 : INVX2 port map( A => memory_7_1_port, Y => n490);
   U980 : MUX2X1 port map( B => n490, A => n536, S => n496, Y => n1566);
   U981 : INVX2 port map( A => memory_7_2_port, Y => n491);
   U982 : MUX2X1 port map( B => n491, A => n537, S => n496, Y => n1567);
   U983 : INVX2 port map( A => memory_7_3_port, Y => n492);
   U984 : MUX2X1 port map( B => n492, A => n538, S => n496, Y => n1568);
   U985 : INVX2 port map( A => memory_7_4_port, Y => n493);
   U986 : MUX2X1 port map( B => n493, A => n539, S => n496, Y => n1569);
   U987 : INVX2 port map( A => memory_7_5_port, Y => n494);
   U988 : MUX2X1 port map( B => n494, A => n154, S => n496, Y => n1570);
   U989 : INVX2 port map( A => memory_7_6_port, Y => n495);
   U990 : MUX2X1 port map( B => n495, A => n541, S => n496, Y => n1571);
   U991 : INVX2 port map( A => memory_7_7_port, Y => n497);
   U992 : MUX2X1 port map( B => n497, A => n159, S => n496, Y => n1572);
   U993 : INVX2 port map( A => memory_6_0_port, Y => n499);
   U994 : MUX2X1 port map( B => n499, A => n535, S => n506, Y => n1575);
   U995 : INVX2 port map( A => memory_6_1_port, Y => n500);
   U996 : MUX2X1 port map( B => n500, A => n536, S => n506, Y => n1576);
   U997 : INVX2 port map( A => memory_6_2_port, Y => n501);
   U998 : MUX2X1 port map( B => n501, A => n537, S => n506, Y => n1577);
   U999 : INVX2 port map( A => memory_6_3_port, Y => n502);
   U1000 : MUX2X1 port map( B => n502, A => n538, S => n506, Y => n1578);
   U1001 : INVX2 port map( A => memory_6_4_port, Y => n503);
   U1002 : MUX2X1 port map( B => n503, A => n539, S => n506, Y => n1579);
   U1003 : INVX2 port map( A => memory_6_5_port, Y => n504);
   U1004 : MUX2X1 port map( B => n504, A => n154, S => n506, Y => n1580);
   U1005 : INVX2 port map( A => memory_6_6_port, Y => n505);
   U1006 : MUX2X1 port map( B => n505, A => n541, S => n506, Y => n1581);
   U1007 : INVX2 port map( A => memory_6_7_port, Y => n507);
   U1008 : MUX2X1 port map( B => n507, A => n158, S => n506, Y => n1582);
   U1009 : INVX2 port map( A => memory_5_0_port, Y => n509);
   U1010 : MUX2X1 port map( B => n509, A => n535, S => n516, Y => n1585);
   U1011 : INVX2 port map( A => memory_5_1_port, Y => n510);
   U1012 : MUX2X1 port map( B => n510, A => n536, S => n516, Y => n1586);
   U1013 : INVX2 port map( A => memory_5_2_port, Y => n511);
   U1014 : MUX2X1 port map( B => n511, A => n537, S => n516, Y => n1587);
   U1015 : INVX2 port map( A => memory_5_3_port, Y => n512);
   U1016 : MUX2X1 port map( B => n512, A => n538, S => n516, Y => n1588);
   U1017 : INVX2 port map( A => memory_5_4_port, Y => n513);
   U1018 : MUX2X1 port map( B => n513, A => n539, S => n516, Y => n1589);
   U1019 : INVX2 port map( A => memory_5_5_port, Y => n514);
   U1020 : MUX2X1 port map( B => n514, A => n154, S => n516, Y => n1590);
   U1021 : INVX2 port map( A => memory_5_6_port, Y => n515);
   U1022 : MUX2X1 port map( B => n515, A => n541, S => n516, Y => n1591);
   U1023 : INVX2 port map( A => memory_5_7_port, Y => n517);
   U1024 : MUX2X1 port map( B => n517, A => n159, S => n516, Y => n1592);
   U1025 : INVX2 port map( A => memory_4_0_port, Y => n519);
   U1026 : MUX2X1 port map( B => n519, A => n535, S => n526, Y => n1595);
   U1027 : INVX2 port map( A => memory_4_1_port, Y => n520);
   U1028 : MUX2X1 port map( B => n520, A => n536, S => n526, Y => n1596);
   U1029 : INVX2 port map( A => memory_4_2_port, Y => n521);
   U1030 : MUX2X1 port map( B => n521, A => n537, S => n526, Y => n1597);
   U1031 : INVX2 port map( A => memory_4_3_port, Y => n522);
   U1032 : MUX2X1 port map( B => n522, A => n538, S => n526, Y => n1598);
   U1033 : INVX2 port map( A => memory_4_4_port, Y => n523);
   U1034 : MUX2X1 port map( B => n523, A => n539, S => n526, Y => n1599);
   U1035 : INVX2 port map( A => memory_4_5_port, Y => n524);
   U1036 : MUX2X1 port map( B => n524, A => n154, S => n526, Y => n1600);
   U1037 : INVX2 port map( A => memory_4_6_port, Y => n525);
   U1038 : MUX2X1 port map( B => n525, A => n541, S => n526, Y => n1601);
   U1039 : INVX2 port map( A => memory_4_7_port, Y => n527);
   U1040 : MUX2X1 port map( B => n527, A => n158, S => n526, Y => n1602);
   U1041 : MUX2X1 port map( B => n693, A => n535, S => n529, Y => n1423);
   U1042 : MUX2X1 port map( B => n694, A => n146, S => n529, Y => n1424);
   U1043 : MUX2X1 port map( B => n695, A => n537, S => n529, Y => n1425);
   U1044 : MUX2X1 port map( B => n696, A => n538, S => n529, Y => n1426);
   U1045 : MUX2X1 port map( B => n697, A => n539, S => n529, Y => n1427);
   U1046 : MUX2X1 port map( B => n698, A => n154, S => n529, Y => n1428);
   U1047 : MUX2X1 port map( B => n699, A => n156, S => n529, Y => n1429);
   U1048 : MUX2X1 port map( B => n700, A => n159, S => n529, Y => n1430);
   U1049 : MUX2X1 port map( B => n685, A => n535, S => n531, Y => n1415);
   U1050 : MUX2X1 port map( B => n686, A => n146, S => n531, Y => n1416);
   U1051 : MUX2X1 port map( B => n687, A => n537, S => n531, Y => n1417);
   U1052 : MUX2X1 port map( B => n688, A => n538, S => n531, Y => n1418);
   U1053 : MUX2X1 port map( B => n689, A => n539, S => n531, Y => n1419);
   U1054 : MUX2X1 port map( B => n690, A => n154, S => n531, Y => n1420);
   U1055 : MUX2X1 port map( B => n691, A => n156, S => n531, Y => n1421);
   U1056 : MUX2X1 port map( B => n692, A => n158, S => n531, Y => n1422);
   U1057 : MUX2X1 port map( B => n677, A => n535, S => n533, Y => n1407);
   U1058 : MUX2X1 port map( B => n678, A => n146, S => n533, Y => n1408);
   U1059 : MUX2X1 port map( B => n679, A => n537, S => n533, Y => n1409);
   U1060 : MUX2X1 port map( B => n680, A => n538, S => n533, Y => n1410);
   U1061 : MUX2X1 port map( B => n681, A => n539, S => n533, Y => n1411);
   U1062 : MUX2X1 port map( B => n682, A => n154, S => n533, Y => n1412);
   U1063 : MUX2X1 port map( B => n683, A => n156, S => n533, Y => n1413);
   U1064 : MUX2X1 port map( B => n684, A => n159, S => n533, Y => n1414);
   U1065 : MUX2X1 port map( B => n669, A => n535, S => n542, Y => n1399);
   U1066 : MUX2X1 port map( B => n670, A => n146, S => n542, Y => n1400);
   U1067 : MUX2X1 port map( B => n671, A => n537, S => n542, Y => n1401);
   U1068 : MUX2X1 port map( B => n672, A => n538, S => n542, Y => n1402);
   U1069 : MUX2X1 port map( B => n673, A => n539, S => n542, Y => n1403);
   U1070 : MUX2X1 port map( B => n674, A => n154, S => n542, Y => n1404);
   U1071 : MUX2X1 port map( B => n675, A => n156, S => n542, Y => n1405);
   U1072 : MUX2X1 port map( B => n676, A => n158, S => n542, Y => n1406);
   U1073 : AND2X2 port map( A => state, B => n543, Y => N338);
   U1074 : XOR2X1 port map( A => n25, B => n88, Y => n544);
   U1075 : INVX2 port map( A => state, Y => n615);
   U1076 : NOR2X1 port map( A => n544, B => n615, Y => N339);
   U1077 : NAND2X1 port map( A => n130, B => n611, Y => n547);
   U1078 : OAI21X1 port map( A => n131, B => n611, C => n25, Y => n546);
   U1079 : AND2X2 port map( A => n547, B => n546, Y => n552);
   U1080 : XNOR2X1 port map( A => n552, B => n548, Y => n549);
   U1081 : AND2X2 port map( A => state, B => n549, Y => N340);
   U1082 : NOR2X1 port map( A => n70, B => n618, Y => n551);
   U1083 : NAND2X1 port map( A => n70, B => n618, Y => n550);
   U1084 : OAI21X1 port map( A => n552, B => n551, C => n550, Y => n556);
   U1085 : XNOR2X1 port map( A => n556, B => n553, Y => n554);
   U1086 : NOR2X1 port map( A => n554, B => n615, Y => N341);
   U1087 : NAND2X1 port map( A => n136, B => n587, Y => n557);
   U1088 : NOR2X1 port map( A => n136, B => n587, Y => n555);
   U1089 : AOI21X1 port map( A => n557, B => n556, C => n555, Y => n559);
   U1090 : XNOR2X1 port map( A => n559, B => n558, Y => n560);
   U1091 : AND2X2 port map( A => state, B => n560, Y => N342);
   U1092 : NOR2X1 port map( A => n41, B => n561, Y => n566);
   U1093 : AND2X2 port map( A => n563, B => n562, Y => n564);
   U1094 : NAND3X1 port map( A => n566, B => n565, C => n564, Y => n567);
   U1095 : MUX2X1 port map( B => n567, A => n701, S => RST, Y => n1431);
   U1096 : NAND2X1 port map( A => n56, B => n161, Y => n583);
   U1097 : INVX2 port map( A => n583, Y => n594);
   U1098 : NAND2X1 port map( A => n594, B => n54, Y => n574);
   U1099 : NAND2X1 port map( A => n29, B => n72, Y => n585);
   U1100 : INVX2 port map( A => n585, Y => n597);
   U1101 : NAND2X1 port map( A => n70, B => n577, Y => n570);
   U1102 : NAND2X1 port map( A => n570, B => n118, Y => n571);
   U1103 : NAND2X1 port map( A => n597, B => n571, Y => n573);
   U1104 : NAND2X1 port map( A => n70, B => n579, Y => n572);
   U1105 : NAND3X1 port map( A => n574, B => n573, C => n572, Y => n1614);
   U1106 : NAND2X1 port map( A => n594, B => n576, Y => n582);
   U1107 : NAND2X1 port map( A => n577, B => n28, Y => n578);
   U1108 : NAND2X1 port map( A => n597, B => n578, Y => n581);
   U1109 : NAND2X1 port map( A => n131, B => n579, Y => n580);
   U1110 : NAND3X1 port map( A => n582, B => n581, C => n580, Y => n1612);
   U1111 : AND2X2 port map( A => n585, B => n583, Y => n584);
   U1112 : MUX2X1 port map( B => n584, A => n56, S => n133, Y => n1610);
   U1113 : OAI21X1 port map( A => n6, B => n585, C => n56, Y => n596);
   U1114 : NAND2X1 port map( A => n100, B => n596, Y => n590);
   U1115 : NAND3X1 port map( A => n597, B => n6, C => n587, Y => n595);
   U1116 : XOR2X1 port map( A => n587, B => n31, Y => n588);
   U1117 : NAND2X1 port map( A => n588, B => n594, Y => n589);
   U1118 : NAND3X1 port map( A => n590, B => n595, C => n589, Y => n1608);
   U1119 : XOR2X1 port map( A => n48, B => n591, Y => n593);
   U1120 : NAND2X1 port map( A => n594, B => n593, Y => n603);
   U1121 : INVX2 port map( A => n595, Y => n601);
   U1122 : INVX2 port map( A => n596, Y => n599);
   U1123 : NAND2X1 port map( A => n597, B => n101, Y => n598);
   U1124 : NAND2X1 port map( A => n599, B => n598, Y => n600);
   U1125 : MUX2X1 port map( B => n601, A => n600, S => n52, Y => n602);
   U1126 : NAND2X1 port map( A => n603, B => n602, Y => n1607);
   U1127 : NAND2X1 port map( A => n87, B => n34, Y => n607);
   U1128 : INVX2 port map( A => n607, Y => n604);
   U1129 : NAND2X1 port map( A => n604, B => n136, Y => n605);
   U1130 : XNOR2X1 port map( A => n605, B => n620, Y => n606);
   U1131 : NOR2X1 port map( A => n615, B => n606, Y => N347);
   U1132 : XNOR2X1 port map( A => n607, B => n619, Y => n608);
   U1133 : NOR2X1 port map( A => n615, B => n608, Y => N346);
   U1134 : NAND2X1 port map( A => n86, B => n34, Y => n610);
   U1135 : OAI21X1 port map( A => n612, B => n611, C => n43, Y => n609);
   U1136 : AOI21X1 port map( A => n610, B => n609, C => n615, Y => N345);
   U1137 : XNOR2X1 port map( A => n612, B => n611, Y => n613);
   U1138 : NOR2X1 port map( A => n615, B => n613, Y => N344);
   U1139 : XNOR2X1 port map( A => n614, B => n57, Y => n616);
   U1140 : NOR2X1 port map( A => n616, B => n615, Y => N343);
   U1141 : INVX1 port map( A => FULL_port, Y => n701);
   U1142 : INVX1 port map( A => EMPTY_port, Y => n702);
   U1143 : NAND2X1 port map( A => n784, B => n785, Y => n783);
   U1144 : NOR2X1 port map( A => n786, B => n787, Y => n785);
   U1145 : NAND3X1 port map( A => n788, B => n789, C => n790, Y => n787);
   U1146 : NOR2X1 port map( A => n791, B => n792, Y => n790);
   U1147 : OAI22X1 port map( A => n735, B => n121, C => n743, D => n120, Y => 
                           n792);
   U1148 : OAI22X1 port map( A => n751, B => n102, C => n759, D => n104, Y => 
                           n791);
   U1149 : AOI22X1 port map( A => n79, B => memory_23_7_port, C => n75, D => 
                           memory_22_7_port, Y => n789);
   U1150 : AOI22X1 port map( A => n795, B => memory_21_7_port, C => n796, D => 
                           memory_20_7_port, Y => n788);
   U1151 : NAND3X1 port map( A => n797, B => n798, C => n799, Y => n786);
   U1152 : NOR2X1 port map( A => n800, B => n801, Y => n799);
   U1153 : OAI22X1 port map( A => n661, B => n123, C => n653, D => n122, Y => 
                           n801);
   U1154 : OAI22X1 port map( A => n645, B => n105, C => n637, D => n107, Y => 
                           n800);
   U1155 : AOI22X1 port map( A => n80, B => memory_31_7_port, C => n77, D => 
                           memory_30_7_port, Y => n798);
   U1156 : AOI22X1 port map( A => n803, B => memory_29_7_port, C => n804, D => 
                           memory_28_7_port, Y => n797);
   U1157 : NOR2X1 port map( A => n805, B => n806, Y => n784);
   U1158 : NAND3X1 port map( A => n807, B => n808, C => n809, Y => n806);
   U1159 : NOR2X1 port map( A => n810, B => n811, Y => n809);
   U1160 : OAI22X1 port map( A => n700, B => n108, C => n692, D => n110, Y => 
                           n811);
   U1161 : OAI22X1 port map( A => n684, B => n125, C => n676, D => n124, Y => 
                           n810);
   U1162 : AOI22X1 port map( A => n813, B => memory_4_7_port, C => n814, D => 
                           memory_5_7_port, Y => n808);
   U1163 : AOI22X1 port map( A => n81, B => memory_6_7_port, C => n76, D => 
                           memory_7_7_port, Y => n807);
   U1164 : NAND3X1 port map( A => n815, B => n816, C => n817, Y => n805);
   U1165 : NOR2X1 port map( A => n818, B => n819, Y => n817);
   U1166 : OAI22X1 port map( A => n703, B => n127, C => n711, D => n126, Y => 
                           n819);
   U1167 : OAI22X1 port map( A => n719, B => n111, C => n727, D => n112, Y => 
                           n818);
   U1168 : AOI22X1 port map( A => n78, B => memory_15_7_port, C => n74, D => 
                           memory_14_7_port, Y => n816);
   U1169 : AOI22X1 port map( A => n820, B => memory_13_7_port, C => n821, D => 
                           memory_12_7_port, Y => n815);
   U1170 : NAND2X1 port map( A => n823, B => n824, Y => n822);
   U1171 : NOR2X1 port map( A => n825, B => n826, Y => n824);
   U1172 : NAND3X1 port map( A => n827, B => n828, C => n829, Y => n826);
   U1173 : NOR2X1 port map( A => n830, B => n831, Y => n829);
   U1174 : OAI22X1 port map( A => n736, B => n121, C => n744, D => n120, Y => 
                           n831);
   U1175 : OAI22X1 port map( A => n752, B => n102, C => n760, D => n104, Y => 
                           n830);
   U1176 : AOI22X1 port map( A => n79, B => memory_23_6_port, C => n75, D => 
                           memory_22_6_port, Y => n828);
   U1177 : AOI22X1 port map( A => n795, B => memory_21_6_port, C => n796, D => 
                           memory_20_6_port, Y => n827);
   U1178 : NAND3X1 port map( A => n832, B => n833, C => n834, Y => n825);
   U1179 : NOR2X1 port map( A => n835, B => n836, Y => n834);
   U1180 : OAI22X1 port map( A => n662, B => n123, C => n654, D => n122, Y => 
                           n836);
   U1181 : OAI22X1 port map( A => n646, B => n105, C => n638, D => n107, Y => 
                           n835);
   U1182 : AOI22X1 port map( A => n80, B => memory_31_6_port, C => n77, D => 
                           memory_30_6_port, Y => n833);
   U1183 : AOI22X1 port map( A => n803, B => memory_29_6_port, C => n804, D => 
                           memory_28_6_port, Y => n832);
   U1184 : NOR2X1 port map( A => n837, B => n838, Y => n823);
   U1185 : NAND3X1 port map( A => n839, B => n840, C => n841, Y => n838);
   U1186 : NOR2X1 port map( A => n842, B => n843, Y => n841);
   U1187 : OAI22X1 port map( A => n699, B => n108, C => n691, D => n110, Y => 
                           n843);
   U1188 : OAI22X1 port map( A => n683, B => n125, C => n675, D => n124, Y => 
                           n842);
   U1189 : AOI22X1 port map( A => n813, B => memory_4_6_port, C => n814, D => 
                           memory_5_6_port, Y => n840);
   U1190 : AOI22X1 port map( A => n81, B => memory_6_6_port, C => n76, D => 
                           memory_7_6_port, Y => n839);
   U1200 : NAND3X1 port map( A => n844, B => n845, C => n846, Y => n837);
   U1201 : NOR2X1 port map( A => n852, B => n861, Y => n846);
   U1203 : OAI22X1 port map( A => n704, B => n127, C => n712, D => n126, Y => 
                           n861);
   U1207 : OAI22X1 port map( A => n720, B => n111, C => n728, D => n112, Y => 
                           n852);
   U1208 : AOI22X1 port map( A => n78, B => memory_15_6_port, C => n74, D => 
                           memory_14_6_port, Y => n845);
   U1209 : AOI22X1 port map( A => n820, B => memory_13_6_port, C => n821, D => 
                           memory_12_6_port, Y => n844);
   U1210 : NAND2X1 port map( A => n865, B => n909, Y => n863);
   U1211 : NOR2X1 port map( A => n910, B => n911, Y => n909);
   U1212 : NAND3X1 port map( A => n912, B => n913, C => n914, Y => n911);
   U1213 : NOR2X1 port map( A => n915, B => n916, Y => n914);
   U1214 : OAI22X1 port map( A => n737, B => n121, C => n745, D => n120, Y => 
                           n916);
   U1215 : OAI22X1 port map( A => n753, B => n102, C => n761, D => n104, Y => 
                           n915);
   U1216 : AOI22X1 port map( A => n79, B => memory_23_5_port, C => n75, D => 
                           memory_22_5_port, Y => n913);
   U1217 : AOI22X1 port map( A => n795, B => memory_21_5_port, C => n796, D => 
                           memory_20_5_port, Y => n912);
   U1218 : NAND3X1 port map( A => n917, B => n918, C => n919, Y => n910);
   U1219 : NOR2X1 port map( A => n920, B => n921, Y => n919);
   U1220 : OAI22X1 port map( A => n663, B => n123, C => n655, D => n122, Y => 
                           n921);
   U1221 : OAI22X1 port map( A => n647, B => n105, C => n639, D => n107, Y => 
                           n920);
   U1222 : AOI22X1 port map( A => n80, B => memory_31_5_port, C => n77, D => 
                           memory_30_5_port, Y => n918);
   U1223 : AOI22X1 port map( A => n803, B => memory_29_5_port, C => n804, D => 
                           memory_28_5_port, Y => n917);
   U1224 : NOR2X1 port map( A => n922, B => n923, Y => n865);
   U1225 : NAND3X1 port map( A => n924, B => n925, C => n926, Y => n923);
   U1226 : NOR2X1 port map( A => n927, B => n928, Y => n926);
   U1227 : OAI22X1 port map( A => n698, B => n108, C => n690, D => n110, Y => 
                           n928);
   U1228 : OAI22X1 port map( A => n682, B => n125, C => n674, D => n124, Y => 
                           n927);
   U1229 : AOI22X1 port map( A => n813, B => memory_4_5_port, C => n814, D => 
                           memory_5_5_port, Y => n925);
   U1230 : AOI22X1 port map( A => n81, B => memory_6_5_port, C => n76, D => 
                           memory_7_5_port, Y => n924);
   U1231 : NAND3X1 port map( A => n929, B => n930, C => n931, Y => n922);
   U1232 : NOR2X1 port map( A => n932, B => n933, Y => n931);
   U1233 : OAI22X1 port map( A => n705, B => n127, C => n713, D => n126, Y => 
                           n933);
   U1234 : OAI22X1 port map( A => n721, B => n111, C => n729, D => n112, Y => 
                           n932);
   U1235 : AOI22X1 port map( A => n78, B => memory_15_5_port, C => n74, D => 
                           memory_14_5_port, Y => n930);
   U1236 : AOI22X1 port map( A => n820, B => memory_13_5_port, C => n821, D => 
                           memory_12_5_port, Y => n929);
   U1237 : NAND2X1 port map( A => n935, B => n936, Y => n934);
   U1238 : NOR2X1 port map( A => n937, B => n938, Y => n936);
   U1239 : NAND3X1 port map( A => n939, B => n940, C => n941, Y => n938);
   U1240 : NOR2X1 port map( A => n942, B => n943, Y => n941);
   U1241 : OAI22X1 port map( A => n738, B => n121, C => n746, D => n120, Y => 
                           n943);
   U1242 : OAI22X1 port map( A => n754, B => n102, C => n762, D => n104, Y => 
                           n942);
   U1243 : AOI22X1 port map( A => n79, B => memory_23_4_port, C => n75, D => 
                           memory_22_4_port, Y => n940);
   U1244 : AOI22X1 port map( A => n795, B => memory_21_4_port, C => n796, D => 
                           memory_20_4_port, Y => n939);
   U1245 : NAND3X1 port map( A => n944, B => n945, C => n946, Y => n937);
   U1246 : NOR2X1 port map( A => n947, B => n948, Y => n946);
   U1247 : OAI22X1 port map( A => n664, B => n123, C => n656, D => n122, Y => 
                           n948);
   U1248 : OAI22X1 port map( A => n648, B => n105, C => n640, D => n107, Y => 
                           n947);
   U1249 : AOI22X1 port map( A => n80, B => memory_31_4_port, C => n77, D => 
                           memory_30_4_port, Y => n945);
   U1250 : AOI22X1 port map( A => n803, B => memory_29_4_port, C => n804, D => 
                           memory_28_4_port, Y => n944);
   U1251 : NOR2X1 port map( A => n949, B => n950, Y => n935);
   U1252 : NAND3X1 port map( A => n951, B => n952, C => n953, Y => n950);
   U1253 : NOR2X1 port map( A => n954, B => n955, Y => n953);
   U1254 : OAI22X1 port map( A => n697, B => n108, C => n689, D => n110, Y => 
                           n955);
   U1255 : OAI22X1 port map( A => n681, B => n125, C => n673, D => n124, Y => 
                           n954);
   U1256 : AOI22X1 port map( A => n813, B => memory_4_4_port, C => n814, D => 
                           memory_5_4_port, Y => n952);
   U1257 : AOI22X1 port map( A => n81, B => memory_6_4_port, C => n76, D => 
                           memory_7_4_port, Y => n951);
   U1258 : NAND3X1 port map( A => n956, B => n957, C => n958, Y => n949);
   U1259 : NOR2X1 port map( A => n959, B => n960, Y => n958);
   U1260 : OAI22X1 port map( A => n706, B => n127, C => n714, D => n126, Y => 
                           n960);
   U1261 : OAI22X1 port map( A => n722, B => n111, C => n730, D => n112, Y => 
                           n959);
   U1262 : AOI22X1 port map( A => n78, B => memory_15_4_port, C => n74, D => 
                           memory_14_4_port, Y => n957);
   U1263 : AOI22X1 port map( A => n820, B => memory_13_4_port, C => n821, D => 
                           memory_12_4_port, Y => n956);
   U1264 : NAND2X1 port map( A => n962, B => n963, Y => n961);
   U1265 : NOR2X1 port map( A => n964, B => n965, Y => n963);
   U1266 : NAND3X1 port map( A => n966, B => n967, C => n968, Y => n965);
   U1267 : NOR2X1 port map( A => n969, B => n970, Y => n968);
   U1268 : OAI22X1 port map( A => n739, B => n121, C => n747, D => n120, Y => 
                           n970);
   U1269 : OAI22X1 port map( A => n755, B => n102, C => n763, D => n104, Y => 
                           n969);
   U1270 : AOI22X1 port map( A => n79, B => memory_23_3_port, C => n75, D => 
                           memory_22_3_port, Y => n967);
   U1271 : AOI22X1 port map( A => n795, B => memory_21_3_port, C => n796, D => 
                           memory_20_3_port, Y => n966);
   U1272 : NAND3X1 port map( A => n971, B => n972, C => n973, Y => n964);
   U1273 : NOR2X1 port map( A => n974, B => n975, Y => n973);
   U1274 : OAI22X1 port map( A => n665, B => n123, C => n657, D => n122, Y => 
                           n975);
   U1275 : OAI22X1 port map( A => n649, B => n105, C => n641, D => n107, Y => 
                           n974);
   U1276 : AOI22X1 port map( A => n80, B => memory_31_3_port, C => n77, D => 
                           memory_30_3_port, Y => n972);
   U1277 : AOI22X1 port map( A => n803, B => memory_29_3_port, C => n804, D => 
                           memory_28_3_port, Y => n971);
   U1278 : NOR2X1 port map( A => n976, B => n977, Y => n962);
   U1279 : NAND3X1 port map( A => n978, B => n979, C => n980, Y => n977);
   U1280 : NOR2X1 port map( A => n981, B => n982, Y => n980);
   U1281 : OAI22X1 port map( A => n696, B => n108, C => n688, D => n110, Y => 
                           n982);
   U1282 : OAI22X1 port map( A => n680, B => n125, C => n672, D => n124, Y => 
                           n981);
   U1283 : AOI22X1 port map( A => n813, B => memory_4_3_port, C => n814, D => 
                           memory_5_3_port, Y => n979);
   U1284 : AOI22X1 port map( A => n81, B => memory_6_3_port, C => n76, D => 
                           memory_7_3_port, Y => n978);
   U1285 : NAND3X1 port map( A => n983, B => n984, C => n985, Y => n976);
   U1286 : NOR2X1 port map( A => n986, B => n987, Y => n985);
   U1287 : OAI22X1 port map( A => n707, B => n127, C => n715, D => n126, Y => 
                           n987);
   U1288 : OAI22X1 port map( A => n723, B => n111, C => n731, D => n112, Y => 
                           n986);
   U1289 : AOI22X1 port map( A => n78, B => memory_15_3_port, C => n74, D => 
                           memory_14_3_port, Y => n984);
   U1290 : AOI22X1 port map( A => n820, B => memory_13_3_port, C => n821, D => 
                           memory_12_3_port, Y => n983);
   U1291 : NAND2X1 port map( A => n989, B => n990, Y => n988);
   U1292 : NOR2X1 port map( A => n991, B => n992, Y => n990);
   U1293 : NAND3X1 port map( A => n993, B => n994, C => n995, Y => n992);
   U1294 : NOR2X1 port map( A => n996, B => n997, Y => n995);
   U1295 : OAI22X1 port map( A => n740, B => n121, C => n748, D => n120, Y => 
                           n997);
   U1296 : OAI22X1 port map( A => n756, B => n102, C => n764, D => n104, Y => 
                           n996);
   U1297 : AOI22X1 port map( A => n79, B => memory_23_2_port, C => n75, D => 
                           memory_22_2_port, Y => n994);
   U1298 : AOI22X1 port map( A => n795, B => memory_21_2_port, C => n796, D => 
                           memory_20_2_port, Y => n993);
   U1299 : NAND3X1 port map( A => n998, B => n999, C => n1000, Y => n991);
   U1300 : NOR2X1 port map( A => n1001, B => n1002, Y => n1000);
   U1301 : OAI22X1 port map( A => n666, B => n123, C => n658, D => n122, Y => 
                           n1002);
   U1302 : OAI22X1 port map( A => n650, B => n105, C => n642, D => n107, Y => 
                           n1001);
   U1303 : AOI22X1 port map( A => n80, B => memory_31_2_port, C => n77, D => 
                           memory_30_2_port, Y => n999);
   U1304 : AOI22X1 port map( A => n803, B => memory_29_2_port, C => n804, D => 
                           memory_28_2_port, Y => n998);
   U1305 : NOR2X1 port map( A => n1003, B => n1004, Y => n989);
   U1306 : NAND3X1 port map( A => n1005, B => n1006, C => n1007, Y => n1004);
   U1307 : NOR2X1 port map( A => n1008, B => n1009, Y => n1007);
   U1308 : OAI22X1 port map( A => n695, B => n108, C => n687, D => n110, Y => 
                           n1009);
   U1309 : OAI22X1 port map( A => n679, B => n125, C => n671, D => n124, Y => 
                           n1008);
   U1310 : AOI22X1 port map( A => n813, B => memory_4_2_port, C => n814, D => 
                           memory_5_2_port, Y => n1006);
   U1311 : AOI22X1 port map( A => n81, B => memory_6_2_port, C => n76, D => 
                           memory_7_2_port, Y => n1005);
   U1312 : NAND3X1 port map( A => n1010, B => n1011, C => n1012, Y => n1003);
   U1313 : NOR2X1 port map( A => n1013, B => n1014, Y => n1012);
   U1314 : OAI22X1 port map( A => n708, B => n127, C => n716, D => n126, Y => 
                           n1014);
   U1315 : OAI22X1 port map( A => n724, B => n111, C => n732, D => n112, Y => 
                           n1013);
   U1316 : AOI22X1 port map( A => n78, B => memory_15_2_port, C => n74, D => 
                           memory_14_2_port, Y => n1011);
   U1317 : AOI22X1 port map( A => n820, B => memory_13_2_port, C => n821, D => 
                           memory_12_2_port, Y => n1010);
   U1318 : NAND2X1 port map( A => n1016, B => n1017, Y => n1015);
   U1319 : NOR2X1 port map( A => n1018, B => n1019, Y => n1017);
   U1320 : NAND3X1 port map( A => n1020, B => n1021, C => n1022, Y => n1019);
   U1321 : NOR2X1 port map( A => n1023, B => n1024, Y => n1022);
   U1322 : OAI22X1 port map( A => n741, B => n121, C => n749, D => n120, Y => 
                           n1024);
   U1323 : OAI22X1 port map( A => n757, B => n102, C => n765, D => n104, Y => 
                           n1023);
   U1324 : AOI22X1 port map( A => n79, B => memory_23_1_port, C => n75, D => 
                           memory_22_1_port, Y => n1021);
   U1325 : AOI22X1 port map( A => n795, B => memory_21_1_port, C => n796, D => 
                           memory_20_1_port, Y => n1020);
   U1326 : NAND3X1 port map( A => n1025, B => n1026, C => n1027, Y => n1018);
   U1327 : NOR2X1 port map( A => n1028, B => n1029, Y => n1027);
   U1328 : OAI22X1 port map( A => n667, B => n123, C => n659, D => n122, Y => 
                           n1029);
   U1329 : OAI22X1 port map( A => n651, B => n105, C => n643, D => n107, Y => 
                           n1028);
   U1330 : AOI22X1 port map( A => n80, B => memory_31_1_port, C => n77, D => 
                           memory_30_1_port, Y => n1026);
   U1331 : AOI22X1 port map( A => n803, B => memory_29_1_port, C => n804, D => 
                           memory_28_1_port, Y => n1025);
   U1332 : NOR2X1 port map( A => n1064, B => n1065, Y => n1016);
   U1333 : NAND3X1 port map( A => n1066, B => n1067, C => n1068, Y => n1065);
   U1334 : NOR2X1 port map( A => n1069, B => n1070, Y => n1068);
   U1335 : OAI22X1 port map( A => n694, B => n108, C => n686, D => n110, Y => 
                           n1070);
   U1336 : OAI22X1 port map( A => n678, B => n125, C => n670, D => n124, Y => 
                           n1069);
   U1337 : AOI22X1 port map( A => n813, B => memory_4_1_port, C => n814, D => 
                           memory_5_1_port, Y => n1067);
   U1338 : AOI22X1 port map( A => n81, B => memory_6_1_port, C => n76, D => 
                           memory_7_1_port, Y => n1066);
   U1339 : NAND3X1 port map( A => n1071, B => n1168, C => n1169, Y => n1064);
   U1340 : NOR2X1 port map( A => n1170, B => n1171, Y => n1169);
   U1341 : OAI22X1 port map( A => n709, B => n127, C => n717, D => n126, Y => 
                           n1171);
   U1342 : OAI22X1 port map( A => n725, B => n111, C => n733, D => n112, Y => 
                           n1170);
   U1343 : AOI22X1 port map( A => n78, B => memory_15_1_port, C => n74, D => 
                           memory_14_1_port, Y => n1168);
   U1344 : AOI22X1 port map( A => n820, B => memory_13_1_port, C => n821, D => 
                           memory_12_1_port, Y => n1071);
   U1345 : NAND2X1 port map( A => n1173, B => n1174, Y => n1172);
   U1346 : NOR2X1 port map( A => n1175, B => n1176, Y => n1174);
   U1347 : NAND3X1 port map( A => n1177, B => n1178, C => n1179, Y => n1176);
   U1348 : NOR2X1 port map( A => n1180, B => n1181, Y => n1179);
   U1349 : OAI22X1 port map( A => n742, B => n121, C => n750, D => n120, Y => 
                           n1181);
   U1350 : OAI22X1 port map( A => n758, B => n102, C => n766, D => n104, Y => 
                           n1180);
   U1351 : AOI22X1 port map( A => n79, B => memory_23_0_port, C => n75, D => 
                           memory_22_0_port, Y => n1178);
   U1352 : AOI22X1 port map( A => n795, B => memory_21_0_port, C => n796, D => 
                           memory_20_0_port, Y => n1177);
   U1353 : NAND3X1 port map( A => n1182, B => n1183, C => n1184, Y => n1175);
   U1354 : NOR2X1 port map( A => n1185, B => n1186, Y => n1184);
   U1355 : OAI22X1 port map( A => n668, B => n123, C => n660, D => n122, Y => 
                           n1186);
   U1356 : OAI22X1 port map( A => n652, B => n105, C => n644, D => n107, Y => 
                           n1185);
   U1357 : AOI22X1 port map( A => n80, B => memory_31_0_port, C => n77, D => 
                           memory_30_0_port, Y => n1183);
   U1358 : AOI22X1 port map( A => n803, B => memory_29_0_port, C => n804, D => 
                           memory_28_0_port, Y => n1182);
   U1359 : NOR2X1 port map( A => n1187, B => n1188, Y => n1173);
   U1360 : NAND3X1 port map( A => n1189, B => n1190, C => n1191, Y => n1188);
   U1361 : NOR2X1 port map( A => n1192, B => n1193, Y => n1191);
   U1362 : OAI22X1 port map( A => n693, B => n108, C => n685, D => n110, Y => 
                           n1193);
   U1363 : OAI22X1 port map( A => n677, B => n125, C => n669, D => n124, Y => 
                           n1192);
   U1364 : AOI22X1 port map( A => n813, B => memory_4_0_port, C => n814, D => 
                           memory_5_0_port, Y => n1190);
   U1365 : AOI22X1 port map( A => n81, B => memory_6_0_port, C => n76, D => 
                           memory_7_0_port, Y => n1189);
   U1366 : NAND3X1 port map( A => n1194, B => n1195, C => n1196, Y => n1187);
   U1367 : NOR2X1 port map( A => n1197, B => n1198, Y => n1196);
   U1368 : OAI22X1 port map( A => n710, B => n127, C => n718, D => n126, Y => 
                           n1198);
   U1369 : OAI22X1 port map( A => n726, B => n111, C => n734, D => n112, Y => 
                           n1197);
   U1370 : AOI22X1 port map( A => n78, B => memory_15_0_port, C => n74, D => 
                           memory_14_0_port, Y => n1195);
   U1371 : AOI22X1 port map( A => n820, B => memory_13_0_port, C => n821, D => 
                           memory_12_0_port, Y => n1194);
   U1372 : NAND2X1 port map( A => n1200, B => n1201, Y => n1199);
   U1373 : NOR2X1 port map( A => n1202, B => n1203, Y => n1201);
   U1374 : NAND3X1 port map( A => n1204, B => n1205, C => n1206, Y => n1203);
   U1375 : NOR2X1 port map( A => n1207, B => n1208, Y => n1206);
   U1376 : OAI22X1 port map( A => n775, B => n121, C => n777, D => n120, Y => 
                           n1208);
   U1377 : OAI22X1 port map( A => n779, B => n102, C => n781, D => n104, Y => 
                           n1207);
   U1378 : AOI22X1 port map( A => n79, B => opcode_23_1_port, C => n75, D => 
                           opcode_22_1_port, Y => n1205);
   U1379 : AOI22X1 port map( A => n795, B => opcode_21_1_port, C => n796, D => 
                           opcode_20_1_port, Y => n1204);
   U1380 : NAND3X1 port map( A => n1209, B => n1210, C => n1211, Y => n1202);
   U1381 : NOR2X1 port map( A => n1212, B => n1213, Y => n1211);
   U1382 : OAI22X1 port map( A => n627, B => n123, C => n625, D => n122, Y => 
                           n1213);
   U1383 : OAI22X1 port map( A => n623, B => n105, C => n621, D => n107, Y => 
                           n1212);
   U1384 : AOI22X1 port map( A => n80, B => opcode_31_1_port, C => n77, D => 
                           opcode_30_1_port, Y => n1210);
   U1385 : AOI22X1 port map( A => n803, B => opcode_29_1_port, C => n804, D => 
                           opcode_28_1_port, Y => n1209);
   U1386 : NOR2X1 port map( A => n1214, B => n1215, Y => n1200);
   U1387 : NAND3X1 port map( A => n1216, B => n1217, C => n1218, Y => n1215);
   U1388 : NOR2X1 port map( A => n1219, B => n1220, Y => n1218);
   U1389 : OAI22X1 port map( A => n636, B => n108, C => n634, D => n110, Y => 
                           n1220);
   U1390 : OAI22X1 port map( A => n632, B => n125, C => n630, D => n124, Y => 
                           n1219);
   U1391 : AOI22X1 port map( A => n813, B => opcode_4_1_port, C => n814, D => 
                           opcode_5_1_port, Y => n1217);
   U1392 : AOI22X1 port map( A => n81, B => opcode_6_1_port, C => n76, D => 
                           opcode_7_1_port, Y => n1216);
   U1393 : NAND3X1 port map( A => n1221, B => n1222, C => n1223, Y => n1214);
   U1394 : NOR2X1 port map( A => n1224, B => n1225, Y => n1223);
   U1395 : OAI22X1 port map( A => n767, B => n127, C => n769, D => n126, Y => 
                           n1225);
   U1396 : OAI22X1 port map( A => n771, B => n111, C => n773, D => n112, Y => 
                           n1224);
   U1397 : AOI22X1 port map( A => n78, B => opcode_15_1_port, C => n74, D => 
                           opcode_14_1_port, Y => n1222);
   U1398 : AOI22X1 port map( A => n820, B => opcode_13_1_port, C => n821, D => 
                           opcode_12_1_port, Y => n1221);
   U1399 : NAND2X1 port map( A => n1227, B => n1228, Y => n1226);
   U1400 : NOR2X1 port map( A => n1229, B => n1230, Y => n1228);
   U1401 : NAND3X1 port map( A => n1231, B => n1232, C => n1233, Y => n1230);
   U1402 : NOR2X1 port map( A => n1234, B => n1235, Y => n1233);
   U1403 : OAI22X1 port map( A => n776, B => n121, C => n778, D => n120, Y => 
                           n1235);
   U1404 : NAND2X1 port map( A => n1236, B => n1237, Y => n793);
   U1405 : OAI22X1 port map( A => n780, B => n102, C => n782, D => n104, Y => 
                           n1234);
   U1406 : AOI22X1 port map( A => n79, B => opcode_23_0_port, C => n75, D => 
                           opcode_22_0_port, Y => n1232);
   U1407 : AOI22X1 port map( A => n795, B => opcode_21_0_port, C => n796, D => 
                           opcode_20_0_port, Y => n1231);
   U1408 : INVX1 port map( A => n1240, Y => n1238);
   U1409 : NAND3X1 port map( A => n57, B => n619, C => n53, Y => n1240);
   U1410 : INVX1 port map( A => n1241, Y => n1236);
   U1411 : NAND3X1 port map( A => n50, B => n619, C => n53, Y => n1241);
   U1412 : NAND3X1 port map( A => n1242, B => n1243, C => n1244, Y => n1229);
   U1413 : NOR2X1 port map( A => n1245, B => n1246, Y => n1244);
   U1414 : OAI22X1 port map( A => n628, B => n123, C => n626, D => n122, Y => 
                           n1246);
   U1415 : OAI22X1 port map( A => n624, B => n105, C => n622, D => n107, Y => 
                           n1245);
   U1416 : AOI22X1 port map( A => n80, B => opcode_31_0_port, C => n77, D => 
                           opcode_30_0_port, Y => n1243);
   U1417 : AOI22X1 port map( A => n803, B => opcode_29_0_port, C => n804, D => 
                           opcode_28_0_port, Y => n1242);
   U1418 : INVX1 port map( A => n1249, Y => n1248);
   U1419 : NAND3X1 port map( A => n136, B => n617, C => n53, Y => n1249);
   U1420 : INVX1 port map( A => n1250, Y => n1247);
   U1421 : NAND3X1 port map( A => n136, B => n50, C => n53, Y => n1250);
   U1422 : NOR2X1 port map( A => n1251, B => n1252, Y => n1227);
   U1423 : NAND3X1 port map( A => n1253, B => n1254, C => n1255, Y => n1252);
   U1424 : NOR2X1 port map( A => n1256, B => n1257, Y => n1255);
   U1425 : OAI22X1 port map( A => n635, B => n108, C => n633, D => n110, Y => 
                           n1257);
   U1426 : OAI22X1 port map( A => n631, B => n125, C => n629, D => n124, Y => 
                           n1256);
   U1427 : AOI22X1 port map( A => n813, B => opcode_4_0_port, C => n814, D => 
                           opcode_5_0_port, Y => n1254);
   U1428 : AOI22X1 port map( A => n81, B => opcode_6_0_port, C => n76, D => 
                           opcode_7_0_port, Y => n1253);
   U1429 : INVX1 port map( A => n1260, Y => n1259);
   U1430 : NAND3X1 port map( A => n619, B => n620, C => n50, Y => n1260);
   U1431 : INVX1 port map( A => n1261, Y => n1258);
   U1432 : NAND3X1 port map( A => n619, B => n620, C => n57, Y => n1261);
   U1433 : NAND3X1 port map( A => n1262, B => n1263, C => n1264, Y => n1251);
   U1434 : NOR2X1 port map( A => n1265, B => n1266, Y => n1264);
   U1435 : OAI22X1 port map( A => n768, B => n127, C => n770, D => n126, Y => 
                           n1266);
   U1436 : NOR2X1 port map( A => n49, B => n43, Y => n1237);
   U1437 : OAI22X1 port map( A => n772, B => n111, C => n774, D => n112, Y => 
                           n1265);
   U1438 : AOI22X1 port map( A => n78, B => opcode_15_0_port, C => n74, D => 
                           opcode_14_0_port, Y => n1263);
   U1439 : AOI22X1 port map( A => n820, B => opcode_13_0_port, C => n821, D => 
                           opcode_12_0_port, Y => n1262);
   U1440 : INVX1 port map( A => n1269, Y => n1268);
   U1441 : NAND3X1 port map( A => n57, B => n620, C => n136, Y => n1269);
   U1442 : NOR2X1 port map( A => n618, B => n49, Y => n1239);
   U1443 : INVX1 port map( A => n1270, Y => n1267);
   U1444 : NAND3X1 port map( A => n50, B => n620, C => n136, Y => n1270);

end SYN_BRFIFO;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RBUFFER_0 is

   port( CLK, RST, NEXT_BYTE : in std_logic;  DATA : in std_logic_vector (7 
         downto 0);  OPCODE : in std_logic_vector (1 downto 0);  BYTE_COUNT : 
         in std_logic_vector (4 downto 0);  EOP : in std_logic;  B_READY, 
         R_ENABLE : out std_logic;  PRGA_IN : out std_logic_vector (7 downto 0)
         ;  PRGA_OPCODE : out std_logic_vector (1 downto 0));

end RBUFFER_0;

architecture SYN_brbuffer of RBUFFER_0 is

   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal B_READY_port, R_ENABLE_port, PRGA_IN_7_port, PRGA_IN_6_port, 
      PRGA_IN_5_port, PRGA_IN_4_port, PRGA_IN_3_port, PRGA_IN_2_port, 
      PRGA_IN_1_port, PRGA_IN_0_port, PRGA_OPCODE_1_port, PRGA_OPCODE_0_port, 
      state_2_port, state_1_port, state_0_port, nextState_2_port, 
      nextState_1_port, nextState_0_port, tempData_7_port, tempData_6_port, 
      tempData_5_port, tempData_4_port, tempData_3_port, tempData_2_port, 
      tempData_1_port, tempData_0_port, tempOpcode_1_port, tempOpcode_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103 : std_logic;

begin
   B_READY <= B_READY_port;
   R_ENABLE <= R_ENABLE_port;
   PRGA_IN <= ( PRGA_IN_7_port, PRGA_IN_6_port, PRGA_IN_5_port, PRGA_IN_4_port,
      PRGA_IN_3_port, PRGA_IN_2_port, PRGA_IN_1_port, PRGA_IN_0_port );
   PRGA_OPCODE <= ( PRGA_OPCODE_1_port, PRGA_OPCODE_0_port );
   
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n1, S => n89, Q => state_0_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n1, S => n90, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n1, S => n91, Q => state_1_port);
   B_READY_reg : DFFPOSX1 port map( D => n92, CLK => CLK, Q => B_READY_port);
   tempData_reg_7_inst : DFFPOSX1 port map( D => n68, CLK => CLK, Q => 
                           tempData_7_port);
   tempData_reg_6_inst : DFFPOSX1 port map( D => n69, CLK => CLK, Q => 
                           tempData_6_port);
   tempData_reg_5_inst : DFFPOSX1 port map( D => n70, CLK => CLK, Q => 
                           tempData_5_port);
   tempData_reg_4_inst : DFFPOSX1 port map( D => n71, CLK => CLK, Q => 
                           tempData_4_port);
   tempData_reg_3_inst : DFFPOSX1 port map( D => n72, CLK => CLK, Q => 
                           tempData_3_port);
   tempData_reg_2_inst : DFFPOSX1 port map( D => n73, CLK => CLK, Q => 
                           tempData_2_port);
   tempData_reg_1_inst : DFFPOSX1 port map( D => n74, CLK => CLK, Q => 
                           tempData_1_port);
   tempData_reg_0_inst : DFFPOSX1 port map( D => n75, CLK => CLK, Q => 
                           tempData_0_port);
   tempOpcode_reg_1_inst : DFFPOSX1 port map( D => n86, CLK => CLK, Q => 
                           tempOpcode_1_port);
   PRGA_OPCODE_reg_1_inst : DFFPOSX1 port map( D => n93, CLK => CLK, Q => 
                           PRGA_OPCODE_1_port);
   tempOpcode_reg_0_inst : DFFPOSX1 port map( D => n88, CLK => CLK, Q => 
                           tempOpcode_0_port);
   PRGA_OPCODE_reg_0_inst : DFFPOSX1 port map( D => n94, CLK => CLK, Q => 
                           PRGA_OPCODE_0_port);
   R_ENABLE_reg : DFFPOSX1 port map( D => n95, CLK => CLK, Q => R_ENABLE_port);
   PRGA_IN_reg_7_inst : DFFPOSX1 port map( D => n96, CLK => CLK, Q => 
                           PRGA_IN_7_port);
   PRGA_IN_reg_6_inst : DFFPOSX1 port map( D => n97, CLK => CLK, Q => 
                           PRGA_IN_6_port);
   PRGA_IN_reg_5_inst : DFFPOSX1 port map( D => n98, CLK => CLK, Q => 
                           PRGA_IN_5_port);
   PRGA_IN_reg_4_inst : DFFPOSX1 port map( D => n99, CLK => CLK, Q => 
                           PRGA_IN_4_port);
   PRGA_IN_reg_3_inst : DFFPOSX1 port map( D => n100, CLK => CLK, Q => 
                           PRGA_IN_3_port);
   PRGA_IN_reg_2_inst : DFFPOSX1 port map( D => n101, CLK => CLK, Q => 
                           PRGA_IN_2_port);
   PRGA_IN_reg_1_inst : DFFPOSX1 port map( D => n102, CLK => CLK, Q => 
                           PRGA_IN_1_port);
   PRGA_IN_reg_0_inst : DFFPOSX1 port map( D => n103, CLK => CLK, Q => 
                           PRGA_IN_0_port);
   n91 <= '1';
   n90 <= '1';
   n89 <= '1';
   U3 : INVX2 port map( A => n41, Y => n28);
   U4 : INVX2 port map( A => RST, Y => n1);
   U5 : OR2X2 port map( A => n39, B => RST, Y => n29);
   U6 : AND2X2 port map( A => n39, B => n1, Y => n44);
   U7 : OAI21X1 port map( A => n2, B => n3, C => n4, Y => nextState_2_port);
   U8 : MUX2X1 port map( B => n5, A => n6, S => state_0_port, Y => n4);
   U9 : NOR2X1 port map( A => state_2_port, B => n7, Y => n6);
   U10 : AND2X1 port map( A => state_2_port, B => n8, Y => n5);
   U11 : OAI21X1 port map( A => NEXT_BYTE, B => n9, C => state_1_port, Y => n8)
                           ;
   U12 : AND2X1 port map( A => n10, B => NEXT_BYTE, Y => n2);
   U13 : OAI21X1 port map( A => state_2_port, B => n11, C => n12, Y => 
                           nextState_1_port);
   U14 : OAI21X1 port map( A => n13, B => n14, C => n15, Y => n12);
   U15 : INVX1 port map( A => n3, Y => n14);
   U16 : OAI21X1 port map( A => state_2_port, B => n16, C => n17, Y => 
                           nextState_0_port);
   U17 : AOI22X1 port map( A => n18, B => n19, C => NEXT_BYTE, D => n20, Y => 
                           n17);
   U18 : OAI21X1 port map( A => n10, B => n3, C => n21, Y => n20);
   U19 : INVX1 port map( A => n13, Y => n21);
   U20 : NOR2X1 port map( A => n16, B => n9, Y => n13);
   U21 : NOR2X1 port map( A => n22, B => BYTE_COUNT(4), Y => n9);
   U22 : NAND3X1 port map( A => state_0_port, B => n7, C => state_2_port, Y => 
                           n3);
   U23 : AND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n10);
   U24 : OAI21X1 port map( A => n23, B => n15, C => n24, Y => n19);
   U25 : INVX1 port map( A => NEXT_BYTE, Y => n15);
   U26 : AOI21X1 port map( A => EOP, B => n22, C => BYTE_COUNT(4), Y => n23);
   U27 : NAND2X1 port map( A => n25, B => n26, Y => n22);
   U28 : NOR2X1 port map( A => BYTE_COUNT(3), B => BYTE_COUNT(2), Y => n26);
   U29 : NOR2X1 port map( A => BYTE_COUNT(1), B => BYTE_COUNT(0), Y => n25);
   U30 : NOR2X1 port map( A => state_1_port, B => state_0_port, Y => n18);
   U31 : INVX1 port map( A => n27, Y => n68);
   U32 : AOI22X1 port map( A => n28, B => DATA(7), C => n29, D => 
                           tempData_7_port, Y => n27);
   U33 : INVX1 port map( A => n30, Y => n69);
   U34 : AOI22X1 port map( A => n28, B => DATA(6), C => n29, D => 
                           tempData_6_port, Y => n30);
   U35 : INVX1 port map( A => n31, Y => n70);
   U36 : AOI22X1 port map( A => n28, B => DATA(5), C => n29, D => 
                           tempData_5_port, Y => n31);
   U37 : INVX1 port map( A => n32, Y => n71);
   U38 : AOI22X1 port map( A => n28, B => DATA(4), C => n29, D => 
                           tempData_4_port, Y => n32);
   U39 : INVX1 port map( A => n33, Y => n72);
   U40 : AOI22X1 port map( A => n28, B => DATA(3), C => n29, D => 
                           tempData_3_port, Y => n33);
   U41 : INVX1 port map( A => n34, Y => n73);
   U42 : AOI22X1 port map( A => n28, B => DATA(2), C => n29, D => 
                           tempData_2_port, Y => n34);
   U43 : INVX1 port map( A => n35, Y => n74);
   U44 : AOI22X1 port map( A => n28, B => DATA(1), C => n29, D => 
                           tempData_1_port, Y => n35);
   U45 : INVX1 port map( A => n36, Y => n75);
   U46 : AOI22X1 port map( A => n28, B => DATA(0), C => n29, D => 
                           tempData_0_port, Y => n36);
   U47 : INVX1 port map( A => n37, Y => n86);
   U48 : AOI22X1 port map( A => OPCODE(1), B => n28, C => n29, D => 
                           tempOpcode_1_port, Y => n37);
   U49 : INVX1 port map( A => n38, Y => n88);
   U50 : AOI22X1 port map( A => OPCODE(0), B => n28, C => n29, D => 
                           tempOpcode_0_port, Y => n38);
   U51 : OAI21X1 port map( A => n1, B => n40, C => n41, Y => n92);
   U52 : INVX1 port map( A => B_READY_port, Y => n40);
   U53 : OAI21X1 port map( A => n1, B => n42, C => n43, Y => n93);
   U54 : AOI22X1 port map( A => n28, B => OPCODE(1), C => n44, D => 
                           tempOpcode_1_port, Y => n43);
   U55 : INVX1 port map( A => PRGA_OPCODE_1_port, Y => n42);
   U56 : OAI21X1 port map( A => n1, B => n45, C => n46, Y => n94);
   U57 : AOI22X1 port map( A => n28, B => OPCODE(0), C => n44, D => 
                           tempOpcode_0_port, Y => n46);
   U58 : INVX1 port map( A => PRGA_OPCODE_0_port, Y => n45);
   U59 : MUX2X1 port map( B => n47, A => n48, S => RST, Y => n95);
   U60 : INVX1 port map( A => R_ENABLE_port, Y => n48);
   U61 : NAND3X1 port map( A => n7, B => n24, C => state_0_port, Y => n47);
   U62 : OAI21X1 port map( A => n1, B => n49, C => n50, Y => n96);
   U63 : AOI22X1 port map( A => DATA(7), B => n28, C => n44, D => 
                           tempData_7_port, Y => n50);
   U64 : INVX1 port map( A => PRGA_IN_7_port, Y => n49);
   U65 : OAI21X1 port map( A => n1, B => n51, C => n52, Y => n97);
   U66 : AOI22X1 port map( A => DATA(6), B => n28, C => n44, D => 
                           tempData_6_port, Y => n52);
   U67 : INVX1 port map( A => PRGA_IN_6_port, Y => n51);
   U68 : OAI21X1 port map( A => n1, B => n53, C => n54, Y => n98);
   U69 : AOI22X1 port map( A => DATA(5), B => n28, C => n44, D => 
                           tempData_5_port, Y => n54);
   U70 : INVX1 port map( A => PRGA_IN_5_port, Y => n53);
   U71 : OAI21X1 port map( A => n1, B => n55, C => n56, Y => n99);
   U72 : AOI22X1 port map( A => DATA(4), B => n28, C => n44, D => 
                           tempData_4_port, Y => n56);
   U73 : INVX1 port map( A => PRGA_IN_4_port, Y => n55);
   U74 : OAI21X1 port map( A => n1, B => n57, C => n58, Y => n100);
   U75 : AOI22X1 port map( A => DATA(3), B => n28, C => n44, D => 
                           tempData_3_port, Y => n58);
   U76 : INVX1 port map( A => PRGA_IN_3_port, Y => n57);
   U77 : OAI21X1 port map( A => n1, B => n59, C => n60, Y => n101);
   U78 : AOI22X1 port map( A => DATA(2), B => n28, C => n44, D => 
                           tempData_2_port, Y => n60);
   U79 : INVX1 port map( A => PRGA_IN_2_port, Y => n59);
   U80 : OAI21X1 port map( A => n1, B => n61, C => n62, Y => n102);
   U81 : AOI22X1 port map( A => DATA(1), B => n28, C => n44, D => 
                           tempData_1_port, Y => n62);
   U82 : INVX1 port map( A => PRGA_IN_1_port, Y => n61);
   U83 : OAI21X1 port map( A => n1, B => n63, C => n64, Y => n103);
   U84 : AOI22X1 port map( A => DATA(0), B => n28, C => n44, D => 
                           tempData_0_port, Y => n64);
   U85 : NAND2X1 port map( A => n11, B => state_2_port, Y => n39);
   U86 : INVX1 port map( A => n65, Y => n11);
   U87 : OAI21X1 port map( A => state_1_port, B => n66, C => n16, Y => n65);
   U88 : NAND2X1 port map( A => state_1_port, B => n66, Y => n16);
   U89 : NAND3X1 port map( A => n66, B => n7, C => n67, Y => n41);
   U90 : NOR2X1 port map( A => RST, B => n24, Y => n67);
   U91 : INVX1 port map( A => state_2_port, Y => n24);
   U92 : INVX1 port map( A => state_1_port, Y => n7);
   U93 : INVX1 port map( A => state_0_port, Y => n66);
   U94 : INVX1 port map( A => PRGA_IN_0_port, Y => n63);

end SYN_brbuffer;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_block_0 is

   port( CLK, RST, SERIAL_IN : in std_logic;  KEY_ERROR, PROG_ERROR : out 
         std_logic;  PLAINKEY : out std_logic_vector (63 downto 0);  RBUF_FULL,
         PARITY_ERROR : out std_logic);

end uart_rcv_block_0;

architecture SYN_struct1 of uart_rcv_block_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component uart_timer_0
      port( CLK, RST, TIMER_TRIG : in std_logic;  STOP_RCVING, SHIFT_STROBE : 
            out std_logic);
   end component;
   
   component keyreg_0
      port( CLK, RST, SBE, OE, RBUF_FULL : in std_logic;  RCV_DATA : in 
            std_logic_vector (7 downto 0);  PLAINKEY : out std_logic_vector (63
            downto 0);  KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR : out 
            std_logic);
   end component;
   
   component uart_sr_10bit_0
      port( CLK, RST, SHIFT_STROBE, SERIAL_IN : in std_logic;  LOAD_DATA : out 
            std_logic_vector (7 downto 0);  STOP_DATA : out std_logic_vector (1
            downto 0));
   end component;
   
   component uart_sb_check_0
      port( RST, CLK, SBC_CLR, SBC_EN : in std_logic;  STOP_DATA : in 
            std_logic_vector (1 downto 0);  SB_DETECT, SBE : out std_logic);
   end component;
   
   component uart_rcv_buf_full_0
      port( CLK, RST, CLR_RBUF, SET_RBUF_FULL : in std_logic;  RBUF_FULL : out 
            std_logic);
   end component;
   
   component uart_rcv_buf_0
      port( CLK, RST, LOAD_RBUF : in std_logic;  LOAD_DATA : in 
            std_logic_vector (7 downto 0);  RCV_DATA : out std_logic_vector (7 
            downto 0));
   end component;
   
   component uart_rcu_0
      port( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT : in std_logic;  
            RBUF_LOAD, TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR : 
            out std_logic);
   end component;
   
   component uart_error_0
      port( RST, CLK, RBUF_FULL, CHK_ERROR : in std_logic;  OE : out std_logic
            );
   end component;
   
   component uart_edge_detector_0
      port( CLK, RST, SERIAL_IN : in std_logic;  START_BIT : out std_logic);
   end component;
   
   signal RBUF_FULL_port, START_BIT, CHK_ERROR, OE, SB_DETECT, STOP_RCVING, 
      RBUF_LOAD, SBC_CLR, SBC_EN, SET_RBUF_FULL, TIMER_TRIG, LOAD_DATA_7_port, 
      LOAD_DATA_6_port, LOAD_DATA_5_port, LOAD_DATA_4_port, LOAD_DATA_3_port, 
      LOAD_DATA_2_port, LOAD_DATA_1_port, LOAD_DATA_0_port, RCV_DATA_7_port, 
      RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, RCV_DATA_3_port, 
      RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, CLR_RBUF, 
      STOP_DATA_1_port, STOP_DATA_0_port, SBE, SHIFT_STROBE, n1, n2 : std_logic
      ;

begin
   RBUF_FULL <= RBUF_FULL_port;
   
   U_0 : uart_edge_detector_0 port map( CLK => CLK, RST => n1, SERIAL_IN => 
                           SERIAL_IN, START_BIT => START_BIT);
   U_1 : uart_error_0 port map( RST => n1, CLK => CLK, RBUF_FULL => 
                           RBUF_FULL_port, CHK_ERROR => CHK_ERROR, OE => OE);
   U_2 : uart_rcu_0 port map( CLK => CLK, RST => n1, START_BIT => START_BIT, 
                           STOP_RCVING => STOP_RCVING, SB_DETECT => SB_DETECT, 
                           RBUF_LOAD => RBUF_LOAD, TIMER_TRIG => TIMER_TRIG, 
                           CHK_ERROR => CHK_ERROR, SET_RBUF_FULL => 
                           SET_RBUF_FULL, SBC_EN => SBC_EN, SBC_CLR => SBC_CLR)
                           ;
   U_3 : uart_rcv_buf_0 port map( CLK => CLK, RST => n1, LOAD_RBUF => RBUF_LOAD
                           , LOAD_DATA(7) => LOAD_DATA_7_port, LOAD_DATA(6) => 
                           LOAD_DATA_6_port, LOAD_DATA(5) => LOAD_DATA_5_port, 
                           LOAD_DATA(4) => LOAD_DATA_4_port, LOAD_DATA(3) => 
                           LOAD_DATA_3_port, LOAD_DATA(2) => LOAD_DATA_2_port, 
                           LOAD_DATA(1) => LOAD_DATA_1_port, LOAD_DATA(0) => 
                           LOAD_DATA_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port);
   U_4 : uart_rcv_buf_full_0 port map( CLK => CLK, RST => n1, CLR_RBUF => 
                           CLR_RBUF, SET_RBUF_FULL => SET_RBUF_FULL, RBUF_FULL 
                           => RBUF_FULL_port);
   U_5 : uart_sb_check_0 port map( RST => n1, CLK => CLK, SBC_CLR => SBC_CLR, 
                           SBC_EN => SBC_EN, STOP_DATA(1) => STOP_DATA_1_port, 
                           STOP_DATA(0) => STOP_DATA_0_port, SB_DETECT => 
                           SB_DETECT, SBE => SBE);
   U_6 : uart_sr_10bit_0 port map( CLK => CLK, RST => n1, SHIFT_STROBE => 
                           SHIFT_STROBE, SERIAL_IN => SERIAL_IN, LOAD_DATA(7) 
                           => LOAD_DATA_7_port, LOAD_DATA(6) => 
                           LOAD_DATA_6_port, LOAD_DATA(5) => LOAD_DATA_5_port, 
                           LOAD_DATA(4) => LOAD_DATA_4_port, LOAD_DATA(3) => 
                           LOAD_DATA_3_port, LOAD_DATA(2) => LOAD_DATA_2_port, 
                           LOAD_DATA(1) => LOAD_DATA_1_port, LOAD_DATA(0) => 
                           LOAD_DATA_0_port, STOP_DATA(1) => STOP_DATA_1_port, 
                           STOP_DATA(0) => STOP_DATA_0_port);
   U_8 : keyreg_0 port map( CLK => CLK, RST => n1, SBE => SBE, OE => OE, 
                           RBUF_FULL => RBUF_FULL_port, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           PLAINKEY(63) => PLAINKEY(63), PLAINKEY(62) => 
                           PLAINKEY(62), PLAINKEY(61) => PLAINKEY(61), 
                           PLAINKEY(60) => PLAINKEY(60), PLAINKEY(59) => 
                           PLAINKEY(59), PLAINKEY(58) => PLAINKEY(58), 
                           PLAINKEY(57) => PLAINKEY(57), PLAINKEY(56) => 
                           PLAINKEY(56), PLAINKEY(55) => PLAINKEY(55), 
                           PLAINKEY(54) => PLAINKEY(54), PLAINKEY(53) => 
                           PLAINKEY(53), PLAINKEY(52) => PLAINKEY(52), 
                           PLAINKEY(51) => PLAINKEY(51), PLAINKEY(50) => 
                           PLAINKEY(50), PLAINKEY(49) => PLAINKEY(49), 
                           PLAINKEY(48) => PLAINKEY(48), PLAINKEY(47) => 
                           PLAINKEY(47), PLAINKEY(46) => PLAINKEY(46), 
                           PLAINKEY(45) => PLAINKEY(45), PLAINKEY(44) => 
                           PLAINKEY(44), PLAINKEY(43) => PLAINKEY(43), 
                           PLAINKEY(42) => PLAINKEY(42), PLAINKEY(41) => 
                           PLAINKEY(41), PLAINKEY(40) => PLAINKEY(40), 
                           PLAINKEY(39) => PLAINKEY(39), PLAINKEY(38) => 
                           PLAINKEY(38), PLAINKEY(37) => PLAINKEY(37), 
                           PLAINKEY(36) => PLAINKEY(36), PLAINKEY(35) => 
                           PLAINKEY(35), PLAINKEY(34) => PLAINKEY(34), 
                           PLAINKEY(33) => PLAINKEY(33), PLAINKEY(32) => 
                           PLAINKEY(32), PLAINKEY(31) => PLAINKEY(31), 
                           PLAINKEY(30) => PLAINKEY(30), PLAINKEY(29) => 
                           PLAINKEY(29), PLAINKEY(28) => PLAINKEY(28), 
                           PLAINKEY(27) => PLAINKEY(27), PLAINKEY(26) => 
                           PLAINKEY(26), PLAINKEY(25) => PLAINKEY(25), 
                           PLAINKEY(24) => PLAINKEY(24), PLAINKEY(23) => 
                           PLAINKEY(23), PLAINKEY(22) => PLAINKEY(22), 
                           PLAINKEY(21) => PLAINKEY(21), PLAINKEY(20) => 
                           PLAINKEY(20), PLAINKEY(19) => PLAINKEY(19), 
                           PLAINKEY(18) => PLAINKEY(18), PLAINKEY(17) => 
                           PLAINKEY(17), PLAINKEY(16) => PLAINKEY(16), 
                           PLAINKEY(15) => PLAINKEY(15), PLAINKEY(14) => 
                           PLAINKEY(14), PLAINKEY(13) => PLAINKEY(13), 
                           PLAINKEY(12) => PLAINKEY(12), PLAINKEY(11) => 
                           PLAINKEY(11), PLAINKEY(10) => PLAINKEY(10), 
                           PLAINKEY(9) => PLAINKEY(9), PLAINKEY(8) => 
                           PLAINKEY(8), PLAINKEY(7) => PLAINKEY(7), PLAINKEY(6)
                           => PLAINKEY(6), PLAINKEY(5) => PLAINKEY(5), 
                           PLAINKEY(4) => PLAINKEY(4), PLAINKEY(3) => 
                           PLAINKEY(3), PLAINKEY(2) => PLAINKEY(2), PLAINKEY(1)
                           => PLAINKEY(1), PLAINKEY(0) => PLAINKEY(0), 
                           KEY_ERROR => KEY_ERROR, PROG_ERROR => PROG_ERROR, 
                           CLR_RBUFF => CLR_RBUF, PARITY_ERROR => PARITY_ERROR)
                           ;
   U_7 : uart_timer_0 port map( CLK => CLK, RST => n1, TIMER_TRIG => TIMER_TRIG
                           , STOP_RCVING => STOP_RCVING, SHIFT_STROBE => 
                           SHIFT_STROBE);
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct1;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0 is

   port( KEY : in std_logic_vector (63 downto 0);  CLK, RST, KEY_ERROR, 
         BYTE_READY : in std_logic;  BYTE : in std_logic_vector (7 downto 0);  
         OPCODE : in std_logic_vector (1 downto 0);  DATA_IN : in 
         std_logic_vector (7 downto 0);  PROCESSED_DATA : out std_logic_vector 
         (7 downto 0);  PDATA_READY, W_ENABLE, R_ENABLE : out std_logic;  ADDR,
         DATA : out std_logic_vector (7 downto 0));

end KSA_0;

architecture SYN_bksa of KSA_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUFX2
      port( A, EN : in std_logic;  Y : out std_logic);
   end component;
   
   component TBUFX1
      port( A, EN : in std_logic;  Y : out std_logic);
   end component;
   
   component KSA_0_DW01_inc_3
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_0_DW01_add_9
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_0_DW01_add_8
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_0_DW01_add_7
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_0_DW01_add_6
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_0_DW01_inc_1
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_0_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, PROCESSED_DATA_5_port, 
      PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, PROCESSED_DATA_2_port, 
      PROCESSED_DATA_1_port, PROCESSED_DATA_0_port, W_ENABLE_port, 
      R_ENABLE_port, ADDR_7_port, ADDR_6_port, ADDR_5_port, ADDR_4_port, 
      ADDR_3_port, ADDR_2_port, ADDR_1_port, ADDR_0_port, DATA_7_port, 
      DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, DATA_2_port, 
      DATA_1_port, DATA_0_port, state_4_port, state_3_port, state_2_port, 
      state_1_port, state_0_port, si_7_port, si_6_port, si_5_port, si_4_port, 
      si_3_port, si_2_port, si_1_port, si_0_port, sj_7_port, sj_6_port, 
      sj_5_port, sj_4_port, sj_3_port, sj_2_port, sj_1_port, sj_0_port, 
      currentProcessedData_7_port, currentProcessedData_6_port, 
      currentProcessedData_5_port, currentProcessedData_4_port, 
      currentProcessedData_3_port, currentProcessedData_2_port, 
      currentProcessedData_1_port, currentProcessedData_0_port, 
      nextState_4_port, nextState_3_port, nextState_2_port, nextState_1_port, 
      nextState_0_port, inti_7_port, inti_6_port, inti_5_port, inti_4_port, 
      inti_3_port, inti_2_port, inti_1_port, inti_0_port, intj_7_port, 
      intj_6_port, intj_5_port, intj_4_port, intj_3_port, intj_2_port, 
      intj_1_port, intj_0_port, keyi_2_port, keyi_1_port, keyi_0_port, 
      permuteComplete, temp_7_port, temp_6_port, temp_5_port, temp_4_port, 
      temp_3_port, temp_2_port, temp_1_port, temp_0_port, extratemp_7_port, 
      extratemp_6_port, extratemp_5_port, extratemp_4_port, extratemp_3_port, 
      extratemp_2_port, extratemp_1_port, extratemp_0_port, 
      nextProcessedData_7_port, nextProcessedData_6_port, 
      nextProcessedData_5_port, nextProcessedData_4_port, 
      nextProcessedData_3_port, nextProcessedData_2_port, 
      nextProcessedData_1_port, nextProcessedData_0_port, keyTable_0_7_port, 
      keyTable_0_6_port, keyTable_0_5_port, keyTable_0_4_port, 
      keyTable_0_3_port, keyTable_0_2_port, keyTable_0_1_port, 
      keyTable_0_0_port, keyTable_1_7_port, keyTable_1_6_port, 
      keyTable_1_5_port, keyTable_1_4_port, keyTable_1_3_port, 
      keyTable_1_2_port, keyTable_1_1_port, keyTable_1_0_port, 
      keyTable_2_7_port, keyTable_2_6_port, keyTable_2_5_port, 
      keyTable_2_4_port, keyTable_2_3_port, keyTable_2_2_port, 
      keyTable_2_1_port, keyTable_2_0_port, keyTable_3_7_port, 
      keyTable_3_6_port, keyTable_3_5_port, keyTable_3_4_port, 
      keyTable_3_3_port, keyTable_3_2_port, keyTable_3_1_port, 
      keyTable_3_0_port, keyTable_4_7_port, keyTable_4_6_port, 
      keyTable_4_5_port, keyTable_4_4_port, keyTable_4_3_port, 
      keyTable_4_2_port, keyTable_4_1_port, keyTable_4_0_port, 
      keyTable_5_7_port, keyTable_5_6_port, keyTable_5_5_port, 
      keyTable_5_4_port, keyTable_5_3_port, keyTable_5_2_port, 
      keyTable_5_1_port, keyTable_5_0_port, keyTable_6_7_port, 
      keyTable_6_6_port, keyTable_6_5_port, keyTable_6_4_port, 
      keyTable_6_3_port, keyTable_6_2_port, keyTable_6_1_port, 
      keyTable_6_0_port, keyTable_7_7_port, keyTable_7_6_port, 
      keyTable_7_5_port, keyTable_7_4_port, keyTable_7_3_port, 
      keyTable_7_2_port, keyTable_7_1_port, keyTable_7_0_port, delaydata_7_port
      , delaydata_6_port, delaydata_5_port, delaydata_4_port, delaydata_3_port,
      delaydata_2_port, delaydata_1_port, delaydata_0_port, 
      prefillCounter_7_port, prefillCounter_6_port, prefillCounter_5_port, 
      prefillCounter_4_port, prefillCounter_3_port, prefillCounter_2_port, 
      prefillCounter_1_port, prefillCounter_0_port, faddr_7_port, faddr_6_port,
      faddr_5_port, faddr_4_port, faddr_3_port, faddr_2_port, faddr_1_port, 
      faddr_0_port, nfaddr_7_port, nfaddr_6_port, nfaddr_5_port, nfaddr_4_port,
      nfaddr_3_port, nfaddr_2_port, nfaddr_1_port, nfaddr_0_port, fdata_7_port,
      fdata_6_port, fdata_5_port, fdata_4_port, fdata_3_port, fdata_2_port, 
      fdata_1_port, fdata_0_port, nfdata_7_port, nfdata_6_port, nfdata_5_port, 
      nfdata_4_port, nfdata_3_port, nfdata_2_port, nfdata_1_port, nfdata_0_port
      , fw_enable, fr_enable, N407, N408, N409, N410, N411, N412, N413, N414, 
      N424, N425, N426, N427, N428, N429, N430, N431, N472, N473, N474, N475, 
      N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, 
      N496, N497, N498, N499, N500, N501, N502, N503, N512, N513, N514, N515, 
      N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, 
      N456, N455, N454, N453, N452, N451, N450, N449, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n125, n127, n129, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n156, n157, n160, n161, n162, n164, 
      n166, n167, n169, n170, n171, n172, n175, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407_port, n408_port, n409_port
      , n410_port, n411_port, n412_port, n413_port, n414_port, n415, n416, n417
      , n418, n419, n420, n421, n422, n423, n424_port, n425_port, n426_port, 
      n427_port, n428_port, n429_port, n430_port, n431_port, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449_port, n450_port, n451_port, n452_port, n453_port, 
      n454_port, n455_port, n456_port, n457, n458, n459, n460, n461, n462, n463
      , n464, n465, n466, n467, n468, n469, n470, n471, n472_port, n473_port, 
      n474_port, n475_port, n476_port, n477_port, n478_port, n479_port, 
      n480_port, n481_port, n482_port, n483_port, n484_port, n485_port, 
      n486_port, n487_port, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496_port, n497_port, n498_port, n499_port, n500_port, n501_port, 
      n502_port, n503_port, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512_port, n513_port, n514_port, n515_port, n516_port, n517_port, 
      n518_port, n519_port, n520_port, n521_port, n522_port, n523_port, 
      n524_port, n525_port, n526_port, n527_port, n528, n529, n530, n531, n532,
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n692, n701, n746, n748, n750, n752, n754, n756, n758, n760, n765, n766, 
      n767, n768, n769, n771, n772, n773, n774, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n864, n865, n866, n867, n868, n869, n870, n871, 
      n883, n884, n885, n886, n887, n888, n889, n890, n898, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n_1024, n_1025, n_1026, n_1027 : std_logic;

begin
   PROCESSED_DATA <= ( PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, 
      PROCESSED_DATA_5_port, PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, 
      PROCESSED_DATA_2_port, PROCESSED_DATA_1_port, PROCESSED_DATA_0_port );
   W_ENABLE <= W_ENABLE_port;
   R_ENABLE <= R_ENABLE_port;
   ADDR <= ( ADDR_7_port, ADDR_6_port, ADDR_5_port, ADDR_4_port, ADDR_3_port, 
      ADDR_2_port, ADDR_1_port, ADDR_0_port );
   DATA <= ( DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, 
      DATA_2_port, DATA_1_port, DATA_0_port );
   
   n1336 <= '0';
   n1335 <= '0';
   prefillCounter_reg_0_inst : DFFPOSX1 port map( D => n1138, CLK => CLK, Q => 
                           prefillCounter_0_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n242, S => n1245, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n242, S => n1246, Q => state_2_port);
   state_reg_4_inst : DFFSR port map( D => nextState_4_port, CLK => CLK, R => 
                           n241, S => n1247, Q => state_4_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n241, S => n1248, Q => state_0_port);
   permuteComplete_reg : DFFPOSX1 port map( D => n1154, CLK => CLK, Q => 
                           permuteComplete);
   state_reg_3_inst : DFFSR port map( D => nextState_3_port, CLK => CLK, R => 
                           n241, S => n1249, Q => state_3_port);
   PDATA_READY_reg : DFFSR port map( D => n1134, CLK => CLK, R => n241, S => 
                           n1250, Q => PDATA_READY);
   extratemp_reg_7_inst : DFFPOSX1 port map( D => n1133, CLK => CLK, Q => 
                           extratemp_7_port);
   extratemp_reg_6_inst : DFFPOSX1 port map( D => n1132, CLK => CLK, Q => 
                           extratemp_6_port);
   extratemp_reg_5_inst : DFFPOSX1 port map( D => n1131, CLK => CLK, Q => 
                           extratemp_5_port);
   extratemp_reg_4_inst : DFFPOSX1 port map( D => n1130, CLK => CLK, Q => 
                           extratemp_4_port);
   extratemp_reg_3_inst : DFFPOSX1 port map( D => n1129, CLK => CLK, Q => 
                           extratemp_3_port);
   extratemp_reg_2_inst : DFFPOSX1 port map( D => n1128, CLK => CLK, Q => 
                           extratemp_2_port);
   extratemp_reg_1_inst : DFFPOSX1 port map( D => n1127, CLK => CLK, Q => 
                           extratemp_1_port);
   extratemp_reg_0_inst : DFFPOSX1 port map( D => n1126, CLK => CLK, Q => 
                           extratemp_0_port);
   keyTable_reg_7_0_inst : DFFPOSX1 port map( D => n1244, CLK => CLK, Q => 
                           keyTable_7_0_port);
   keyTable_reg_7_1_inst : DFFPOSX1 port map( D => n1243, CLK => CLK, Q => 
                           keyTable_7_1_port);
   keyTable_reg_7_2_inst : DFFPOSX1 port map( D => n1242, CLK => CLK, Q => 
                           keyTable_7_2_port);
   keyTable_reg_7_3_inst : DFFPOSX1 port map( D => n1241, CLK => CLK, Q => 
                           keyTable_7_3_port);
   keyTable_reg_7_4_inst : DFFPOSX1 port map( D => n1240, CLK => CLK, Q => 
                           keyTable_7_4_port);
   keyTable_reg_7_5_inst : DFFPOSX1 port map( D => n1239, CLK => CLK, Q => 
                           keyTable_7_5_port);
   keyTable_reg_7_6_inst : DFFPOSX1 port map( D => n1238, CLK => CLK, Q => 
                           keyTable_7_6_port);
   keyTable_reg_7_7_inst : DFFPOSX1 port map( D => n1237, CLK => CLK, Q => 
                           keyTable_7_7_port);
   keyTable_reg_6_0_inst : DFFPOSX1 port map( D => n1236, CLK => CLK, Q => 
                           keyTable_6_0_port);
   keyTable_reg_6_1_inst : DFFPOSX1 port map( D => n1235, CLK => CLK, Q => 
                           keyTable_6_1_port);
   keyTable_reg_6_2_inst : DFFPOSX1 port map( D => n1234, CLK => CLK, Q => 
                           keyTable_6_2_port);
   keyTable_reg_6_3_inst : DFFPOSX1 port map( D => n1233, CLK => CLK, Q => 
                           keyTable_6_3_port);
   keyTable_reg_6_4_inst : DFFPOSX1 port map( D => n1232, CLK => CLK, Q => 
                           keyTable_6_4_port);
   keyTable_reg_6_5_inst : DFFPOSX1 port map( D => n1231, CLK => CLK, Q => 
                           keyTable_6_5_port);
   keyTable_reg_6_6_inst : DFFPOSX1 port map( D => n1230, CLK => CLK, Q => 
                           keyTable_6_6_port);
   keyTable_reg_6_7_inst : DFFPOSX1 port map( D => n1229, CLK => CLK, Q => 
                           keyTable_6_7_port);
   keyTable_reg_5_0_inst : DFFPOSX1 port map( D => n1228, CLK => CLK, Q => 
                           keyTable_5_0_port);
   keyTable_reg_5_1_inst : DFFPOSX1 port map( D => n1227, CLK => CLK, Q => 
                           keyTable_5_1_port);
   keyTable_reg_5_2_inst : DFFPOSX1 port map( D => n1226, CLK => CLK, Q => 
                           keyTable_5_2_port);
   keyTable_reg_5_3_inst : DFFPOSX1 port map( D => n1225, CLK => CLK, Q => 
                           keyTable_5_3_port);
   keyTable_reg_5_4_inst : DFFPOSX1 port map( D => n1224, CLK => CLK, Q => 
                           keyTable_5_4_port);
   keyTable_reg_5_5_inst : DFFPOSX1 port map( D => n1223, CLK => CLK, Q => 
                           keyTable_5_5_port);
   keyTable_reg_5_6_inst : DFFPOSX1 port map( D => n1222, CLK => CLK, Q => 
                           keyTable_5_6_port);
   keyTable_reg_5_7_inst : DFFPOSX1 port map( D => n1221, CLK => CLK, Q => 
                           keyTable_5_7_port);
   keyTable_reg_4_0_inst : DFFPOSX1 port map( D => n1220, CLK => CLK, Q => 
                           keyTable_4_0_port);
   keyTable_reg_4_1_inst : DFFPOSX1 port map( D => n1219, CLK => CLK, Q => 
                           keyTable_4_1_port);
   keyTable_reg_4_2_inst : DFFPOSX1 port map( D => n1218, CLK => CLK, Q => 
                           keyTable_4_2_port);
   keyTable_reg_4_3_inst : DFFPOSX1 port map( D => n1217, CLK => CLK, Q => 
                           keyTable_4_3_port);
   keyTable_reg_4_4_inst : DFFPOSX1 port map( D => n1216, CLK => CLK, Q => 
                           keyTable_4_4_port);
   keyTable_reg_4_5_inst : DFFPOSX1 port map( D => n1215, CLK => CLK, Q => 
                           keyTable_4_5_port);
   keyTable_reg_4_6_inst : DFFPOSX1 port map( D => n1214, CLK => CLK, Q => 
                           keyTable_4_6_port);
   keyTable_reg_4_7_inst : DFFPOSX1 port map( D => n1213, CLK => CLK, Q => 
                           keyTable_4_7_port);
   keyTable_reg_3_0_inst : DFFPOSX1 port map( D => n1212, CLK => CLK, Q => 
                           keyTable_3_0_port);
   keyTable_reg_3_1_inst : DFFPOSX1 port map( D => n1211, CLK => CLK, Q => 
                           keyTable_3_1_port);
   keyTable_reg_3_2_inst : DFFPOSX1 port map( D => n1210, CLK => CLK, Q => 
                           keyTable_3_2_port);
   keyTable_reg_3_3_inst : DFFPOSX1 port map( D => n1209, CLK => CLK, Q => 
                           keyTable_3_3_port);
   keyTable_reg_3_4_inst : DFFPOSX1 port map( D => n1208, CLK => CLK, Q => 
                           keyTable_3_4_port);
   keyTable_reg_3_5_inst : DFFPOSX1 port map( D => n1207, CLK => CLK, Q => 
                           keyTable_3_5_port);
   keyTable_reg_3_6_inst : DFFPOSX1 port map( D => n1206, CLK => CLK, Q => 
                           keyTable_3_6_port);
   keyTable_reg_3_7_inst : DFFPOSX1 port map( D => n1205, CLK => CLK, Q => 
                           keyTable_3_7_port);
   keyTable_reg_2_0_inst : DFFPOSX1 port map( D => n1204, CLK => CLK, Q => 
                           keyTable_2_0_port);
   keyTable_reg_2_1_inst : DFFPOSX1 port map( D => n1203, CLK => CLK, Q => 
                           keyTable_2_1_port);
   keyTable_reg_2_2_inst : DFFPOSX1 port map( D => n1202, CLK => CLK, Q => 
                           keyTable_2_2_port);
   keyTable_reg_2_3_inst : DFFPOSX1 port map( D => n1201, CLK => CLK, Q => 
                           keyTable_2_3_port);
   keyTable_reg_2_4_inst : DFFPOSX1 port map( D => n1200, CLK => CLK, Q => 
                           keyTable_2_4_port);
   keyTable_reg_2_5_inst : DFFPOSX1 port map( D => n1199, CLK => CLK, Q => 
                           keyTable_2_5_port);
   keyTable_reg_2_6_inst : DFFPOSX1 port map( D => n1198, CLK => CLK, Q => 
                           keyTable_2_6_port);
   keyTable_reg_2_7_inst : DFFPOSX1 port map( D => n1197, CLK => CLK, Q => 
                           keyTable_2_7_port);
   keyTable_reg_1_0_inst : DFFPOSX1 port map( D => n1196, CLK => CLK, Q => 
                           keyTable_1_0_port);
   keyTable_reg_1_1_inst : DFFPOSX1 port map( D => n1195, CLK => CLK, Q => 
                           keyTable_1_1_port);
   keyTable_reg_1_2_inst : DFFPOSX1 port map( D => n1194, CLK => CLK, Q => 
                           keyTable_1_2_port);
   keyTable_reg_1_3_inst : DFFPOSX1 port map( D => n1193, CLK => CLK, Q => 
                           keyTable_1_3_port);
   keyTable_reg_1_4_inst : DFFPOSX1 port map( D => n1192, CLK => CLK, Q => 
                           keyTable_1_4_port);
   keyTable_reg_1_5_inst : DFFPOSX1 port map( D => n1191, CLK => CLK, Q => 
                           keyTable_1_5_port);
   keyTable_reg_1_6_inst : DFFPOSX1 port map( D => n1190, CLK => CLK, Q => 
                           keyTable_1_6_port);
   keyTable_reg_0_6_inst : DFFPOSX1 port map( D => n1189, CLK => CLK, Q => 
                           keyTable_0_6_port);
   keyTable_reg_0_5_inst : DFFPOSX1 port map( D => n1188, CLK => CLK, Q => 
                           keyTable_0_5_port);
   keyTable_reg_0_4_inst : DFFPOSX1 port map( D => n1187, CLK => CLK, Q => 
                           keyTable_0_4_port);
   keyTable_reg_0_3_inst : DFFPOSX1 port map( D => n1186, CLK => CLK, Q => 
                           keyTable_0_3_port);
   keyTable_reg_0_2_inst : DFFPOSX1 port map( D => n1185, CLK => CLK, Q => 
                           keyTable_0_2_port);
   keyTable_reg_0_1_inst : DFFPOSX1 port map( D => n1184, CLK => CLK, Q => 
                           keyTable_0_1_port);
   keyTable_reg_0_0_inst : DFFPOSX1 port map( D => n1183, CLK => CLK, Q => 
                           keyTable_0_0_port);
   keyTable_reg_1_7_inst : DFFPOSX1 port map( D => n1182, CLK => CLK, Q => 
                           keyTable_1_7_port);
   keyTable_reg_0_7_inst : DFFPOSX1 port map( D => n1181, CLK => CLK, Q => 
                           keyTable_0_7_port);
   prefillCounter_reg_7_inst : DFFPOSX1 port map( D => n1139, CLK => CLK, Q => 
                           prefillCounter_7_port);
   prefillCounter_reg_1_inst : DFFPOSX1 port map( D => n1140, CLK => CLK, Q => 
                           prefillCounter_1_port);
   prefillCounter_reg_2_inst : DFFPOSX1 port map( D => n1141, CLK => CLK, Q => 
                           prefillCounter_2_port);
   prefillCounter_reg_3_inst : DFFPOSX1 port map( D => n1142, CLK => CLK, Q => 
                           prefillCounter_3_port);
   prefillCounter_reg_4_inst : DFFPOSX1 port map( D => n1143, CLK => CLK, Q => 
                           prefillCounter_4_port);
   prefillCounter_reg_5_inst : DFFPOSX1 port map( D => n1144, CLK => CLK, Q => 
                           prefillCounter_5_port);
   prefillCounter_reg_6_inst : DFFPOSX1 port map( D => n1145, CLK => CLK, Q => 
                           prefillCounter_6_port);
   temp_reg_7_inst : DFFPOSX1 port map( D => n1180, CLK => CLK, Q => 
                           temp_7_port);
   temp_reg_0_inst : DFFPOSX1 port map( D => n1173, CLK => CLK, Q => 
                           temp_0_port);
   temp_reg_1_inst : DFFPOSX1 port map( D => n1174, CLK => CLK, Q => 
                           temp_1_port);
   temp_reg_2_inst : DFFPOSX1 port map( D => n1175, CLK => CLK, Q => 
                           temp_2_port);
   temp_reg_3_inst : DFFPOSX1 port map( D => n1176, CLK => CLK, Q => 
                           temp_3_port);
   temp_reg_4_inst : DFFPOSX1 port map( D => n1177, CLK => CLK, Q => 
                           temp_4_port);
   temp_reg_5_inst : DFFPOSX1 port map( D => n1178, CLK => CLK, Q => 
                           temp_5_port);
   temp_reg_6_inst : DFFPOSX1 port map( D => n1179, CLK => CLK, Q => 
                           temp_6_port);
   si_reg_0_inst : DFFSR port map( D => n1146, CLK => CLK, R => n241, S => 
                           n1251, Q => si_0_port);
   si_reg_1_inst : DFFSR port map( D => n1147, CLK => CLK, R => n240, S => 
                           n1252, Q => si_1_port);
   si_reg_6_inst : DFFSR port map( D => n1152, CLK => CLK, R => n240, S => 
                           n1253, Q => si_6_port);
   delaydata_reg_7_inst : DFFPOSX1 port map( D => n1110, CLK => CLK, Q => 
                           delaydata_7_port);
   delaydata_reg_0_inst : DFFPOSX1 port map( D => n1117, CLK => CLK, Q => 
                           delaydata_0_port);
   delaydata_reg_1_inst : DFFPOSX1 port map( D => n1116, CLK => CLK, Q => 
                           delaydata_1_port);
   delaydata_reg_2_inst : DFFPOSX1 port map( D => n1115, CLK => CLK, Q => 
                           delaydata_2_port);
   delaydata_reg_3_inst : DFFPOSX1 port map( D => n1114, CLK => CLK, Q => 
                           delaydata_3_port);
   delaydata_reg_4_inst : DFFPOSX1 port map( D => n1113, CLK => CLK, Q => 
                           delaydata_4_port);
   delaydata_reg_5_inst : DFFPOSX1 port map( D => n1112, CLK => CLK, Q => 
                           delaydata_5_port);
   delaydata_reg_6_inst : DFFPOSX1 port map( D => n1111, CLK => CLK, Q => 
                           delaydata_6_port);
   intj_reg_7_inst : DFFPOSX1 port map( D => n1169, CLK => CLK, Q => 
                           intj_7_port);
   intj_reg_0_inst : DFFPOSX1 port map( D => n1162, CLK => CLK, Q => 
                           intj_0_port);
   intj_reg_1_inst : DFFPOSX1 port map( D => n1163, CLK => CLK, Q => 
                           intj_1_port);
   intj_reg_2_inst : DFFPOSX1 port map( D => n1164, CLK => CLK, Q => 
                           intj_2_port);
   intj_reg_3_inst : DFFPOSX1 port map( D => n1165, CLK => CLK, Q => 
                           intj_3_port);
   intj_reg_4_inst : DFFPOSX1 port map( D => n1166, CLK => CLK, Q => 
                           intj_4_port);
   intj_reg_5_inst : DFFPOSX1 port map( D => n1167, CLK => CLK, Q => 
                           intj_5_port);
   intj_reg_6_inst : DFFPOSX1 port map( D => n1168, CLK => CLK, Q => 
                           intj_6_port);
   sj_reg_3_inst : DFFSR port map( D => n1158, CLK => CLK, R => n239, S => 
                           n1254, Q => sj_3_port);
   sj_reg_2_inst : DFFSR port map( D => n1159, CLK => CLK, R => n239, S => 
                           n1255, Q => sj_2_port);
   sj_reg_1_inst : DFFSR port map( D => n1160, CLK => CLK, R => n239, S => 
                           n1256, Q => sj_1_port);
   sj_reg_0_inst : DFFSR port map( D => n1161, CLK => CLK, R => n236, S => 
                           n1257, Q => sj_0_port);
   keyi_reg_2_inst : DFFPOSX1 port map( D => n1170, CLK => CLK, Q => 
                           keyi_2_port);
   keyi_reg_1_inst : DFFPOSX1 port map( D => n1171, CLK => CLK, Q => 
                           keyi_1_port);
   keyi_reg_0_inst : DFFPOSX1 port map( D => n1172, CLK => CLK, Q => 
                           keyi_0_port);
   inti_reg_7_inst : DFFPOSX1 port map( D => n1125, CLK => CLK, Q => 
                           inti_7_port);
   inti_reg_0_inst : DFFPOSX1 port map( D => n1118, CLK => CLK, Q => 
                           inti_0_port);
   inti_reg_1_inst : DFFPOSX1 port map( D => n1119, CLK => CLK, Q => 
                           inti_1_port);
   inti_reg_2_inst : DFFPOSX1 port map( D => n1120, CLK => CLK, Q => 
                           inti_2_port);
   inti_reg_3_inst : DFFPOSX1 port map( D => n1121, CLK => CLK, Q => 
                           inti_3_port);
   inti_reg_4_inst : DFFPOSX1 port map( D => n1122, CLK => CLK, Q => 
                           inti_4_port);
   inti_reg_5_inst : DFFPOSX1 port map( D => n1123, CLK => CLK, Q => 
                           inti_5_port);
   inti_reg_6_inst : DFFPOSX1 port map( D => n1124, CLK => CLK, Q => 
                           inti_6_port);
   PROCESSED_DATA_reg_0_inst : DFFPOSX1 port map( D => n1258, CLK => CLK, Q => 
                           PROCESSED_DATA_0_port);
   PROCESSED_DATA_reg_1_inst : DFFPOSX1 port map( D => n1259, CLK => CLK, Q => 
                           PROCESSED_DATA_1_port);
   PROCESSED_DATA_reg_2_inst : DFFPOSX1 port map( D => n1260, CLK => CLK, Q => 
                           PROCESSED_DATA_2_port);
   PROCESSED_DATA_reg_3_inst : DFFPOSX1 port map( D => n1261, CLK => CLK, Q => 
                           PROCESSED_DATA_3_port);
   PROCESSED_DATA_reg_4_inst : DFFPOSX1 port map( D => n1262, CLK => CLK, Q => 
                           PROCESSED_DATA_4_port);
   PROCESSED_DATA_reg_5_inst : DFFPOSX1 port map( D => n1263, CLK => CLK, Q => 
                           PROCESSED_DATA_5_port);
   PROCESSED_DATA_reg_6_inst : DFFPOSX1 port map( D => n1264, CLK => CLK, Q => 
                           PROCESSED_DATA_6_port);
   PROCESSED_DATA_reg_7_inst : DFFPOSX1 port map( D => n1265, CLK => CLK, Q => 
                           PROCESSED_DATA_7_port);
   faddr_reg_7_inst : DFFPOSX1 port map( D => n1266, CLK => CLK, Q => 
                           faddr_7_port);
   ADDR_reg_7_inst : DFFPOSX1 port map( D => n1267, CLK => CLK, Q => 
                           ADDR_7_port);
   faddr_reg_6_inst : DFFPOSX1 port map( D => n1268, CLK => CLK, Q => 
                           faddr_6_port);
   ADDR_reg_6_inst : DFFPOSX1 port map( D => n1269, CLK => CLK, Q => 
                           ADDR_6_port);
   faddr_reg_5_inst : DFFPOSX1 port map( D => n1270, CLK => CLK, Q => 
                           faddr_5_port);
   ADDR_reg_5_inst : DFFPOSX1 port map( D => n1271, CLK => CLK, Q => 
                           ADDR_5_port);
   faddr_reg_4_inst : DFFPOSX1 port map( D => n1272, CLK => CLK, Q => 
                           faddr_4_port);
   ADDR_reg_4_inst : DFFPOSX1 port map( D => n1273, CLK => CLK, Q => 
                           ADDR_4_port);
   faddr_reg_3_inst : DFFPOSX1 port map( D => n1274, CLK => CLK, Q => 
                           faddr_3_port);
   ADDR_reg_3_inst : DFFPOSX1 port map( D => n1275, CLK => CLK, Q => 
                           ADDR_3_port);
   faddr_reg_2_inst : DFFPOSX1 port map( D => n1276, CLK => CLK, Q => 
                           faddr_2_port);
   ADDR_reg_2_inst : DFFPOSX1 port map( D => n1277, CLK => CLK, Q => 
                           ADDR_2_port);
   faddr_reg_1_inst : DFFPOSX1 port map( D => n1278, CLK => CLK, Q => 
                           faddr_1_port);
   ADDR_reg_1_inst : DFFPOSX1 port map( D => n1279, CLK => CLK, Q => 
                           ADDR_1_port);
   faddr_reg_0_inst : DFFPOSX1 port map( D => n1280, CLK => CLK, Q => 
                           faddr_0_port);
   ADDR_reg_0_inst : DFFPOSX1 port map( D => n1281, CLK => CLK, Q => 
                           ADDR_0_port);
   fdata_reg_7_inst : DFFPOSX1 port map( D => n1282, CLK => CLK, Q => 
                           fdata_7_port);
   fdata_reg_6_inst : DFFPOSX1 port map( D => n1283, CLK => CLK, Q => 
                           fdata_6_port);
   fdata_reg_5_inst : DFFPOSX1 port map( D => n1284, CLK => CLK, Q => 
                           fdata_5_port);
   fdata_reg_4_inst : DFFPOSX1 port map( D => n1285, CLK => CLK, Q => 
                           fdata_4_port);
   fdata_reg_3_inst : DFFPOSX1 port map( D => n1286, CLK => CLK, Q => 
                           fdata_3_port);
   fdata_reg_2_inst : DFFPOSX1 port map( D => n1287, CLK => CLK, Q => 
                           fdata_2_port);
   fdata_reg_1_inst : DFFPOSX1 port map( D => n1288, CLK => CLK, Q => 
                           fdata_1_port);
   fdata_reg_0_inst : DFFPOSX1 port map( D => n1289, CLK => CLK, Q => 
                           fdata_0_port);
   fw_enable_reg : DFFPOSX1 port map( D => n1290, CLK => CLK, Q => fw_enable);
   fr_enable_reg : DFFPOSX1 port map( D => n1291, CLK => CLK, Q => fr_enable);
   W_ENABLE_reg : DFFPOSX1 port map( D => n1292, CLK => CLK, Q => W_ENABLE_port
                           );
   R_ENABLE_reg : DFFPOSX1 port map( D => n1293, CLK => CLK, Q => R_ENABLE_port
                           );
   DATA_reg_7_inst : DFFPOSX1 port map( D => n1294, CLK => CLK, Q => 
                           DATA_7_port);
   DATA_reg_6_inst : DFFPOSX1 port map( D => n1295, CLK => CLK, Q => 
                           DATA_6_port);
   DATA_reg_5_inst : DFFPOSX1 port map( D => n1296, CLK => CLK, Q => 
                           DATA_5_port);
   DATA_reg_4_inst : DFFPOSX1 port map( D => n1297, CLK => CLK, Q => 
                           DATA_4_port);
   DATA_reg_3_inst : DFFPOSX1 port map( D => n1298, CLK => CLK, Q => 
                           DATA_3_port);
   DATA_reg_2_inst : DFFPOSX1 port map( D => n1299, CLK => CLK, Q => 
                           DATA_2_port);
   DATA_reg_1_inst : DFFPOSX1 port map( D => n1300, CLK => CLK, Q => 
                           DATA_1_port);
   DATA_reg_0_inst : DFFPOSX1 port map( D => n1301, CLK => CLK, Q => 
                           DATA_0_port);
   U110 : NOR2X1 port map( A => KEY_ERROR, B => n1332, Y => n1333);
   U111 : OAI21X1 port map( A => n1106, B => n1331, C => n1105, Y => n1334);
   U123 : NOR2X1 port map( A => n1328, B => n1106, Y => n1330);
   U126 : NAND3X1 port map( A => n1327, B => n1100, C => n1326, Y => 
                           nextState_1_port);
   U130 : NOR2X1 port map( A => prefillCounter_2_port, B => 
                           prefillCounter_1_port, Y => n1324);
   U131 : NAND3X1 port map( A => n1323, B => n1135, C => n1322, Y => n1325);
   U132 : NOR2X1 port map( A => prefillCounter_4_port, B => 
                           prefillCounter_3_port, Y => n1322);
   U133 : NOR2X1 port map( A => prefillCounter_7_port, B => 
                           prefillCounter_6_port, Y => n1323);
   U143 : NAND3X1 port map( A => n1109, B => n1108, C => BYTE_READY, Y => n1329
                           );
   U156 : NAND2X1 port map( A => OPCODE(0), B => n1108, Y => n1331);
   U158 : NAND2X1 port map( A => BYTE_READY, B => n1320, Y => n1332);
   U159 : OAI21X1 port map( A => OPCODE(0), B => OPCODE(1), C => n1321, Y => 
                           n1320);
   U160 : NAND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n1321);
   U669 : NOR2X1 port map( A => n1103, B => n1104, Y => n1319);
   U673 : NOR2X1 port map( A => n1101, B => n1102, Y => n1318);
   n1257 <= '1';
   n1256 <= '1';
   n1255 <= '1';
   n1254 <= '1';
   n1253 <= '1';
   n1252 <= '1';
   n1251 <= '1';
   n1250 <= '1';
   n1249 <= '1';
   n1248 <= '1';
   n1247 <= '1';
   n1246 <= '1';
   n1245 <= '1';
   U142 : AND2X2 port map( A => n1331, B => n1321, Y => n1328);
   add_289 : KSA_0_DW01_inc_0 port map( A(7) => si_7_port, A(6) => si_6_port, 
                           A(5) => si_5_port, A(4) => si_4_port, A(3) => 
                           si_3_port, A(2) => si_2_port, A(1) => si_1_port, 
                           A(0) => si_0_port, SUM(7) => N431, SUM(6) => N430, 
                           SUM(5) => N429, SUM(4) => N428, SUM(3) => N427, 
                           SUM(2) => N426, SUM(1) => N425, SUM(0) => N424);
   add_263 : KSA_0_DW01_inc_1 port map( A(7) => prefillCounter_7_port, A(6) => 
                           prefillCounter_6_port, A(5) => prefillCounter_5_port
                           , A(4) => prefillCounter_4_port, A(3) => 
                           prefillCounter_3_port, A(2) => prefillCounter_2_port
                           , A(1) => prefillCounter_1_port, A(0) => 
                           prefillCounter_0_port, SUM(7) => N414, SUM(6) => 
                           N413, SUM(5) => N412, SUM(4) => N411, SUM(3) => N410
                           , SUM(2) => N409, SUM(1) => N408, SUM(0) => N407);
   add_377 : KSA_0_DW01_add_6 port map( A(7) => temp_7_port, A(6) => 
                           temp_6_port, A(5) => temp_5_port, A(4) => 
                           temp_4_port, A(3) => temp_3_port, A(2) => 
                           temp_2_port, A(1) => temp_1_port, A(0) => 
                           temp_0_port, B(7) => extratemp_7_port, B(6) => 
                           extratemp_6_port, B(5) => extratemp_5_port, B(4) => 
                           extratemp_4_port, B(3) => extratemp_3_port, B(2) => 
                           extratemp_2_port, B(1) => extratemp_1_port, B(0) => 
                           extratemp_0_port, CI => n1336, SUM(7) => N527, 
                           SUM(6) => N526, SUM(5) => N525, SUM(4) => N524, 
                           SUM(3) => N523, SUM(2) => N522, SUM(1) => N521, 
                           SUM(0) => N520, CO => n_1024);
   add_337 : KSA_0_DW01_add_7 port map( A(7) => intj_7_port, A(6) => 
                           intj_6_port, A(5) => intj_5_port, A(4) => 
                           intj_4_port, A(3) => intj_3_port, A(2) => 
                           intj_2_port, A(1) => intj_1_port, A(0) => 
                           intj_0_port, B(7) => DATA_IN(7), B(6) => DATA_IN(6),
                           B(5) => DATA_IN(5), B(4) => DATA_IN(4), B(3) => 
                           DATA_IN(3), B(2) => DATA_IN(2), B(1) => DATA_IN(1), 
                           B(0) => DATA_IN(0), CI => n1335, SUM(7) => N519, 
                           SUM(6) => N518, SUM(5) => N517, SUM(4) => N516, 
                           SUM(3) => N515, SUM(2) => N514, SUM(1) => N513, 
                           SUM(0) => N512, CO => n_1025);
   add_1_root_add_0_root_add_302_2 : KSA_0_DW01_add_8 port map( A(7) => 
                           DATA_IN(7), A(6) => DATA_IN(6), A(5) => DATA_IN(5), 
                           A(4) => DATA_IN(4), A(3) => DATA_IN(3), A(2) => 
                           DATA_IN(2), A(1) => DATA_IN(1), A(0) => DATA_IN(0), 
                           B(7) => sj_7_port, B(6) => sj_6_port, B(5) => 
                           sj_5_port, B(4) => sj_4_port, B(3) => sj_3_port, 
                           B(2) => sj_2_port, B(1) => sj_1_port, B(0) => n58, 
                           CI => n1136, SUM(7) => N456, SUM(6) => N455, SUM(5) 
                           => N454, SUM(4) => N453, SUM(3) => N452, SUM(2) => 
                           N451, SUM(1) => N450, SUM(0) => N449, CO => n_1026);
   add_0_root_add_0_root_add_302_2 : KSA_0_DW01_add_9 port map( A(7) => N472, 
                           A(6) => N473, A(5) => N474, A(4) => N475, A(3) => 
                           N476, A(2) => N477, A(1) => N478, A(0) => N479, B(7)
                           => N456, B(6) => N455, B(5) => N454, B(4) => N453, 
                           B(3) => N452, B(2) => N451, B(1) => N450, B(0) => 
                           N449, CI => n1137, SUM(7) => N487, SUM(6) => N486, 
                           SUM(5) => N485, SUM(4) => N484, SUM(3) => N483, 
                           SUM(2) => N482, SUM(1) => N481, SUM(0) => N480, CO 
                           => n_1027);
   r126 : KSA_0_DW01_inc_3 port map( A(7) => inti_7_port, A(6) => inti_6_port, 
                           A(5) => inti_5_port, A(4) => inti_4_port, A(3) => 
                           inti_3_port, A(2) => inti_2_port, A(1) => 
                           inti_1_port, A(0) => inti_0_port, SUM(7) => N503, 
                           SUM(6) => N502, SUM(5) => N501, SUM(4) => N500, 
                           SUM(3) => N499, SUM(2) => N498, SUM(1) => N497, 
                           SUM(0) => N496);
   nfdata_tri_0_inst : TBUFX1 port map( A => n1310, EN => n77, Y => 
                           nfdata_0_port);
   nfdata_tri_1_inst : TBUFX1 port map( A => n1311, EN => n77, Y => 
                           nfdata_1_port);
   nfdata_tri_2_inst : TBUFX1 port map( A => n1312, EN => n77, Y => 
                           nfdata_2_port);
   nfdata_tri_3_inst : TBUFX1 port map( A => n1313, EN => n77, Y => 
                           nfdata_3_port);
   nfdata_tri_4_inst : TBUFX1 port map( A => n1314, EN => n77, Y => 
                           nfdata_4_port);
   nfdata_tri_5_inst : TBUFX1 port map( A => n1315, EN => n77, Y => 
                           nfdata_5_port);
   nfdata_tri_6_inst : TBUFX1 port map( A => n1316, EN => n77, Y => 
                           nfdata_6_port);
   nfdata_tri_7_inst : TBUFX1 port map( A => n1317, EN => n77, Y => 
                           nfdata_7_port);
   nfaddr_tri_4_inst : TBUFX1 port map( A => n1306, EN => n1099, Y => 
                           nfaddr_4_port);
   nfaddr_tri_1_inst : TBUFX1 port map( A => n1303, EN => n1099, Y => 
                           nfaddr_1_port);
   nfaddr_tri_2_inst : TBUFX1 port map( A => n1304, EN => n1099, Y => 
                           nfaddr_2_port);
   nfaddr_tri_3_inst : TBUFX1 port map( A => n1305, EN => n1099, Y => 
                           nfaddr_3_port);
   nfaddr_tri_0_inst : TBUFX1 port map( A => n1302, EN => n1099, Y => 
                           nfaddr_0_port);
   nfaddr_tri_7_inst : TBUFX2 port map( A => n1309, EN => n1099, Y => 
                           nfaddr_7_port);
   nfaddr_tri_6_inst : TBUFX1 port map( A => n1308, EN => n1099, Y => 
                           nfaddr_6_port);
   nfaddr_tri_5_inst : TBUFX2 port map( A => n1307, EN => n1099, Y => 
                           nfaddr_5_port);
   si_reg_7_inst : DFFSR port map( D => n1153, CLK => CLK, R => n231, S => n30,
                           Q => si_7_port);
   si_reg_3_inst : DFFSR port map( D => n1149, CLK => CLK, R => n231, S => n29,
                           Q => si_3_port);
   si_reg_2_inst : DFFSR port map( D => n1148, CLK => CLK, R => n231, S => n28,
                           Q => si_2_port);
   si_reg_5_inst : DFFSR port map( D => n1151, CLK => CLK, R => n231, S => n27,
                           Q => si_5_port);
   si_reg_4_inst : DFFSR port map( D => n1150, CLK => CLK, R => n231, S => n26,
                           Q => si_4_port);
   sj_reg_4_inst : DFFSR port map( D => n1157, CLK => CLK, R => n231, S => n25,
                           Q => sj_4_port);
   currentProcessedData_reg_6_inst : DFFSR port map( D => 
                           nextProcessedData_6_port, CLK => CLK, R => n231, S 
                           => n24, Q => currentProcessedData_6_port);
   currentProcessedData_reg_4_inst : DFFSR port map( D => 
                           nextProcessedData_4_port, CLK => CLK, R => n231, S 
                           => n23, Q => currentProcessedData_4_port);
   currentProcessedData_reg_1_inst : DFFSR port map( D => 
                           nextProcessedData_1_port, CLK => CLK, R => n231, S 
                           => n22, Q => currentProcessedData_1_port);
   sj_reg_6_inst : DFFSR port map( D => n1155, CLK => CLK, R => n231, S => n21,
                           Q => sj_6_port);
   currentProcessedData_reg_7_inst : DFFSR port map( D => 
                           nextProcessedData_7_port, CLK => CLK, R => n231, S 
                           => n20, Q => currentProcessedData_7_port);
   currentProcessedData_reg_5_inst : DFFSR port map( D => 
                           nextProcessedData_5_port, CLK => CLK, R => n231, S 
                           => n19, Q => currentProcessedData_5_port);
   currentProcessedData_reg_3_inst : DFFSR port map( D => 
                           nextProcessedData_3_port, CLK => CLK, R => n231, S 
                           => n18, Q => currentProcessedData_3_port);
   currentProcessedData_reg_2_inst : DFFSR port map( D => 
                           nextProcessedData_2_port, CLK => CLK, R => n231, S 
                           => n17, Q => currentProcessedData_2_port);
   currentProcessedData_reg_0_inst : DFFSR port map( D => 
                           nextProcessedData_0_port, CLK => CLK, R => n231, S 
                           => n16, Q => currentProcessedData_0_port);
   sj_reg_5_inst : DFFSR port map( D => n1156, CLK => CLK, R => n231, S => n15,
                           Q => sj_5_port);
   sj_reg_7_inst : DFFSR port map( D => n1098, CLK => CLK, R => n231, S => n14,
                           Q => sj_7_port);
   U3 : AND2X1 port map( A => n1063, B => n236, Y => n3);
   U4 : AND2X2 port map( A => n175, B => n144, Y => n4);
   U7 : INVX2 port map( A => n701, Y => n73);
   U8 : AND2X2 port map( A => n303, B => n689, Y => n5);
   U9 : NAND2X1 port map( A => n185, B => n1088, Y => n6);
   U10 : AND2X2 port map( A => n153, B => n71, Y => n7);
   U11 : INVX1 port map( A => n701, Y => n452_port);
   U12 : AND2X2 port map( A => n1053, B => n1051, Y => n8);
   U13 : INVX2 port map( A => n225, Y => n342);
   U14 : INVX2 port map( A => n265, Y => n269);
   U15 : OR2X1 port map( A => n325, B => n324, Y => n9);
   U16 : OR2X2 port map( A => n361, B => n360, Y => n10);
   U17 : NAND2X1 port map( A => n33, B => n36, Y => n11);
   U18 : AND2X1 port map( A => n311, B => n312, Y => n12);
   U19 : AND2X2 port map( A => n65, B => n68, Y => n13);
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   n18 <= '1';
   n19 <= '1';
   n20 <= '1';
   n21 <= '1';
   n22 <= '1';
   n23 <= '1';
   n24 <= '1';
   n25 <= '1';
   n26 <= '1';
   n27 <= '1';
   n28 <= '1';
   n29 <= '1';
   n30 <= '1';
   U37 : NAND2X1 port map( A => n153, B => n71, Y => n31);
   U38 : INVX2 port map( A => n214, Y => n71);
   U39 : BUFX4 port map( A => n34, Y => n32);
   U40 : AND2X2 port map( A => n208, B => n144, Y => n33);
   U41 : NAND3X1 port map( A => keyi_1_port, B => keyi_0_port, C => n520_port, 
                           Y => n34);
   U42 : INVX1 port map( A => n169, Y => n35);
   U43 : BUFX4 port map( A => n216, Y => n169);
   U44 : INVX2 port map( A => n169, Y => n117);
   U45 : AND2X2 port map( A => n213, B => n299, Y => n36);
   U46 : INVX2 port map( A => state_2_port, Y => n299);
   U47 : NAND3X1 port map( A => n54, B => n267, C => n84, Y => n37);
   U48 : INVX1 port map( A => n171, Y => n38);
   U49 : NAND2X1 port map( A => n214, B => n299, Y => n39);
   U50 : XNOR2X1 port map( A => n49, B => n1069, Y => n254);
   U51 : NOR2X1 port map( A => n229, B => n1039, Y => n40);
   U52 : BUFX2 port map( A => n486_port, Y => n46);
   U53 : INVX1 port map( A => n215, Y => n1087);
   U54 : AND2X2 port map( A => n149, B => n252, Y => n208);
   U55 : INVX4 port map( A => keyi_1_port, Y => n519_port);
   U56 : INVX4 port map( A => keyi_0_port, Y => n521_port);
   U57 : INVX4 port map( A => keyi_2_port, Y => n520_port);
   U58 : BUFX4 port map( A => n36, Y => n41);
   U59 : AND2X2 port map( A => n229, B => n244, Y => n42);
   U60 : INVX4 port map( A => n83, Y => n171);
   U61 : INVX1 port map( A => n420, Y => n43);
   U62 : INVX2 port map( A => n43, Y => n44);
   U63 : BUFX4 port map( A => n486_port, Y => n45);
   U64 : BUFX2 port map( A => n175, Y => n47);
   U65 : INVX2 port map( A => n299, Y => n153);
   U66 : BUFX2 port map( A => n1063, Y => n48);
   U67 : BUFX4 port map( A => state_4_port, Y => n49);
   U68 : OAI21X1 port map( A => n52, B => n171, C => n300, Y => n50);
   U69 : INVX1 port map( A => n1073, Y => n226);
   U70 : INVX1 port map( A => n66, Y => n252);
   U71 : BUFX2 port map( A => n72, Y => n51);
   U72 : INVX2 port map( A => n36, Y => n52);
   U73 : NAND2X1 port map( A => n98, B => n1020, Y => n53);
   U74 : INVX2 port map( A => n97, Y => n98);
   U75 : NAND2X1 port map( A => n40, B => n41, Y => n54);
   U76 : INVX1 port map( A => n178, Y => n55);
   U77 : INVX1 port map( A => n55, Y => n56);
   U78 : INVX1 port map( A => n692, Y => n57);
   U79 : BUFX2 port map( A => state_1_port, Y => n149);
   U80 : BUFX4 port map( A => sj_0_port, Y => n58);
   U81 : INVX1 port map( A => n442, Y => n1274);
   U82 : INVX1 port map( A => n441, Y => n1275);
   U83 : AND2X2 port map( A => n639, B => n59, Y => n123);
   U84 : NOR2X1 port map( A => n180, B => n166, Y => n59);
   U85 : AND2X2 port map( A => n187, B => n679, Y => n60);
   U86 : BUFX4 port map( A => n1097, Y => n61);
   U87 : BUFX4 port map( A => n1097, Y => n62);
   U88 : AND2X2 port map( A => n210, B => n1057, Y => n147);
   U89 : INVX1 port map( A => n216, Y => n656);
   U90 : INVX2 port map( A => n1053, Y => n63);
   U91 : INVX1 port map( A => n60, Y => n64);
   U92 : INVX1 port map( A => n64, Y => n65);
   U93 : INVX2 port map( A => n211, Y => n66);
   U94 : INVX1 port map( A => n211, Y => n212);
   U95 : NAND2X1 port map( A => n154, B => n41, Y => n67);
   U96 : NAND2X1 port map( A => n154, B => n41, Y => n68);
   U97 : INVX1 port map( A => n310, Y => n99);
   U98 : BUFX2 port map( A => n196, Y => n69);
   U99 : NOR2X1 port map( A => n638, B => n180, Y => n70);
   U100 : INVX2 port map( A => n67, Y => n89);
   U101 : AND2X2 port map( A => n271, B => n270, Y => n187);
   U102 : INVX1 port map( A => n458, Y => n489);
   U103 : INVX2 port map( A => n39, Y => n72);
   U104 : INVX4 port map( A => n86, Y => n616);
   U105 : INVX2 port map( A => n211, Y => n74);
   U106 : INVX1 port map( A => n54, Y => n1053);
   U107 : AND2X2 port map( A => n271, B => n270, Y => n75);
   U108 : BUFX4 port map( A => n683, Y => n76);
   U109 : INVX1 port map( A => n683, Y => n228);
   U112 : INVX2 port map( A => n1061, Y => n77);
   U113 : INVX1 port map( A => n171, Y => n78);
   U114 : NOR2X1 port map( A => n364, B => si_3_port, Y => n79);
   U115 : INVX1 port map( A => n79, Y => n349);
   U116 : NAND2X1 port map( A => n109, B => n314, Y => n80);
   U117 : NOR2X1 port map( A => n80, B => n81, Y => n182);
   U118 : OR2X2 port map( A => n82, B => n497_port, Y => n81);
   U119 : INVX1 port map( A => n68, Y => n82);
   U120 : INVX2 port map( A => n214, Y => n1069);
   U121 : AND2X2 port map( A => n49, B => n196, Y => n83);
   U122 : AND2X2 port map( A => n210, B => n1057, Y => n84);
   U124 : INVX1 port map( A => n214, Y => n164);
   U125 : NOR2X1 port map( A => n215, B => n262, Y => n85);
   U127 : NOR2X1 port map( A => n359, B => n10, Y => n1305);
   U128 : MUX2X1 port map( B => faddr_6_port, A => nfaddr_6_port, S => n237, Y 
                           => n448);
   U129 : AND2X2 port map( A => n253, B => n617, Y => n86);
   U134 : BUFX2 port map( A => n221, Y => n87);
   U135 : INVX2 port map( A => n157, Y => n179);
   U136 : INVX1 port map( A => n118, Y => n88);
   U137 : NAND2X1 port map( A => n11, B => n3, Y => n690);
   U138 : MUX2X1 port map( B => ADDR_6_port, A => nfaddr_6_port, S => n238, Y 
                           => n447);
   U139 : NAND2X1 port map( A => n185, B => n1088, Y => n90);
   U140 : INVX2 port map( A => n104, Y => n1094);
   U141 : INVX1 port map( A => n228, Y => n91);
   U144 : AND2X2 port map( A => n79, B => n1103, Y => n92);
   U145 : INVX1 port map( A => n92, Y => n330);
   U146 : INVX1 port map( A => n445, Y => n1271);
   U147 : INVX8 port map( A => n76, Y => n93);
   U148 : INVX1 port map( A => n448, Y => n1268);
   U149 : INVX1 port map( A => n179, Y => n94);
   U150 : INVX1 port map( A => n447, Y => n1269);
   U151 : AND2X2 port map( A => n13, B => n221, Y => n223);
   U152 : INVX1 port map( A => n1020, Y => n95);
   U153 : INVX1 port map( A => n95, Y => n96);
   U154 : NAND2X1 port map( A => n150, B => n60, Y => n97);
   U155 : NAND2X1 port map( A => n98, B => n1020, Y => n773);
   U157 : INVX1 port map( A => n657, Y => n496_port);
   U161 : AND2X2 port map( A => n100, B => n99, Y => n311);
   U162 : NAND2X1 port map( A => n656, B => faddr_7_port, Y => n100);
   U163 : NAND2X1 port map( A => n109, B => n314, Y => n101);
   U164 : INVX1 port map( A => n151, Y => n102);
   U165 : NAND2X1 port map( A => n679, B => n75, Y => n103);
   U166 : AND2X2 port map( A => n746, B => n87, Y => n104);
   U167 : INVX1 port map( A => n75, Y => n105);
   U168 : INVX1 port map( A => n105, Y => n106);
   U169 : INVX1 port map( A => n5, Y => n225);
   U170 : NOR2X1 port map( A => n188, B => n108, Y => n107);
   U171 : NAND2X1 port map( A => n303, B => n305, Y => n108);
   U172 : INVX1 port map( A => n11, Y => n1061);
   U173 : BUFX2 port map( A => n185, Y => n109);
   U174 : INVX1 port map( A => si_0_port, Y => n1101);
   U175 : BUFX2 port map( A => n225, Y => n110);
   U176 : INVX2 port map( A => n1076, Y => n111);
   U177 : INVX1 port map( A => n182, Y => n112);
   U178 : INVX1 port map( A => n112, Y => n113);
   U179 : AND2X2 port map( A => n7, B => n175, Y => n114);
   U180 : AND2X1 port map( A => n7, B => n208, Y => n219);
   U181 : INVX1 port map( A => n228, Y => n115);
   U182 : INVX1 port map( A => n153, Y => n116);
   U183 : NOR2X1 port map( A => n118, B => n119, Y => n120);
   U184 : NOR2X1 port map( A => n120, B => n103, Y => n314);
   U185 : INVX1 port map( A => n33, Y => n118);
   U186 : INVX1 port map( A => n164, Y => n119);
   U187 : BUFX2 port map( A => n222, Y => n121);
   U188 : INVX1 port map( A => n1039, Y => n1040);
   U189 : INVX1 port map( A => n53, Y => n746);
   U190 : NOR2X1 port map( A => n326, B => n9, Y => n1308);
   U191 : AND2X2 port map( A => n491, B => n490, Y => n122);
   U192 : INVX1 port map( A => n122, Y => nextProcessedData_0_port);
   U193 : AND2X2 port map( A => n12, B => n313, Y => n1309);
   U194 : INVX1 port map( A => n123, Y => n1054);
   U195 : AND2X2 port map( A => n484_port, B => n483_port, Y => n125);
   U196 : INVX1 port map( A => n125, Y => nextProcessedData_1_port);
   U197 : AND2X2 port map( A => n480_port, B => n479_port, Y => n127);
   U198 : INVX1 port map( A => n127, Y => nextProcessedData_2_port);
   U199 : AND2X2 port map( A => n476_port, B => n475_port, Y => n129);
   U200 : INVX1 port map( A => n129, Y => nextProcessedData_3_port);
   U201 : AND2X2 port map( A => n472_port, B => n471, Y => n131);
   U202 : INVX1 port map( A => n131, Y => nextProcessedData_4_port);
   U203 : AND2X2 port map( A => n468, B => n467, Y => n132);
   U204 : INVX1 port map( A => n132, Y => nextProcessedData_5_port);
   U205 : AND2X2 port map( A => n464, B => n463, Y => n133);
   U206 : INVX1 port map( A => n133, Y => nextProcessedData_6_port);
   U207 : AND2X2 port map( A => n460, B => n459, Y => n134);
   U208 : INVX1 port map( A => n134, Y => nextProcessedData_7_port);
   U209 : AND2X2 port map( A => n1068, B => n206, Y => n135);
   U210 : INVX1 port map( A => n135, Y => n596);
   U211 : INVX1 port map( A => n92, Y => n136);
   U212 : INVX1 port map( A => n136, Y => n137);
   U213 : BUFX4 port map( A => n184, Y => n138);
   U214 : BUFX4 port map( A => n184, Y => n139);
   U215 : BUFX4 port map( A => n184, Y => n140);
   U216 : BUFX4 port map( A => n184, Y => n141);
   U217 : BUFX4 port map( A => n184, Y => n142);
   U218 : BUFX4 port map( A => n184, Y => n143);
   U219 : INVX2 port map( A => n49, Y => n144);
   U220 : INVX1 port map( A => n434, Y => n1282);
   U221 : INVX1 port map( A => n433, Y => n1283);
   U222 : INVX1 port map( A => n431_port, Y => n1285);
   U223 : INVX1 port map( A => n430_port, Y => n1286);
   U224 : INVX1 port map( A => n429_port, Y => n1287);
   U225 : INVX1 port map( A => n428_port, Y => n1288);
   U226 : INVX1 port map( A => n427_port, Y => n1289);
   U227 : INVX1 port map( A => n410_port, Y => n1294);
   U228 : INVX1 port map( A => n409_port, Y => n1295);
   U229 : INVX1 port map( A => n407_port, Y => n1297);
   U230 : INVX1 port map( A => n406, Y => n1298);
   U231 : INVX1 port map( A => n405, Y => n1299);
   U232 : INVX1 port map( A => n404, Y => n1300);
   U233 : INVX1 port map( A => n403, Y => n1301);
   U234 : INVX1 port map( A => n229, Y => n145);
   U235 : NOR2X1 port map( A => n229, B => n1039, Y => n189);
   U236 : BUFX2 port map( A => n329, Y => n146);
   U237 : INVX1 port map( A => n84, Y => n1046);
   U238 : AND2X2 port map( A => n329, B => n302, Y => n148);
   U239 : AND2X1 port map( A => n146, B => n302, Y => n199);
   U240 : BUFX2 port map( A => state_1_port, Y => n230);
   U241 : BUFX2 port map( A => n701, Y => n150);
   U242 : INVX1 port map( A => n450_port, Y => n1266);
   U243 : INVX1 port map( A => n449_port, Y => n1267);
   U244 : INVX1 port map( A => n160, Y => n151);
   U245 : NOR2X1 port map( A => n229, B => n152, Y => n160);
   U246 : NAND2X1 port map( A => n74, B => n243, Y => n152);
   U247 : INVX2 port map( A => n230, Y => n243);
   U248 : AND2X2 port map( A => n212, B => n243, Y => n196);
   U249 : BUFX2 port map( A => n190, Y => n154);
   U250 : AND2X2 port map( A => n259, B => n74, Y => n156);
   U251 : AND2X2 port map( A => n451_port, B => n458, Y => n157);
   U252 : INVX1 port map( A => n94, Y => n1134);
   U253 : INVX1 port map( A => n270, Y => n1042);
   U254 : INVX1 port map( A => n156, Y => n263);
   U255 : BUFX2 port map( A => n493, Y => n161);
   U256 : NAND3X1 port map( A => n54, B => n267, C => n84, Y => n162);
   U257 : NAND2X1 port map( A => n121, B => n1072, Y => n166);
   U258 : INVX1 port map( A => n101, Y => n1099);
   U259 : BUFX2 port map( A => n114, Y => n167);
   U260 : NAND2X1 port map( A => n85, B => n107, Y => n420);
   U261 : INVX4 port map( A => n188, Y => n222);
   U262 : AND2X2 port map( A => n153, B => n214, Y => n192);
   U263 : INVX2 port map( A => n590, Y => n170);
   U264 : NOR2X1 port map( A => n172, B => n162, Y => n216);
   U265 : NAND2X1 port map( A => n157, B => n67, Y => n172);
   U266 : AND2X2 port map( A => n149, B => n252, Y => n175);
   U267 : INVX2 port map( A => n253, Y => n177);
   U268 : INVX4 port map( A => n223, Y => n224);
   U269 : NOR2X1 port map( A => n1061, B => n655, Y => n660);
   U270 : AND2X1 port map( A => n96, B => n1019, Y => n181);
   U271 : OR2X1 port map( A => n568, B => n569, Y => n183);
   U272 : AND2X1 port map( A => keyi_2_port, B => keyi_1_port, Y => n200);
   U273 : INVX2 port map( A => n237, Y => n234);
   U274 : INVX2 port map( A => n238, Y => n233);
   U275 : INVX2 port map( A => n236, Y => n235);
   U276 : INVX2 port map( A => n654, Y => n1018);
   U277 : BUFX2 port map( A => n613, Y => n201);
   U278 : NOR2X1 port map( A => n179, B => n455_port, Y => n178);
   U279 : BUFX2 port map( A => n231, Y => n236);
   U280 : BUFX2 port map( A => n231, Y => n237);
   U281 : BUFX2 port map( A => n231, Y => n238);
   U282 : BUFX2 port map( A => n236, Y => n239);
   U283 : BUFX2 port map( A => n237, Y => n240);
   U284 : BUFX2 port map( A => n238, Y => n241);
   U285 : BUFX2 port map( A => n231, Y => n242);
   U286 : OR2X2 port map( A => n101, B => n232, Y => n180);
   U287 : AND2X2 port map( A => n221, B => n774, Y => n184);
   U288 : AND2X2 port map( A => n135, B => n1044, Y => n185);
   U289 : AND2X2 port map( A => n192, B => n156, Y => n188);
   U290 : AND2X2 port map( A => n197, B => n144, Y => n190);
   U291 : INVX2 port map( A => RST, Y => n231);
   U292 : AND2X2 port map( A => n200, B => n521_port, Y => n191);
   U293 : MUX2X1 port map( B => n1101, A => n521_port, S => n193, Y => n1172);
   U294 : NAND2X1 port map( A => n123, B => n68, Y => n193);
   U295 : MUX2X1 port map( B => n1102, A => n519_port, S => n194, Y => n1171);
   U296 : NAND2X1 port map( A => n123, B => n68, Y => n194);
   U297 : MUX2X1 port map( B => n650, A => n520_port, S => n195, Y => n1170);
   U298 : NAND2X1 port map( A => n123, B => n68, Y => n195);
   U299 : NOR2X1 port map( A => n149, B => n212, Y => n197);
   U300 : AND2X2 port map( A => n200, B => keyi_0_port, Y => n198);
   U301 : INVX1 port map( A => n638, Y => n639);
   U302 : INVX1 port map( A => n1057, Y => n1082);
   U303 : NAND2X1 port map( A => n272, B => n78, Y => n202);
   U304 : INVX1 port map( A => n689, Y => n294);
   U305 : BUFX2 port map( A => n1068, Y => n203);
   U306 : NAND2X1 port map( A => n205, B => n269, Y => n206);
   U307 : INVX1 port map( A => n31, Y => n205);
   U308 : NAND2X1 port map( A => n244, B => n229, Y => n207);
   U309 : BUFX2 port map( A => n149, Y => n209);
   U310 : INVX1 port map( A => n227, Y => n1074);
   U311 : INVX4 port map( A => n226, Y => n227);
   U312 : AND2X2 port map( A => n1072, B => n493, Y => n210);
   U313 : INVX1 port map( A => n210, Y => n1083);
   U314 : INVX2 port map( A => state_0_port, Y => n211);
   U315 : INVX2 port map( A => state_3_port, Y => n213);
   U316 : INVX4 port map( A => n213, Y => n214);
   U317 : AND2X2 port map( A => n219, B => n49, Y => n215);
   U318 : BUFX4 port map( A => state_4_port, Y => n229);
   U319 : AND2X1 port map( A => n1087, B => n150, Y => n255);
   U320 : INVX1 port map( A => n114, Y => n340);
   U321 : INVX1 port map( A => n1044, Y => n253);
   U322 : AND2X2 port map( A => n617, B => n111, Y => n217);
   U323 : AND2X2 port map( A => n617, B => n111, Y => n218);
   U324 : OR2X2 port map( A => n1080, B => n207, Y => n1063);
   U325 : INVX1 port map( A => n31, Y => n272);
   U326 : INVX1 port map( A => n1072, Y => n1076);
   U327 : INVX1 port map( A => n1088, Y => n590);
   U328 : INVX1 port map( A => n1080, Y => n1041);
   U329 : NAND2X1 port map( A => n181, B => n223, Y => n1021);
   U330 : NOR2X1 port map( A => n657, B => n183, Y => n574);
   U331 : INVX1 port map( A => n689, Y => n692);
   U332 : NOR2X1 port map( A => n638, B => n180, Y => n516_port);
   U333 : BUFX2 port map( A => n657, Y => n220);
   U334 : INVX2 port map( A => n242, Y => n232);
   U335 : AND2X2 port map( A => n178, B => n268, Y => n221);
   U336 : INVX1 port map( A => n87, Y => n423);
   U337 : INVX1 port map( A => n1063, Y => n295);
   U338 : INVX4 port map( A => n1021, Y => n1036);
   U339 : INVX8 port map( A => n76, Y => n684);
   U340 : INVX2 port map( A => si_1_port, Y => n1102);
   U341 : INVX2 port map( A => si_4_port, Y => n1103);
   U342 : INVX2 port map( A => si_5_port, Y => n1104);
   U343 : INVX2 port map( A => prefillCounter_5_port, Y => n1135);
   U344 : NAND3X1 port map( A => n197, B => n145, C => n192, Y => n1072);
   U345 : NOR2X1 port map( A => n230, B => n66, Y => n244);
   U346 : NAND2X1 port map( A => n42, B => n192, Y => n493);
   U347 : INVX2 port map( A => n1329, Y => n245);
   U348 : NAND2X1 port map( A => n1083, B => n245, Y => n250);
   U349 : NAND2X1 port map( A => n49, B => n196, Y => n264);
   U350 : NAND2X1 port map( A => n78, B => n245, Y => n247);
   U351 : NAND3X1 port map( A => n149, B => n74, C => n229, Y => n265);
   U352 : OAI21X1 port map( A => n1328, B => n1106, C => n269, Y => n246);
   U353 : NAND2X1 port map( A => n247, B => n246, Y => n248);
   U354 : NAND2X1 port map( A => n51, B => n248, Y => n249);
   U355 : NAND2X1 port map( A => n250, B => n249, Y => n251);
   U356 : AOI22X1 port map( A => n69, B => n41, C => n1105, D => n251, Y => 
                           n1327);
   U357 : NAND2X1 port map( A => n114, B => n145, Y => n1088);
   U358 : NAND2X1 port map( A => n149, B => n74, Y => n1039);
   U359 : NAND2X1 port map( A => n189, B => n72, Y => n270);
   U360 : INVX2 port map( A => permuteComplete, Y => n1050);
   U361 : NAND2X1 port map( A => n192, B => n33, Y => n1044);
   U362 : AOI21X1 port map( A => n1042, B => n1050, C => n253, Y => n256);
   U363 : NAND3X1 port map( A => n254, B => n175, C => n116, Y => n701);
   U364 : NAND3X1 port map( A => n1088, B => n256, C => n255, Y => n1065);
   U365 : INVX2 port map( A => n1065, Y => n1100);
   U366 : NOR2X1 port map( A => prefillCounter_0_port, B => n1325, Y => n257);
   U367 : NAND3X1 port map( A => n1324, B => n1061, C => n257, Y => n258);
   U368 : NAND3X1 port map( A => n72, B => n175, C => n49, Y => n458);
   U369 : NAND2X1 port map( A => n258, B => n458, Y => n261);
   U370 : NAND2X1 port map( A => n83, B => n7, Y => n679);
   U371 : NOR2X1 port map( A => n229, B => n149, Y => n259);
   U372 : NAND2X1 port map( A => n202, B => n263, Y => n260);
   U373 : NOR2X1 port map( A => n261, B => n260, Y => n1326);
   U374 : NAND2X1 port map( A => n42, B => n72, Y => n451_port);
   U375 : NAND2X1 port map( A => n42, B => n36, Y => n1068);
   U376 : NAND2X1 port map( A => n153, B => n1069, Y => n1080);
   U377 : NAND2X1 port map( A => n189, B => n7, Y => n300);
   U378 : OAI21X1 port map( A => n52, B => n171, C => n300, Y => n262);
   U379 : NOR2X1 port map( A => n215, B => n50, Y => n454_port);
   U380 : NAND2X1 port map( A => n190, B => n272, Y => n303);
   U381 : NAND2X1 port map( A => n40, B => n192, Y => n305);
   U382 : NOR2X1 port map( A => n90, B => n420, Y => n268);
   U383 : NAND2X1 port map( A => n40, B => n36, Y => n634);
   U384 : NAND2X1 port map( A => n102, B => n272, Y => n267);
   U385 : NAND2X1 port map( A => n265, B => n264, Y => n266);
   U386 : NAND2X1 port map( A => n72, B => n266, Y => n1057);
   U387 : NAND3X1 port map( A => n634, B => n267, C => n147, Y => n455_port);
   U388 : AOI22X1 port map( A => n160, B => n72, C => n269, D => n36, Y => n271
                           );
   U389 : NAND2X1 port map( A => n679, B => n187, Y => n569);
   U390 : NAND2X1 port map( A => n190, B => n72, Y => n689);
   U391 : NAND2X1 port map( A => n294, B => DATA_IN(7), Y => n274);
   U392 : NAND2X1 port map( A => n36, B => n156, Y => n654);
   U393 : NAND2X1 port map( A => prefillCounter_7_port, B => n1018, Y => n309);
   U394 : AOI22X1 port map( A => extratemp_7_port, B => n295, C => n73, D => 
                           temp_7_port, Y => n273);
   U395 : NAND3X1 port map( A => n274, B => n309, C => n273, Y => n275);
   U396 : AOI21X1 port map( A => fdata_7_port, B => n224, C => n275, Y => n1317
                           );
   U397 : NAND2X1 port map( A => n294, B => DATA_IN(6), Y => n277);
   U398 : NAND2X1 port map( A => prefillCounter_6_port, B => n1018, Y => n320);
   U399 : AOI22X1 port map( A => extratemp_6_port, B => n295, C => n73, D => 
                           temp_6_port, Y => n276);
   U400 : NAND3X1 port map( A => n277, B => n320, C => n276, Y => n278);
   U401 : AOI21X1 port map( A => fdata_6_port, B => n224, C => n278, Y => n1316
                           );
   U402 : NAND2X1 port map( A => n294, B => DATA_IN(5), Y => n280);
   U403 : NAND2X1 port map( A => n1018, B => prefillCounter_5_port, Y => n327);
   U404 : AOI22X1 port map( A => extratemp_5_port, B => n295, C => n73, D => 
                           temp_5_port, Y => n279);
   U405 : NAND3X1 port map( A => n280, B => n327, C => n279, Y => n281);
   U406 : AOI21X1 port map( A => n224, B => fdata_5_port, C => n281, Y => n1315
                           );
   U407 : NAND2X1 port map( A => n294, B => DATA_IN(4), Y => n283);
   U408 : NAND2X1 port map( A => prefillCounter_4_port, B => n1018, Y => n338);
   U409 : AOI22X1 port map( A => extratemp_4_port, B => n295, C => n73, D => 
                           temp_4_port, Y => n282);
   U410 : NAND3X1 port map( A => n283, B => n338, C => n282, Y => n284);
   U411 : AOI21X1 port map( A => fdata_4_port, B => n224, C => n284, Y => n1314
                           );
   U412 : NAND2X1 port map( A => n294, B => DATA_IN(3), Y => n286);
   U413 : NAND2X1 port map( A => prefillCounter_3_port, B => n1018, Y => n355);
   U414 : AOI22X1 port map( A => extratemp_3_port, B => n295, C => n73, D => 
                           temp_3_port, Y => n285);
   U415 : NAND3X1 port map( A => n286, B => n355, C => n285, Y => n287);
   U416 : AOI21X1 port map( A => fdata_3_port, B => n224, C => n287, Y => n1313
                           );
   U417 : NAND2X1 port map( A => n294, B => DATA_IN(2), Y => n289);
   U418 : NAND2X1 port map( A => prefillCounter_2_port, B => n1018, Y => n369);
   U419 : AOI22X1 port map( A => extratemp_2_port, B => n295, C => n73, D => 
                           temp_2_port, Y => n288);
   U420 : NAND3X1 port map( A => n289, B => n369, C => n288, Y => n290);
   U421 : AOI21X1 port map( A => fdata_2_port, B => n224, C => n290, Y => n1312
                           );
   U422 : NAND2X1 port map( A => n294, B => DATA_IN(1), Y => n292);
   U423 : NAND2X1 port map( A => prefillCounter_1_port, B => n1018, Y => n383);
   U424 : AOI22X1 port map( A => extratemp_1_port, B => n295, C => n73, D => 
                           temp_1_port, Y => n291);
   U425 : NAND3X1 port map( A => n292, B => n383, C => n291, Y => n293);
   U426 : AOI21X1 port map( A => fdata_1_port, B => n224, C => n293, Y => n1311
                           );
   U427 : NAND2X1 port map( A => n294, B => DATA_IN(0), Y => n297);
   U428 : NAND2X1 port map( A => prefillCounter_0_port, B => n1018, Y => n395);
   U429 : AOI22X1 port map( A => extratemp_0_port, B => n295, C => n73, D => 
                           temp_0_port, Y => n296);
   U430 : NAND3X1 port map( A => n297, B => n395, C => n296, Y => n298);
   U431 : AOI21X1 port map( A => n224, B => fdata_0_port, C => n298, Y => n1310
                           );
   U432 : NAND2X1 port map( A => n4, B => n116, Y => n411_port);
   U433 : NAND2X1 port map( A => n411_port, B => n300, Y => n390);
   U434 : OR2X2 port map( A => si_1_port, B => si_0_port, Y => n378);
   U435 : INVX2 port map( A => n378, Y => n301);
   U436 : INVX2 port map( A => si_2_port, Y => n650);
   U437 : NAND2X1 port map( A => n301, B => n650, Y => n364);
   U438 : INVX2 port map( A => si_3_port, Y => n648);
   U439 : NAND2X1 port map( A => n92, B => n1104, Y => n315);
   U440 : INVX2 port map( A => n315, Y => n329);
   U441 : INVX2 port map( A => si_6_port, Y => n302);
   U442 : XOR2X1 port map( A => n148, B => si_7_port, Y => n304);
   U443 : AOI22X1 port map( A => sj_7_port, B => n390, C => n304, D => n110, Y 
                           => n313);
   U444 : INVX2 port map( A => n222, Y => n497_port);
   U445 : NAND2X1 port map( A => n305, B => n1063, Y => n1073);
   U446 : AOI22X1 port map( A => N503, B => n497_port, C => intj_7_port, D => 
                           n227, Y => n312);
   U447 : NAND2X1 port map( A => temp_7_port, B => n167, Y => n308);
   U448 : OAI21X1 port map( A => n47, B => n38, C => n41, Y => n306);
   U449 : INVX2 port map( A => n306, Y => n397);
   U450 : NAND2X1 port map( A => n397, B => inti_7_port, Y => n307);
   U451 : NAND3X1 port map( A => n309, B => n308, C => n307, Y => n310);
   U452 : NAND2X1 port map( A => sj_6_port, B => n390, Y => n319);
   U453 : AND2X2 port map( A => si_6_port, B => n315, Y => n316);
   U454 : OAI21X1 port map( A => n199, B => n316, C => n110, Y => n318);
   U455 : AOI22X1 port map( A => intj_6_port, B => n227, C => N502, D => 
                           n497_port, Y => n317);
   U456 : NAND3X1 port map( A => n319, B => n318, C => n317, Y => n326);
   U457 : NAND2X1 port map( A => temp_6_port, B => n167, Y => n321);
   U458 : NAND2X1 port map( A => n321, B => n320, Y => n325);
   U459 : INVX2 port map( A => faddr_6_port, Y => n323);
   U460 : NAND2X1 port map( A => n397, B => inti_6_port, Y => n322);
   U461 : OAI21X1 port map( A => n169, B => n323, C => n322, Y => n324);
   U462 : INVX2 port map( A => temp_5_port, Y => n328);
   U463 : OAI21X1 port map( A => n340, B => n328, C => n327, Y => n335);
   U464 : AND2X2 port map( A => sj_5_port, B => n390, Y => n334);
   U465 : AOI21X1 port map( A => n330, B => si_5_port, C => n146, Y => n332);
   U466 : AOI22X1 port map( A => N501, B => n497_port, C => intj_5_port, D => 
                           n227, Y => n331);
   U467 : OAI21X1 port map( A => n332, B => n342, C => n331, Y => n333);
   U468 : NOR3X1 port map( A => n335, B => n334, C => n333, Y => n337);
   U469 : AOI22X1 port map( A => n117, B => faddr_5_port, C => n397, D => 
                           inti_5_port, Y => n336);
   U470 : AND2X2 port map( A => n337, B => n336, Y => n1307);
   U471 : INVX2 port map( A => temp_4_port, Y => n339);
   U472 : OAI21X1 port map( A => n340, B => n339, C => n338, Y => n346);
   U473 : AND2X2 port map( A => sj_4_port, B => n390, Y => n345);
   U474 : AOI21X1 port map( A => n349, B => si_4_port, C => n137, Y => n343);
   U475 : AOI22X1 port map( A => N500, B => n497_port, C => intj_4_port, D => 
                           n227, Y => n341);
   U476 : OAI21X1 port map( A => n343, B => n342, C => n341, Y => n344);
   U477 : NOR3X1 port map( A => n346, B => n345, C => n344, Y => n348);
   U478 : AOI22X1 port map( A => faddr_4_port, B => n117, C => n397, D => 
                           inti_4_port, Y => n347);
   U479 : AND2X2 port map( A => n348, B => n347, Y => n1306);
   U480 : NAND2X1 port map( A => sj_3_port, B => n390, Y => n354);
   U481 : NAND2X1 port map( A => si_3_port, B => n364, Y => n350);
   U482 : NAND2X1 port map( A => n350, B => n349, Y => n351);
   U483 : NAND2X1 port map( A => n351, B => n225, Y => n353);
   U484 : AOI22X1 port map( A => intj_3_port, B => n227, C => N499, D => 
                           n497_port, Y => n352);
   U485 : NAND3X1 port map( A => n354, B => n353, C => n352, Y => n361);
   U486 : NAND2X1 port map( A => temp_3_port, B => n167, Y => n356);
   U487 : NAND2X1 port map( A => n356, B => n355, Y => n360);
   U488 : INVX2 port map( A => faddr_3_port, Y => n358);
   U489 : NAND2X1 port map( A => n397, B => inti_3_port, Y => n357);
   U490 : OAI21X1 port map( A => n169, B => n358, C => n357, Y => n359);
   U491 : NAND2X1 port map( A => n397, B => inti_2_port, Y => n363);
   U492 : NAND2X1 port map( A => faddr_2_port, B => n35, Y => n362);
   U493 : NAND2X1 port map( A => n363, B => n362, Y => n375);
   U494 : NAND2X1 port map( A => si_2_port, B => n378, Y => n365);
   U495 : NAND2X1 port map( A => n365, B => n364, Y => n368);
   U496 : INVX2 port map( A => N498, Y => n507);
   U497 : NAND2X1 port map( A => intj_2_port, B => n227, Y => n366);
   U498 : OAI21X1 port map( A => n121, B => n507, C => n366, Y => n367);
   U499 : AOI21X1 port map( A => n368, B => n110, C => n367, Y => n373);
   U500 : NAND2X1 port map( A => sj_2_port, B => n390, Y => n372);
   U501 : INVX2 port map( A => n369, Y => n370);
   U502 : AOI21X1 port map( A => temp_2_port, B => n167, C => n370, Y => n371);
   U503 : NAND3X1 port map( A => n373, B => n372, C => n371, Y => n374);
   U504 : NOR2X1 port map( A => n375, B => n374, Y => n1304);
   U505 : NAND2X1 port map( A => n397, B => inti_1_port, Y => n377);
   U506 : NAND2X1 port map( A => faddr_1_port, B => n117, Y => n376);
   U507 : NAND2X1 port map( A => n377, B => n376, Y => n389);
   U508 : NAND2X1 port map( A => si_0_port, B => si_1_port, Y => n379);
   U509 : NAND2X1 port map( A => n379, B => n378, Y => n382);
   U510 : INVX2 port map( A => N497, Y => n509);
   U511 : NAND2X1 port map( A => intj_1_port, B => n227, Y => n380);
   U512 : OAI21X1 port map( A => n121, B => n509, C => n380, Y => n381);
   U513 : AOI21X1 port map( A => n382, B => n110, C => n381, Y => n387);
   U514 : NAND2X1 port map( A => sj_1_port, B => n390, Y => n386);
   U515 : INVX2 port map( A => n383, Y => n384);
   U516 : AOI21X1 port map( A => temp_1_port, B => n167, C => n384, Y => n385);
   U517 : NAND3X1 port map( A => n387, B => n386, C => n385, Y => n388);
   U518 : NOR2X1 port map( A => n389, B => n388, Y => n1303);
   U519 : NAND2X1 port map( A => n58, B => n390, Y => n394);
   U520 : NAND2X1 port map( A => n225, B => n1101, Y => n393);
   U521 : INVX2 port map( A => N496, Y => n511);
   U522 : NOR2X1 port map( A => n222, B => n511, Y => n391);
   U523 : AOI21X1 port map( A => intj_0_port, B => n227, C => n391, Y => n392);
   U524 : NAND3X1 port map( A => n394, B => n393, C => n392, Y => n402);
   U525 : NAND2X1 port map( A => temp_0_port, B => n167, Y => n396);
   U526 : NAND2X1 port map( A => n396, B => n395, Y => n401);
   U527 : INVX2 port map( A => faddr_0_port, Y => n399);
   U528 : NAND2X1 port map( A => n397, B => inti_0_port, Y => n398);
   U529 : OAI21X1 port map( A => n169, B => n399, C => n398, Y => n400);
   U530 : NOR3X1 port map( A => n402, B => n401, C => n400, Y => n1302);
   U531 : MUX2X1 port map( B => nfdata_0_port, A => DATA_0_port, S => n232, Y 
                           => n403);
   U532 : MUX2X1 port map( B => nfdata_1_port, A => DATA_1_port, S => n234, Y 
                           => n404);
   U533 : MUX2X1 port map( B => nfdata_2_port, A => DATA_2_port, S => n235, Y 
                           => n405);
   U534 : MUX2X1 port map( B => nfdata_3_port, A => DATA_3_port, S => n235, Y 
                           => n406);
   U535 : MUX2X1 port map( B => nfdata_4_port, A => DATA_4_port, S => n235, Y 
                           => n407_port);
   U536 : MUX2X1 port map( B => nfdata_5_port, A => DATA_5_port, S => n235, Y 
                           => n408_port);
   U537 : INVX2 port map( A => n408_port, Y => n1296);
   U538 : MUX2X1 port map( B => nfdata_6_port, A => DATA_6_port, S => n234, Y 
                           => n409_port);
   U539 : MUX2X1 port map( B => nfdata_7_port, A => DATA_7_port, S => n234, Y 
                           => n410_port);
   U540 : NOR2X1 port map( A => n1018, B => n103, Y => n413_port);
   U541 : AND2X2 port map( A => n411_port, B => n48, Y => n412_port);
   U542 : NAND3X1 port map( A => n413_port, B => n56, C => n412_port, Y => n419
                           );
   U543 : AOI21X1 port map( A => fr_enable, B => n419, C => n44, Y => n415);
   U544 : INVX2 port map( A => R_ENABLE_port, Y => n414_port);
   U545 : MUX2X1 port map( B => n415, A => n414_port, S => n234, Y => n1293);
   U546 : AND2X2 port map( A => n150, B => n654, Y => n416);
   U547 : NAND3X1 port map( A => n57, B => n48, C => n416, Y => n424_port);
   U548 : AOI21X1 port map( A => fw_enable, B => n423, C => n424_port, Y => 
                           n418);
   U549 : INVX2 port map( A => W_ENABLE_port, Y => n417);
   U550 : MUX2X1 port map( B => n418, A => n417, S => n234, Y => n1292);
   U551 : OAI21X1 port map( A => n235, B => n419, C => fr_enable, Y => n422);
   U552 : NAND2X1 port map( A => n44, B => n240, Y => n421);
   U553 : NAND2X1 port map( A => n422, B => n421, Y => n1291);
   U554 : OAI21X1 port map( A => n235, B => n423, C => fw_enable, Y => 
                           n426_port);
   U555 : NAND2X1 port map( A => n424_port, B => n238, Y => n425_port);
   U556 : NAND2X1 port map( A => n426_port, B => n425_port, Y => n1290);
   U557 : MUX2X1 port map( B => nfdata_0_port, A => fdata_0_port, S => n234, Y 
                           => n427_port);
   U558 : MUX2X1 port map( B => nfdata_1_port, A => fdata_1_port, S => n234, Y 
                           => n428_port);
   U559 : MUX2X1 port map( B => nfdata_2_port, A => fdata_2_port, S => n234, Y 
                           => n429_port);
   U560 : MUX2X1 port map( B => nfdata_3_port, A => fdata_3_port, S => n234, Y 
                           => n430_port);
   U561 : MUX2X1 port map( B => nfdata_4_port, A => fdata_4_port, S => n234, Y 
                           => n431_port);
   U562 : MUX2X1 port map( B => nfdata_5_port, A => fdata_5_port, S => n234, Y 
                           => n432);
   U563 : INVX2 port map( A => n432, Y => n1284);
   U564 : MUX2X1 port map( B => nfdata_6_port, A => fdata_6_port, S => n234, Y 
                           => n433);
   U565 : MUX2X1 port map( B => nfdata_7_port, A => fdata_7_port, S => n234, Y 
                           => n434);
   U566 : MUX2X1 port map( B => nfaddr_0_port, A => ADDR_0_port, S => n233, Y 
                           => n435);
   U567 : INVX2 port map( A => n435, Y => n1281);
   U568 : MUX2X1 port map( B => nfaddr_0_port, A => faddr_0_port, S => n233, Y 
                           => n436);
   U569 : INVX2 port map( A => n436, Y => n1280);
   U570 : MUX2X1 port map( B => nfaddr_1_port, A => ADDR_1_port, S => n233, Y 
                           => n437);
   U571 : INVX2 port map( A => n437, Y => n1279);
   U572 : MUX2X1 port map( B => nfaddr_1_port, A => faddr_1_port, S => n233, Y 
                           => n438);
   U573 : INVX2 port map( A => n438, Y => n1278);
   U574 : MUX2X1 port map( B => nfaddr_2_port, A => ADDR_2_port, S => n233, Y 
                           => n439);
   U575 : INVX2 port map( A => n439, Y => n1277);
   U576 : MUX2X1 port map( B => nfaddr_2_port, A => faddr_2_port, S => n233, Y 
                           => n440);
   U577 : INVX2 port map( A => n440, Y => n1276);
   U578 : MUX2X1 port map( B => nfaddr_3_port, A => ADDR_3_port, S => n233, Y 
                           => n441);
   U579 : MUX2X1 port map( B => nfaddr_3_port, A => faddr_3_port, S => n233, Y 
                           => n442);
   U580 : MUX2X1 port map( B => nfaddr_4_port, A => ADDR_4_port, S => n233, Y 
                           => n443);
   U581 : INVX2 port map( A => n443, Y => n1273);
   U582 : MUX2X1 port map( B => nfaddr_4_port, A => faddr_4_port, S => n233, Y 
                           => n444);
   U583 : INVX2 port map( A => n444, Y => n1272);
   U584 : MUX2X1 port map( B => nfaddr_5_port, A => ADDR_5_port, S => n233, Y 
                           => n445);
   U585 : MUX2X1 port map( B => nfaddr_5_port, A => faddr_5_port, S => n233, Y 
                           => n446);
   U586 : INVX2 port map( A => n446, Y => n1270);
   U587 : MUX2X1 port map( B => nfaddr_7_port, A => ADDR_7_port, S => n232, Y 
                           => n449_port);
   U588 : MUX2X1 port map( B => nfaddr_7_port, A => faddr_7_port, S => n233, Y 
                           => n450_port);
   U589 : INVX2 port map( A => n451_port, Y => n488);
   U590 : XOR2X1 port map( A => delaydata_7_port, B => temp_7_port, Y => n457);
   U591 : NOR2X1 port map( A => n452_port, B => n1073, Y => n453_port);
   U592 : NAND3X1 port map( A => n5, B => n454_port, C => n453_port, Y => n657)
                           ;
   U593 : NOR2X1 port map( A => n37, B => n220, Y => n456_port);
   U594 : NAND3X1 port map( A => n654, B => n182, C => n456_port, Y => 
                           n486_port);
   U595 : AOI22X1 port map( A => n488, B => n457, C => n45, D => 
                           currentProcessedData_7_port, Y => n460);
   U596 : NAND2X1 port map( A => BYTE(7), B => n489, Y => n459);
   U597 : INVX2 port map( A => PROCESSED_DATA_7_port, Y => n461);
   U598 : MUX2X1 port map( B => n134, A => n461, S => n232, Y => n1265);
   U599 : XOR2X1 port map( A => delaydata_6_port, B => temp_6_port, Y => n462);
   U600 : AOI22X1 port map( A => n488, B => n462, C => n46, D => 
                           currentProcessedData_6_port, Y => n464);
   U601 : NAND2X1 port map( A => BYTE(6), B => n489, Y => n463);
   U602 : INVX2 port map( A => PROCESSED_DATA_6_port, Y => n465);
   U603 : MUX2X1 port map( B => n133, A => n465, S => n232, Y => n1264);
   U604 : XOR2X1 port map( A => delaydata_5_port, B => temp_5_port, Y => n466);
   U605 : AOI22X1 port map( A => n488, B => n466, C => n45, D => 
                           currentProcessedData_5_port, Y => n468);
   U606 : NAND2X1 port map( A => BYTE(5), B => n489, Y => n467);
   U607 : INVX2 port map( A => PROCESSED_DATA_5_port, Y => n469);
   U608 : MUX2X1 port map( B => n132, A => n469, S => n232, Y => n1263);
   U609 : XOR2X1 port map( A => delaydata_4_port, B => temp_4_port, Y => n470);
   U610 : AOI22X1 port map( A => n488, B => n470, C => n46, D => 
                           currentProcessedData_4_port, Y => n472_port);
   U611 : NAND2X1 port map( A => BYTE(4), B => n489, Y => n471);
   U612 : INVX2 port map( A => PROCESSED_DATA_4_port, Y => n473_port);
   U613 : MUX2X1 port map( B => n131, A => n473_port, S => n232, Y => n1262);
   U614 : XOR2X1 port map( A => delaydata_3_port, B => temp_3_port, Y => 
                           n474_port);
   U615 : AOI22X1 port map( A => n488, B => n474_port, C => n45, D => 
                           currentProcessedData_3_port, Y => n476_port);
   U616 : NAND2X1 port map( A => BYTE(3), B => n489, Y => n475_port);
   U617 : INVX2 port map( A => PROCESSED_DATA_3_port, Y => n477_port);
   U618 : MUX2X1 port map( B => n129, A => n477_port, S => n232, Y => n1261);
   U619 : XOR2X1 port map( A => delaydata_2_port, B => temp_2_port, Y => 
                           n478_port);
   U620 : AOI22X1 port map( A => n488, B => n478_port, C => n45, D => 
                           currentProcessedData_2_port, Y => n480_port);
   U621 : NAND2X1 port map( A => BYTE(2), B => n489, Y => n479_port);
   U622 : INVX2 port map( A => PROCESSED_DATA_2_port, Y => n481_port);
   U623 : MUX2X1 port map( B => n127, A => n481_port, S => n232, Y => n1260);
   U624 : XOR2X1 port map( A => delaydata_1_port, B => temp_1_port, Y => 
                           n482_port);
   U625 : AOI22X1 port map( A => n488, B => n482_port, C => n46, D => 
                           currentProcessedData_1_port, Y => n484_port);
   U626 : NAND2X1 port map( A => BYTE(1), B => n489, Y => n483_port);
   U627 : INVX2 port map( A => PROCESSED_DATA_1_port, Y => n485_port);
   U628 : MUX2X1 port map( B => n125, A => n485_port, S => n232, Y => n1259);
   U629 : XOR2X1 port map( A => delaydata_0_port, B => temp_0_port, Y => 
                           n487_port);
   U630 : AOI22X1 port map( A => n488, B => n487_port, C => n45, D => 
                           currentProcessedData_0_port, Y => n491);
   U631 : NAND2X1 port map( A => BYTE(0), B => n489, Y => n490);
   U632 : INVX2 port map( A => PROCESSED_DATA_0_port, Y => n492);
   U633 : MUX2X1 port map( B => n122, A => n492, S => n232, Y => n1258);
   U634 : NAND2X1 port map( A => n102, B => n164, Y => n570);
   U635 : NAND2X1 port map( A => n161, B => n1057, Y => n1071);
   U636 : INVX2 port map( A => n1071, Y => n494);
   U637 : NAND2X1 port map( A => n494, B => n157, Y => n571);
   U638 : INVX2 port map( A => n571, Y => n495);
   U639 : NAND3X1 port map( A => n495, B => n570, C => n496_port, Y => n638);
   U640 : NAND2X1 port map( A => n497_port, B => n516_port, Y => n515_port);
   U641 : INVX2 port map( A => N502, Y => n499_port);
   U642 : NAND3X1 port map( A => n68, B => n63, C => n70, Y => n512_port);
   U643 : NAND2X1 port map( A => inti_6_port, B => n512_port, Y => n498_port);
   U644 : OAI21X1 port map( A => n515_port, B => n499_port, C => n498_port, Y 
                           => n1124);
   U645 : INVX2 port map( A => N501, Y => n501_port);
   U646 : NAND2X1 port map( A => inti_5_port, B => n512_port, Y => n500_port);
   U647 : OAI21X1 port map( A => n515_port, B => n501_port, C => n500_port, Y 
                           => n1123);
   U648 : INVX2 port map( A => N500, Y => n503_port);
   U649 : NAND2X1 port map( A => inti_4_port, B => n512_port, Y => n502_port);
   U650 : OAI21X1 port map( A => n515_port, B => n503_port, C => n502_port, Y 
                           => n1122);
   U651 : INVX2 port map( A => N499, Y => n505);
   U652 : NAND2X1 port map( A => inti_3_port, B => n512_port, Y => n504);
   U653 : OAI21X1 port map( A => n515_port, B => n505, C => n504, Y => n1121);
   U654 : NAND2X1 port map( A => inti_2_port, B => n512_port, Y => n506);
   U655 : OAI21X1 port map( A => n515_port, B => n507, C => n506, Y => n1120);
   U656 : NAND2X1 port map( A => inti_1_port, B => n512_port, Y => n508);
   U657 : OAI21X1 port map( A => n515_port, B => n509, C => n508, Y => n1119);
   U658 : NAND2X1 port map( A => inti_0_port, B => n512_port, Y => n510);
   U659 : OAI21X1 port map( A => n515_port, B => n511, C => n510, Y => n1118);
   U660 : INVX2 port map( A => N503, Y => n514_port);
   U661 : NAND2X1 port map( A => inti_7_port, B => n512_port, Y => n513_port);
   U662 : OAI21X1 port map( A => n515_port, B => n514_port, C => n513_port, Y 
                           => n1125);
   U663 : NAND3X1 port map( A => keyi_2_port, B => n519_port, C => n521_port, Y
                           => n517_port);
   U664 : INVX2 port map( A => n517_port, Y => n559);
   U665 : NAND3X1 port map( A => keyi_2_port, B => keyi_0_port, C => n519_port,
                           Y => n518_port);
   U666 : INVX2 port map( A => n518_port, Y => n558);
   U667 : AOI22X1 port map( A => keyTable_4_7_port, B => n559, C => 
                           keyTable_5_7_port, D => n558, Y => n527_port);
   U668 : AOI22X1 port map( A => keyTable_6_7_port, B => n191, C => 
                           keyTable_7_7_port, D => n198, Y => n526_port);
   U670 : INVX2 port map( A => keyTable_3_7_port, Y => n939);
   U671 : NAND3X1 port map( A => keyi_1_port, B => n520_port, C => n521_port, Y
                           => n560);
   U672 : INVX2 port map( A => keyTable_2_7_port, Y => n923);
   U674 : OAI22X1 port map( A => n32, B => n939, C => n560, D => n923, Y => 
                           n524_port);
   U675 : NAND3X1 port map( A => keyi_0_port, B => n520_port, C => n519_port, Y
                           => n562);
   U676 : INVX2 port map( A => keyTable_1_7_port, Y => n786);
   U677 : NOR2X1 port map( A => keyi_2_port, B => keyi_1_port, Y => n522_port);
   U678 : NAND2X1 port map( A => n522_port, B => n521_port, Y => n561);
   U679 : INVX2 port map( A => keyTable_0_7_port, Y => n784);
   U680 : OAI22X1 port map( A => n562, B => n786, C => n561, D => n784, Y => 
                           n523_port);
   U681 : NOR2X1 port map( A => n524_port, B => n523_port, Y => n525_port);
   U682 : NAND3X1 port map( A => n527_port, B => n526_port, C => n525_port, Y 
                           => N472);
   U683 : AOI22X1 port map( A => keyTable_4_6_port, B => n559, C => 
                           keyTable_5_6_port, D => n558, Y => n532);
   U684 : AOI22X1 port map( A => keyTable_6_6_port, B => n191, C => 
                           keyTable_7_6_port, D => n198, Y => n531);
   U685 : INVX2 port map( A => keyTable_3_6_port, Y => n941);
   U686 : INVX2 port map( A => keyTable_2_6_port, Y => n925);
   U687 : OAI22X1 port map( A => n32, B => n941, C => n560, D => n925, Y => 
                           n529);
   U688 : INVX2 port map( A => keyTable_1_6_port, Y => n885);
   U689 : INVX2 port map( A => keyTable_0_6_port, Y => n883);
   U690 : OAI22X1 port map( A => n562, B => n885, C => n561, D => n883, Y => 
                           n528);
   U691 : NOR2X1 port map( A => n529, B => n528, Y => n530);
   U692 : NAND3X1 port map( A => n532, B => n531, C => n530, Y => N473);
   U693 : AOI22X1 port map( A => keyTable_4_5_port, B => n559, C => 
                           keyTable_5_5_port, D => n558, Y => n537);
   U694 : AOI22X1 port map( A => keyTable_6_5_port, B => n191, C => 
                           keyTable_7_5_port, D => n198, Y => n536);
   U695 : INVX2 port map( A => keyTable_3_5_port, Y => n943);
   U696 : INVX2 port map( A => keyTable_2_5_port, Y => n927);
   U697 : OAI22X1 port map( A => n32, B => n943, C => n560, D => n927, Y => 
                           n534);
   U698 : INVX2 port map( A => keyTable_1_5_port, Y => n887);
   U699 : INVX2 port map( A => keyTable_0_5_port, Y => n870);
   U700 : OAI22X1 port map( A => n562, B => n887, C => n561, D => n870, Y => 
                           n533);
   U701 : NOR2X1 port map( A => n534, B => n533, Y => n535);
   U702 : NAND3X1 port map( A => n537, B => n536, C => n535, Y => N474);
   U703 : AOI22X1 port map( A => keyTable_4_4_port, B => n559, C => 
                           keyTable_5_4_port, D => n558, Y => n542);
   U704 : AOI22X1 port map( A => keyTable_6_4_port, B => n191, C => 
                           keyTable_7_4_port, D => n198, Y => n541);
   U705 : INVX2 port map( A => keyTable_3_4_port, Y => n945);
   U706 : INVX2 port map( A => keyTable_2_4_port, Y => n929);
   U707 : OAI22X1 port map( A => n32, B => n945, C => n560, D => n929, Y => 
                           n539);
   U708 : INVX2 port map( A => keyTable_1_4_port, Y => n889);
   U709 : INVX2 port map( A => keyTable_0_4_port, Y => n868);
   U710 : OAI22X1 port map( A => n562, B => n889, C => n561, D => n868, Y => 
                           n538);
   U711 : NOR2X1 port map( A => n539, B => n538, Y => n540);
   U712 : NAND3X1 port map( A => n542, B => n541, C => n540, Y => N475);
   U713 : AOI22X1 port map( A => keyTable_4_3_port, B => n559, C => 
                           keyTable_5_3_port, D => n558, Y => n547);
   U714 : AOI22X1 port map( A => keyTable_6_3_port, B => n191, C => 
                           keyTable_7_3_port, D => n198, Y => n546);
   U715 : INVX2 port map( A => keyTable_3_3_port, Y => n947);
   U716 : INVX2 port map( A => keyTable_2_3_port, Y => n931);
   U717 : OAI22X1 port map( A => n32, B => n947, C => n560, D => n931, Y => 
                           n544);
   U718 : INVX2 port map( A => keyTable_1_3_port, Y => n898);
   U719 : INVX2 port map( A => keyTable_0_3_port, Y => n866);
   U720 : OAI22X1 port map( A => n562, B => n898, C => n561, D => n866, Y => 
                           n543);
   U721 : NOR2X1 port map( A => n544, B => n543, Y => n545);
   U722 : NAND3X1 port map( A => n547, B => n546, C => n545, Y => N476);
   U723 : AOI22X1 port map( A => keyTable_4_2_port, B => n559, C => 
                           keyTable_5_2_port, D => n558, Y => n552);
   U724 : AOI22X1 port map( A => keyTable_6_2_port, B => n191, C => 
                           keyTable_7_2_port, D => n198, Y => n551);
   U725 : INVX2 port map( A => keyTable_3_2_port, Y => n949);
   U726 : INVX2 port map( A => keyTable_2_2_port, Y => n933);
   U727 : OAI22X1 port map( A => n32, B => n949, C => n560, D => n933, Y => 
                           n549);
   U728 : INVX2 port map( A => keyTable_1_2_port, Y => n917);
   U729 : INVX2 port map( A => keyTable_0_2_port, Y => n864);
   U730 : OAI22X1 port map( A => n562, B => n917, C => n561, D => n864, Y => 
                           n548);
   U731 : NOR2X1 port map( A => n549, B => n548, Y => n550);
   U732 : NAND3X1 port map( A => n552, B => n551, C => n550, Y => N477);
   U733 : AOI22X1 port map( A => keyTable_4_1_port, B => n559, C => 
                           keyTable_5_1_port, D => n558, Y => n557);
   U734 : AOI22X1 port map( A => keyTable_6_1_port, B => n191, C => 
                           keyTable_7_1_port, D => n198, Y => n556);
   U735 : INVX2 port map( A => keyTable_3_1_port, Y => n951);
   U736 : INVX2 port map( A => keyTable_2_1_port, Y => n935);
   U737 : OAI22X1 port map( A => n32, B => n951, C => n560, D => n935, Y => 
                           n554);
   U738 : INVX2 port map( A => keyTable_1_1_port, Y => n919);
   U739 : INVX2 port map( A => keyTable_0_1_port, Y => n790);
   U740 : OAI22X1 port map( A => n562, B => n919, C => n561, D => n790, Y => 
                           n553);
   U741 : NOR2X1 port map( A => n554, B => n553, Y => n555);
   U742 : NAND3X1 port map( A => n557, B => n556, C => n555, Y => N478);
   U743 : AOI22X1 port map( A => keyTable_4_0_port, B => n559, C => 
                           keyTable_5_0_port, D => n558, Y => n567);
   U744 : AOI22X1 port map( A => keyTable_6_0_port, B => n191, C => 
                           keyTable_7_0_port, D => n198, Y => n566);
   U745 : INVX2 port map( A => keyTable_3_0_port, Y => n953);
   U746 : INVX2 port map( A => keyTable_2_0_port, Y => n937);
   U747 : OAI22X1 port map( A => n32, B => n953, C => n560, D => n937, Y => 
                           n564);
   U748 : INVX2 port map( A => keyTable_1_0_port, Y => n921);
   U749 : INVX2 port map( A => keyTable_0_0_port, Y => n788);
   U750 : OAI22X1 port map( A => n562, B => n921, C => n561, D => n788, Y => 
                           n563);
   U751 : NOR2X1 port map( A => n564, B => n563, Y => n565);
   U752 : NAND3X1 port map( A => n567, B => n566, C => n565, Y => N479);
   U753 : NAND3X1 port map( A => n634, B => n11, C => n222, Y => n568);
   U754 : INVX2 port map( A => n570, Y => n572);
   U755 : NOR3X1 port map( A => n572, B => n89, C => n571, Y => n573);
   U756 : AND2X2 port map( A => n574, B => n573, Y => n597);
   U757 : NAND2X1 port map( A => n597, B => n109, Y => n593);
   U758 : INVX2 port map( A => n593, Y => n579);
   U759 : INVX2 port map( A => n58, Y => n576);
   U760 : NAND2X1 port map( A => N480, B => n590, Y => n575);
   U761 : OAI21X1 port map( A => n579, B => n576, C => n575, Y => n1161);
   U762 : INVX2 port map( A => sj_1_port, Y => n578);
   U763 : NAND2X1 port map( A => N481, B => n590, Y => n577);
   U764 : OAI21X1 port map( A => n579, B => n578, C => n577, Y => n1160);
   U765 : NAND2X1 port map( A => sj_2_port, B => n593, Y => n581);
   U766 : NAND2X1 port map( A => N482, B => n590, Y => n580);
   U767 : NAND2X1 port map( A => n581, B => n580, Y => n1159);
   U768 : NAND2X1 port map( A => sj_3_port, B => n593, Y => n583);
   U769 : NAND2X1 port map( A => N483, B => n590, Y => n582);
   U770 : NAND2X1 port map( A => n583, B => n582, Y => n1158);
   U771 : NAND2X1 port map( A => sj_4_port, B => n593, Y => n585);
   U772 : NAND2X1 port map( A => N484, B => n590, Y => n584);
   U773 : NAND2X1 port map( A => n585, B => n584, Y => n1157);
   U774 : NAND2X1 port map( A => sj_5_port, B => n593, Y => n587);
   U775 : NAND2X1 port map( A => N485, B => n590, Y => n586);
   U776 : NAND2X1 port map( A => n587, B => n586, Y => n1156);
   U777 : NAND2X1 port map( A => sj_6_port, B => n593, Y => n592);
   U778 : NAND2X1 port map( A => N486, B => n590, Y => n591);
   U779 : NAND2X1 port map( A => n592, B => n591, Y => n1155);
   U780 : NAND2X1 port map( A => sj_7_port, B => n593, Y => n595);
   U781 : INVX2 port map( A => N487, Y => n594);
   U782 : AOI22X1 port map( A => n595, B => n170, C => n595, D => n594, Y => 
                           n1098);
   U783 : NOR2X1 port map( A => n235, B => n596, Y => n598);
   U784 : NAND3X1 port map( A => n598, B => n1088, C => n597, Y => n613);
   U785 : INVX2 port map( A => n613, Y => n617);
   U786 : INVX2 port map( A => N518, Y => n600);
   U787 : NAND2X1 port map( A => intj_6_port, B => n201, Y => n599);
   U788 : OAI21X1 port map( A => n616, B => n600, C => n599, Y => n1168);
   U789 : INVX2 port map( A => N517, Y => n602);
   U790 : NAND2X1 port map( A => intj_5_port, B => n201, Y => n601);
   U791 : OAI21X1 port map( A => n616, B => n602, C => n601, Y => n1167);
   U792 : INVX2 port map( A => N516, Y => n604);
   U793 : NAND2X1 port map( A => intj_4_port, B => n201, Y => n603);
   U794 : OAI21X1 port map( A => n616, B => n604, C => n603, Y => n1166);
   U795 : INVX2 port map( A => N515, Y => n606);
   U796 : NAND2X1 port map( A => intj_3_port, B => n201, Y => n605);
   U797 : OAI21X1 port map( A => n616, B => n606, C => n605, Y => n1165);
   U798 : INVX2 port map( A => N514, Y => n608);
   U799 : NAND2X1 port map( A => intj_2_port, B => n201, Y => n607);
   U800 : OAI21X1 port map( A => n616, B => n608, C => n607, Y => n1164);
   U801 : INVX2 port map( A => N513, Y => n610);
   U802 : NAND2X1 port map( A => intj_1_port, B => n201, Y => n609);
   U803 : OAI21X1 port map( A => n616, B => n610, C => n609, Y => n1163);
   U804 : INVX2 port map( A => N512, Y => n612);
   U805 : NAND2X1 port map( A => intj_0_port, B => n201, Y => n611);
   U806 : OAI21X1 port map( A => n616, B => n612, C => n611, Y => n1162);
   U807 : INVX2 port map( A => N519, Y => n615);
   U808 : NAND2X1 port map( A => intj_7_port, B => n201, Y => n614);
   U809 : OAI21X1 port map( A => n616, B => n615, C => n614, Y => n1169);
   U810 : INVX2 port map( A => delaydata_6_port, Y => n619);
   U811 : INVX2 port map( A => BYTE(6), Y => n618);
   U812 : MUX2X1 port map( B => n619, A => n618, S => n218, Y => n1111);
   U813 : INVX2 port map( A => delaydata_5_port, Y => n621);
   U814 : INVX2 port map( A => BYTE(5), Y => n620);
   U815 : MUX2X1 port map( B => n621, A => n620, S => n217, Y => n1112);
   U816 : INVX2 port map( A => delaydata_4_port, Y => n623);
   U817 : INVX2 port map( A => BYTE(4), Y => n622);
   U818 : MUX2X1 port map( B => n623, A => n622, S => n218, Y => n1113);
   U819 : INVX2 port map( A => delaydata_3_port, Y => n625);
   U820 : INVX2 port map( A => BYTE(3), Y => n624);
   U821 : MUX2X1 port map( B => n625, A => n624, S => n217, Y => n1114);
   U822 : INVX2 port map( A => delaydata_2_port, Y => n627);
   U823 : INVX2 port map( A => BYTE(2), Y => n626);
   U824 : MUX2X1 port map( B => n627, A => n626, S => n218, Y => n1115);
   U825 : INVX2 port map( A => delaydata_1_port, Y => n629);
   U826 : INVX2 port map( A => BYTE(1), Y => n628);
   U827 : MUX2X1 port map( B => n629, A => n628, S => n217, Y => n1116);
   U828 : INVX2 port map( A => delaydata_0_port, Y => n631);
   U829 : INVX2 port map( A => BYTE(0), Y => n630);
   U830 : MUX2X1 port map( B => n631, A => n630, S => n218, Y => n1117);
   U831 : INVX2 port map( A => delaydata_7_port, Y => n633);
   U832 : INVX2 port map( A => BYTE(7), Y => n632);
   U833 : MUX2X1 port map( B => n633, A => n632, S => n217, Y => n1110);
   U834 : NAND3X1 port map( A => si_3_port, B => si_2_port, C => si_6_port, Y 
                           => n636);
   U835 : NAND2X1 port map( A => n1319, B => si_7_port, Y => n635);
   U836 : NOR2X1 port map( A => n636, B => n635, Y => n637);
   U837 : NAND2X1 port map( A => n637, B => n1318, Y => n1051);
   U838 : NAND2X1 port map( A => N431, B => n8, Y => n641);
   U839 : NAND2X1 port map( A => n113, B => n639, Y => n644);
   U840 : NAND2X1 port map( A => si_7_port, B => n644, Y => n640);
   U841 : NAND2X1 port map( A => n641, B => n640, Y => n1153);
   U842 : NAND2X1 port map( A => N430, B => n8, Y => n643);
   U843 : NAND2X1 port map( A => si_6_port, B => n644, Y => n642);
   U844 : NAND2X1 port map( A => n643, B => n642, Y => n1152);
   U845 : INVX2 port map( A => n644, Y => n653);
   U846 : NAND2X1 port map( A => N429, B => n8, Y => n645);
   U847 : OAI21X1 port map( A => n1104, B => n653, C => n645, Y => n1151);
   U848 : NAND2X1 port map( A => N428, B => n8, Y => n646);
   U849 : OAI21X1 port map( A => n1103, B => n653, C => n646, Y => n1150);
   U850 : NAND2X1 port map( A => N427, B => n8, Y => n647);
   U851 : OAI21X1 port map( A => n653, B => n648, C => n647, Y => n1149);
   U852 : NAND2X1 port map( A => N426, B => n8, Y => n649);
   U853 : OAI21X1 port map( A => n653, B => n650, C => n649, Y => n1148);
   U854 : NAND2X1 port map( A => N425, B => n8, Y => n651);
   U855 : OAI21X1 port map( A => n1102, B => n653, C => n651, Y => n1147);
   U856 : NAND2X1 port map( A => N424, B => n8, Y => n652);
   U857 : OAI21X1 port map( A => n1101, B => n653, C => n652, Y => n1146);
   U858 : NAND2X1 port map( A => n222, B => n654, Y => n655);
   U859 : NAND2X1 port map( A => n106, B => n237, Y => n658);
   U860 : NOR3X1 port map( A => n658, B => n220, C => n656, Y => n659);
   U861 : NAND2X1 port map( A => n660, B => n659, Y => n683);
   U862 : NAND2X1 port map( A => temp_6_port, B => n115, Y => n663);
   U863 : NAND3X1 port map( A => DATA_IN(6), B => n6, C => n684, Y => n662);
   U864 : INVX2 port map( A => n202, Y => n685);
   U865 : NAND3X1 port map( A => N526, B => n685, C => n684, Y => n661);
   U866 : NAND3X1 port map( A => n663, B => n662, C => n661, Y => n1179);
   U867 : NAND2X1 port map( A => temp_5_port, B => n115, Y => n666);
   U868 : NAND3X1 port map( A => DATA_IN(5), B => n6, C => n684, Y => n665);
   U869 : NAND3X1 port map( A => N525, B => n685, C => n93, Y => n664);
   U870 : NAND3X1 port map( A => n666, B => n665, C => n664, Y => n1178);
   U871 : NAND2X1 port map( A => temp_4_port, B => n91, Y => n669);
   U872 : NAND3X1 port map( A => DATA_IN(4), B => n6, C => n93, Y => n668);
   U873 : NAND3X1 port map( A => N524, B => n685, C => n684, Y => n667);
   U874 : NAND3X1 port map( A => n669, B => n668, C => n667, Y => n1177);
   U875 : NAND2X1 port map( A => temp_3_port, B => n91, Y => n672);
   U876 : NAND3X1 port map( A => DATA_IN(3), B => n6, C => n93, Y => n671);
   U877 : NAND3X1 port map( A => N523, B => n685, C => n93, Y => n670);
   U878 : NAND3X1 port map( A => n672, B => n671, C => n670, Y => n1176);
   U879 : NAND2X1 port map( A => temp_2_port, B => n115, Y => n675);
   U880 : NAND3X1 port map( A => DATA_IN(2), B => n6, C => n684, Y => n674);
   U881 : NAND3X1 port map( A => N522, B => n685, C => n93, Y => n673);
   U882 : NAND3X1 port map( A => n675, B => n674, C => n673, Y => n1175);
   U883 : NAND2X1 port map( A => temp_1_port, B => n91, Y => n678);
   U884 : NAND3X1 port map( A => DATA_IN(1), B => n6, C => n93, Y => n677);
   U885 : NAND3X1 port map( A => N521, B => n685, C => n684, Y => n676);
   U886 : NAND3X1 port map( A => n678, B => n677, C => n676, Y => n1174);
   U887 : NAND2X1 port map( A => temp_0_port, B => n76, Y => n682);
   U888 : NAND3X1 port map( A => DATA_IN(0), B => n6, C => n684, Y => n681);
   U889 : NAND3X1 port map( A => N520, B => n685, C => n93, Y => n680);
   U890 : NAND3X1 port map( A => n682, B => n681, C => n680, Y => n1173);
   U891 : NAND2X1 port map( A => temp_7_port, B => n115, Y => n688);
   U892 : NAND3X1 port map( A => DATA_IN(7), B => n6, C => n93, Y => n687);
   U893 : NAND3X1 port map( A => N527, B => n685, C => n684, Y => n686);
   U894 : NAND3X1 port map( A => n688, B => n687, C => n686, Y => n1180);
   U895 : NOR2X1 port map( A => n692, B => n690, Y => n1020);
   U896 : NAND2X1 port map( A => n104, B => n1018, Y => n1097);
   U897 : INVX2 port map( A => N413, Y => n750);
   U898 : NAND2X1 port map( A => prefillCounter_6_port, B => n1094, Y => n748);
   U899 : OAI21X1 port map( A => n61, B => n750, C => n748, Y => n1145);
   U900 : INVX2 port map( A => N412, Y => n754);
   U901 : NAND2X1 port map( A => n1094, B => prefillCounter_5_port, Y => n752);
   U902 : OAI21X1 port map( A => n61, B => n754, C => n752, Y => n1144);
   U903 : INVX2 port map( A => N411, Y => n758);
   U904 : NAND2X1 port map( A => prefillCounter_4_port, B => n1094, Y => n756);
   U905 : OAI21X1 port map( A => n62, B => n758, C => n756, Y => n1143);
   U906 : INVX2 port map( A => N410, Y => n765);
   U907 : NAND2X1 port map( A => prefillCounter_3_port, B => n1094, Y => n760);
   U908 : OAI21X1 port map( A => n62, B => n765, C => n760, Y => n1142);
   U909 : INVX2 port map( A => N409, Y => n767);
   U914 : NAND2X1 port map( A => prefillCounter_2_port, B => n1094, Y => n766);
   U915 : OAI21X1 port map( A => n62, B => n767, C => n766, Y => n1141);
   U916 : INVX2 port map( A => N408, Y => n769);
   U917 : NAND2X1 port map( A => prefillCounter_1_port, B => n1094, Y => n768);
   U918 : OAI21X1 port map( A => n62, B => n769, C => n768, Y => n1140);
   U920 : INVX2 port map( A => N414, Y => n772);
   U921 : NAND2X1 port map( A => prefillCounter_7_port, B => n1094, Y => n771);
   U922 : OAI21X1 port map( A => n61, B => n772, C => n771, Y => n1139);
   U923 : INVX2 port map( A => KEY(7), Y => n783);
   U932 : NOR2X1 port map( A => n89, B => n773, Y => n774);
   U933 : MUX2X1 port map( B => n784, A => n783, S => n138, Y => n1181);
   U934 : INVX2 port map( A => KEY(15), Y => n785);
   U935 : MUX2X1 port map( B => n786, A => n785, S => n141, Y => n1182);
   U936 : INVX2 port map( A => KEY(0), Y => n787);
   U937 : MUX2X1 port map( B => n788, A => n787, S => n138, Y => n1183);
   U938 : INVX2 port map( A => KEY(1), Y => n789);
   U939 : MUX2X1 port map( B => n790, A => n789, S => n138, Y => n1184);
   U940 : INVX2 port map( A => KEY(2), Y => n791);
   U941 : MUX2X1 port map( B => n864, A => n791, S => n143, Y => n1185);
   U942 : INVX2 port map( A => KEY(3), Y => n865);
   U943 : MUX2X1 port map( B => n866, A => n865, S => n138, Y => n1186);
   U944 : INVX2 port map( A => KEY(4), Y => n867);
   U945 : MUX2X1 port map( B => n868, A => n867, S => n142, Y => n1187);
   U946 : INVX2 port map( A => KEY(5), Y => n869);
   U947 : MUX2X1 port map( B => n870, A => n869, S => n142, Y => n1188);
   U948 : INVX2 port map( A => KEY(6), Y => n871);
   U949 : MUX2X1 port map( B => n883, A => n871, S => n140, Y => n1189);
   U950 : INVX2 port map( A => KEY(14), Y => n884);
   U951 : MUX2X1 port map( B => n885, A => n884, S => n143, Y => n1190);
   U952 : INVX2 port map( A => KEY(13), Y => n886);
   U953 : MUX2X1 port map( B => n887, A => n886, S => n139, Y => n1191);
   U954 : INVX2 port map( A => KEY(12), Y => n888);
   U955 : MUX2X1 port map( B => n889, A => n888, S => n139, Y => n1192);
   U956 : INVX2 port map( A => KEY(11), Y => n890);
   U957 : MUX2X1 port map( B => n898, A => n890, S => n139, Y => n1193);
   U958 : INVX2 port map( A => KEY(10), Y => n916);
   U959 : MUX2X1 port map( B => n917, A => n916, S => n140, Y => n1194);
   U960 : INVX2 port map( A => KEY(9), Y => n918);
   U961 : MUX2X1 port map( B => n919, A => n918, S => n142, Y => n1195);
   U962 : INVX2 port map( A => KEY(8), Y => n920);
   U963 : MUX2X1 port map( B => n921, A => n920, S => n140, Y => n1196);
   U964 : INVX2 port map( A => KEY(23), Y => n922);
   U965 : MUX2X1 port map( B => n923, A => n922, S => n138, Y => n1197);
   U966 : INVX2 port map( A => KEY(22), Y => n924);
   U967 : MUX2X1 port map( B => n925, A => n924, S => n138, Y => n1198);
   U968 : INVX2 port map( A => KEY(21), Y => n926);
   U969 : MUX2X1 port map( B => n927, A => n926, S => n138, Y => n1199);
   U970 : INVX2 port map( A => KEY(20), Y => n928);
   U971 : MUX2X1 port map( B => n929, A => n928, S => n138, Y => n1200);
   U972 : INVX2 port map( A => KEY(19), Y => n930);
   U973 : MUX2X1 port map( B => n931, A => n930, S => n138, Y => n1201);
   U974 : INVX2 port map( A => KEY(18), Y => n932);
   U975 : MUX2X1 port map( B => n933, A => n932, S => n141, Y => n1202);
   U976 : INVX2 port map( A => KEY(17), Y => n934);
   U977 : MUX2X1 port map( B => n935, A => n934, S => n139, Y => n1203);
   U978 : INVX2 port map( A => KEY(16), Y => n936);
   U979 : MUX2X1 port map( B => n937, A => n936, S => n138, Y => n1204);
   U980 : INVX2 port map( A => KEY(31), Y => n938);
   U981 : MUX2X1 port map( B => n939, A => n938, S => n139, Y => n1205);
   U982 : INVX2 port map( A => KEY(30), Y => n940);
   U983 : MUX2X1 port map( B => n941, A => n940, S => n143, Y => n1206);
   U984 : INVX2 port map( A => KEY(29), Y => n942);
   U985 : MUX2X1 port map( B => n943, A => n942, S => n141, Y => n1207);
   U986 : INVX2 port map( A => KEY(28), Y => n944);
   U987 : MUX2X1 port map( B => n945, A => n944, S => n143, Y => n1208);
   U988 : INVX2 port map( A => KEY(27), Y => n946);
   U989 : MUX2X1 port map( B => n947, A => n946, S => n141, Y => n1209);
   U990 : INVX2 port map( A => KEY(26), Y => n948);
   U991 : MUX2X1 port map( B => n949, A => n948, S => n140, Y => n1210);
   U992 : INVX2 port map( A => KEY(25), Y => n950);
   U993 : MUX2X1 port map( B => n951, A => n950, S => n143, Y => n1211);
   U994 : INVX2 port map( A => KEY(24), Y => n952);
   U995 : MUX2X1 port map( B => n953, A => n952, S => n142, Y => n1212);
   U996 : INVX2 port map( A => keyTable_4_7_port, Y => n955);
   U997 : INVX2 port map( A => KEY(39), Y => n954);
   U998 : MUX2X1 port map( B => n955, A => n954, S => n142, Y => n1213);
   U999 : INVX2 port map( A => keyTable_4_6_port, Y => n957);
   U1000 : INVX2 port map( A => KEY(38), Y => n956);
   U1001 : MUX2X1 port map( B => n957, A => n956, S => n140, Y => n1214);
   U1002 : INVX2 port map( A => keyTable_4_5_port, Y => n959);
   U1003 : INVX2 port map( A => KEY(37), Y => n958);
   U1004 : MUX2X1 port map( B => n959, A => n958, S => n142, Y => n1215);
   U1005 : INVX2 port map( A => keyTable_4_4_port, Y => n961);
   U1006 : INVX2 port map( A => KEY(36), Y => n960);
   U1007 : MUX2X1 port map( B => n961, A => n960, S => n140, Y => n1216);
   U1008 : INVX2 port map( A => keyTable_4_3_port, Y => n963);
   U1009 : INVX2 port map( A => KEY(35), Y => n962);
   U1010 : MUX2X1 port map( B => n963, A => n962, S => n139, Y => n1217);
   U1011 : INVX2 port map( A => keyTable_4_2_port, Y => n965);
   U1012 : INVX2 port map( A => KEY(34), Y => n964);
   U1013 : MUX2X1 port map( B => n965, A => n964, S => n143, Y => n1218);
   U1014 : INVX2 port map( A => keyTable_4_1_port, Y => n967);
   U1015 : INVX2 port map( A => KEY(33), Y => n966);
   U1016 : MUX2X1 port map( B => n967, A => n966, S => n142, Y => n1219);
   U1017 : INVX2 port map( A => keyTable_4_0_port, Y => n969);
   U1018 : INVX2 port map( A => KEY(32), Y => n968);
   U1019 : MUX2X1 port map( B => n969, A => n968, S => n141, Y => n1220);
   U1020 : INVX2 port map( A => keyTable_5_7_port, Y => n971);
   U1021 : INVX2 port map( A => KEY(47), Y => n970);
   U1022 : MUX2X1 port map( B => n971, A => n970, S => n139, Y => n1221);
   U1023 : INVX2 port map( A => keyTable_5_6_port, Y => n973);
   U1024 : INVX2 port map( A => KEY(46), Y => n972);
   U1025 : MUX2X1 port map( B => n973, A => n972, S => n141, Y => n1222);
   U1026 : INVX2 port map( A => keyTable_5_5_port, Y => n975);
   U1027 : INVX2 port map( A => KEY(45), Y => n974);
   U1028 : MUX2X1 port map( B => n975, A => n974, S => n141, Y => n1223);
   U1029 : INVX2 port map( A => keyTable_5_4_port, Y => n977);
   U1030 : INVX2 port map( A => KEY(44), Y => n976);
   U1031 : MUX2X1 port map( B => n977, A => n976, S => n139, Y => n1224);
   U1032 : INVX2 port map( A => keyTable_5_3_port, Y => n979);
   U1033 : INVX2 port map( A => KEY(43), Y => n978);
   U1034 : MUX2X1 port map( B => n979, A => n978, S => n141, Y => n1225);
   U1035 : INVX2 port map( A => keyTable_5_2_port, Y => n981);
   U1036 : INVX2 port map( A => KEY(42), Y => n980);
   U1037 : MUX2X1 port map( B => n981, A => n980, S => n141, Y => n1226);
   U1038 : INVX2 port map( A => keyTable_5_1_port, Y => n983);
   U1039 : INVX2 port map( A => KEY(41), Y => n982);
   U1040 : MUX2X1 port map( B => n983, A => n982, S => n141, Y => n1227);
   U1041 : INVX2 port map( A => keyTable_5_0_port, Y => n985);
   U1042 : INVX2 port map( A => KEY(40), Y => n984);
   U1043 : MUX2X1 port map( B => n985, A => n984, S => n143, Y => n1228);
   U1044 : INVX2 port map( A => keyTable_6_7_port, Y => n987);
   U1045 : INVX2 port map( A => KEY(55), Y => n986);
   U1046 : MUX2X1 port map( B => n987, A => n986, S => n140, Y => n1229);
   U1047 : INVX2 port map( A => keyTable_6_6_port, Y => n989);
   U1048 : INVX2 port map( A => KEY(54), Y => n988);
   U1049 : MUX2X1 port map( B => n989, A => n988, S => n143, Y => n1230);
   U1050 : INVX2 port map( A => keyTable_6_5_port, Y => n991);
   U1051 : INVX2 port map( A => KEY(53), Y => n990);
   U1052 : MUX2X1 port map( B => n991, A => n990, S => n141, Y => n1231);
   U1053 : INVX2 port map( A => keyTable_6_4_port, Y => n993);
   U1054 : INVX2 port map( A => KEY(52), Y => n992);
   U1055 : MUX2X1 port map( B => n993, A => n992, S => n139, Y => n1232);
   U1056 : INVX2 port map( A => keyTable_6_3_port, Y => n995);
   U1057 : INVX2 port map( A => KEY(51), Y => n994);
   U1058 : MUX2X1 port map( B => n995, A => n994, S => n143, Y => n1233);
   U1059 : INVX2 port map( A => keyTable_6_2_port, Y => n997);
   U1060 : INVX2 port map( A => KEY(50), Y => n996);
   U1061 : MUX2X1 port map( B => n997, A => n996, S => n142, Y => n1234);
   U1062 : INVX2 port map( A => keyTable_6_1_port, Y => n999);
   U1063 : INVX2 port map( A => KEY(49), Y => n998);
   U1064 : MUX2X1 port map( B => n999, A => n998, S => n140, Y => n1235);
   U1065 : INVX2 port map( A => keyTable_6_0_port, Y => n1001);
   U1066 : INVX2 port map( A => KEY(48), Y => n1000);
   U1067 : MUX2X1 port map( B => n1001, A => n1000, S => n140, Y => n1236);
   U1068 : INVX2 port map( A => keyTable_7_7_port, Y => n1003);
   U1069 : INVX2 port map( A => KEY(63), Y => n1002);
   U1070 : MUX2X1 port map( B => n1003, A => n1002, S => n140, Y => n1237);
   U1071 : INVX2 port map( A => keyTable_7_6_port, Y => n1005);
   U1072 : INVX2 port map( A => KEY(62), Y => n1004);
   U1073 : MUX2X1 port map( B => n1005, A => n1004, S => n139, Y => n1238);
   U1074 : INVX2 port map( A => keyTable_7_5_port, Y => n1007);
   U1075 : INVX2 port map( A => KEY(61), Y => n1006);
   U1076 : MUX2X1 port map( B => n1007, A => n1006, S => n142, Y => n1239);
   U1077 : INVX2 port map( A => keyTable_7_4_port, Y => n1009);
   U1078 : INVX2 port map( A => KEY(60), Y => n1008);
   U1079 : MUX2X1 port map( B => n1009, A => n1008, S => n143, Y => n1240);
   U1080 : INVX2 port map( A => keyTable_7_3_port, Y => n1011);
   U1081 : INVX2 port map( A => KEY(59), Y => n1010);
   U1082 : MUX2X1 port map( B => n1011, A => n1010, S => n143, Y => n1241);
   U1083 : INVX2 port map( A => keyTable_7_2_port, Y => n1013);
   U1084 : INVX2 port map( A => KEY(58), Y => n1012);
   U1085 : MUX2X1 port map( B => n1013, A => n1012, S => n139, Y => n1242);
   U1086 : INVX2 port map( A => keyTable_7_1_port, Y => n1015);
   U1087 : INVX2 port map( A => KEY(57), Y => n1014);
   U1088 : MUX2X1 port map( B => n1015, A => n1014, S => n140, Y => n1243);
   U1089 : INVX2 port map( A => keyTable_7_0_port, Y => n1017);
   U1090 : INVX2 port map( A => KEY(56), Y => n1016);
   U1091 : MUX2X1 port map( B => n1017, A => n1016, S => n142, Y => n1244);
   U1092 : INVX2 port map( A => extratemp_0_port, Y => n1023);
   U1093 : INVX2 port map( A => DATA_IN(0), Y => n1022);
   U1094 : AOI21X1 port map( A => n88, B => n51, C => n1018, Y => n1019);
   U1095 : MUX2X1 port map( B => n1023, A => n1022, S => n1036, Y => n1126);
   U1096 : INVX2 port map( A => extratemp_1_port, Y => n1025);
   U1097 : INVX2 port map( A => DATA_IN(1), Y => n1024);
   U1098 : MUX2X1 port map( B => n1025, A => n1024, S => n1036, Y => n1127);
   U1099 : INVX2 port map( A => extratemp_2_port, Y => n1027);
   U1100 : INVX2 port map( A => DATA_IN(2), Y => n1026);
   U1101 : MUX2X1 port map( B => n1027, A => n1026, S => n1036, Y => n1128);
   U1102 : INVX2 port map( A => extratemp_3_port, Y => n1029);
   U1103 : INVX2 port map( A => DATA_IN(3), Y => n1028);
   U1104 : MUX2X1 port map( B => n1029, A => n1028, S => n1036, Y => n1129);
   U1105 : INVX2 port map( A => extratemp_4_port, Y => n1031);
   U1106 : INVX2 port map( A => DATA_IN(4), Y => n1030);
   U1107 : MUX2X1 port map( B => n1031, A => n1030, S => n1036, Y => n1130);
   U1108 : INVX2 port map( A => extratemp_5_port, Y => n1033);
   U1109 : INVX2 port map( A => DATA_IN(5), Y => n1032);
   U1110 : MUX2X1 port map( B => n1033, A => n1032, S => n1036, Y => n1131);
   U1111 : INVX2 port map( A => extratemp_6_port, Y => n1035);
   U1112 : INVX2 port map( A => DATA_IN(6), Y => n1034);
   U1113 : MUX2X1 port map( B => n1035, A => n1034, S => n1036, Y => n1132);
   U1114 : INVX2 port map( A => extratemp_7_port, Y => n1038);
   U1115 : INVX2 port map( A => DATA_IN(7), Y => n1037);
   U1116 : MUX2X1 port map( B => n1038, A => n1037, S => n1036, Y => n1133);
   U1117 : AOI21X1 port map( A => n1041, B => n1040, C => n1134, Y => n1049);
   U1118 : NAND2X1 port map( A => permuteComplete, B => n1042, Y => n1043);
   U1119 : NAND3X1 port map( A => n177, B => n121, C => n1043, Y => n1089);
   U1120 : INVX2 port map( A => n1089, Y => n1048);
   U1121 : OAI21X1 port map( A => n49, B => n209, C => n118, Y => n1045);
   U1122 : AOI22X1 port map( A => n1105, B => n1046, C => n51, D => n1045, Y =>
                           n1047);
   U1123 : NAND3X1 port map( A => n1049, B => n1048, C => n1047, Y => 
                           nextState_3_port);
   U1124 : OAI21X1 port map( A => n1054, B => n1051, C => n1050, Y => n1052);
   U1125 : NAND2X1 port map( A => n1053, B => n1052, Y => n1056);
   U1126 : NAND2X1 port map( A => permuteComplete, B => n1054, Y => n1055);
   U1127 : NAND2X1 port map( A => n1056, B => n1055, Y => n1154);
   U1128 : NAND3X1 port map( A => n1107, B => BYTE_READY, C => n1083, Y => 
                           n1060);
   U1129 : NAND2X1 port map( A => n1332, B => n1082, Y => n1059);
   U1130 : NAND2X1 port map( A => n154, B => n164, Y => n1058);
   U1131 : NAND3X1 port map( A => n1060, B => n1059, C => n1058, Y => n1062);
   U1132 : AOI21X1 port map( A => n1062, B => n1105, C => n1061, Y => n1067);
   U1133 : NAND2X1 port map( A => n342, B => n48, Y => n1064);
   U1134 : NOR3X1 port map( A => n1065, B => n1064, C => n1134, Y => n1066);
   U1135 : NAND3X1 port map( A => n203, B => n1067, C => n1066, Y => 
                           nextState_0_port);
   U1136 : NAND2X1 port map( A => n49, B => n164, Y => n1079);
   U1137 : INVX2 port map( A => n1334, Y => n1070);
   U1138 : NAND2X1 port map( A => n1071, B => n1070, Y => n1078);
   U1139 : NAND2X1 port map( A => n1074, B => n94, Y => n1075);
   U1140 : AOI21X1 port map( A => n1333, B => n1076, C => n1075, Y => n1077);
   U1141 : NAND3X1 port map( A => n1079, B => n1078, C => n1077, Y => 
                           nextState_4_port);
   U1142 : AND2X2 port map( A => n41, B => n74, Y => n1081);
   U1143 : MUX2X1 port map( B => n1041, A => n1081, S => n209, Y => n1093);
   U1144 : NAND2X1 port map( A => n1330, B => n1082, Y => n1085);
   U1145 : NAND2X1 port map( A => n1329, B => n1083, Y => n1084);
   U1146 : NAND2X1 port map( A => n1085, B => n1084, Y => n1086);
   U1147 : NAND2X1 port map( A => n1086, B => n1105, Y => n1092);
   U1148 : NAND2X1 port map( A => n170, B => n1087, Y => n1090);
   U1149 : NOR2X1 port map( A => n1090, B => n1089, Y => n1091);
   U1150 : NAND3X1 port map( A => n1093, B => n1092, C => n1091, Y => 
                           nextState_2_port);
   U1151 : INVX2 port map( A => N407, Y => n1096);
   U1152 : NAND2X1 port map( A => prefillCounter_0_port, B => n1094, Y => n1095
                           );
   U1153 : OAI21X1 port map( A => n61, B => n1096, C => n1095, Y => n1138);
   U1154 : INVX2 port map( A => KEY_ERROR, Y => n1105);
   U1155 : INVX2 port map( A => BYTE_READY, Y => n1106);
   U1156 : INVX2 port map( A => n1331, Y => n1107);
   U1157 : INVX2 port map( A => OPCODE(1), Y => n1108);
   U1158 : INVX2 port map( A => OPCODE(0), Y => n1109);
   n1136 <= '0';
   n1137 <= '0';

end SYN_bksa;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity transmitter_block_0 is

   port( PRGA_OUT : in std_logic_vector (7 downto 0);  clk, p_ready : in 
         std_logic;  prga_opcode : in std_logic_vector (1 downto 0);  rst : in 
         std_logic;  SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE : out std_logic);

end transmitter_block_0;

architecture SYN_struct of transmitter_block_0 is

   component tx_timer_0
      port( CLK, RST, SENDING : in std_logic;  SHIFT_ENABLE_R, SHIFT_ENABLE_E :
            out std_logic);
   end component;
   
   component tx_tcu_0
      port( clk, rst, p_ready, t_bitstuff : in std_logic;  PRGA_OUT : in 
            std_logic_vector (7 downto 0);  prga_opcode : in std_logic_vector 
            (1 downto 0);  t_crc : in std_logic_vector (15 downto 0);  sending,
            EOP, next_byte : out std_logic;  send_data : out std_logic_vector 
            (7 downto 0);  t_strobe : out std_logic);
   end component;
   
   component tx_shiftreg_0
      port( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe : in std_logic;  
            send_data : in std_logic_vector (7 downto 0);  d_encode : out 
            std_logic);
   end component;
   
   component tx_encode_0
      port( clk, rst, SHIFT_ENABLE_E, d_encode, EOP : in std_logic;  t_bitstuff
            , dp_tx_out, dm_tx_out : out std_logic);
   end component;
   
   component tx_CRC_CALC_0
      port( CLK, RST, EOP, T_STROBE : in std_logic;  PRGA_OPCODE : in 
            std_logic_vector (1 downto 0);  PRGA_OUT : in std_logic_vector (7 
            downto 0);  TX_CRC : out std_logic_vector (15 downto 0));
   end component;
   
   signal SENDING_port, t_strobe, EOP, TX_CRC_15_port, TX_CRC_14_port, 
      TX_CRC_13_port, TX_CRC_12_port, TX_CRC_11_port, TX_CRC_10_port, 
      TX_CRC_9_port, TX_CRC_8_port, TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port
      , TX_CRC_4_port, TX_CRC_3_port, TX_CRC_2_port, TX_CRC_1_port, 
      TX_CRC_0_port, SHIFT_ENABLE_E, d_encode, t_bitstuff, SHIFT_ENABLE_R, 
      send_data_7_port, send_data_6_port, send_data_5_port, send_data_4_port, 
      send_data_3_port, send_data_2_port, send_data_1_port, send_data_0_port : 
      std_logic;

begin
   SENDING <= SENDING_port;
   
   U_1 : tx_CRC_CALC_0 port map( CLK => clk, RST => rst, EOP => EOP, T_STROBE 
                           => t_strobe, PRGA_OPCODE(1) => prga_opcode(1), 
                           PRGA_OPCODE(0) => prga_opcode(0), PRGA_OUT(7) => 
                           PRGA_OUT(7), PRGA_OUT(6) => PRGA_OUT(6), PRGA_OUT(5)
                           => PRGA_OUT(5), PRGA_OUT(4) => PRGA_OUT(4), 
                           PRGA_OUT(3) => PRGA_OUT(3), PRGA_OUT(2) => 
                           PRGA_OUT(2), PRGA_OUT(1) => PRGA_OUT(1), PRGA_OUT(0)
                           => PRGA_OUT(0), TX_CRC(15) => TX_CRC_15_port, 
                           TX_CRC(14) => TX_CRC_14_port, TX_CRC(13) => 
                           TX_CRC_13_port, TX_CRC(12) => TX_CRC_12_port, 
                           TX_CRC(11) => TX_CRC_11_port, TX_CRC(10) => 
                           TX_CRC_10_port, TX_CRC(9) => TX_CRC_9_port, 
                           TX_CRC(8) => TX_CRC_8_port, TX_CRC(7) => 
                           TX_CRC_7_port, TX_CRC(6) => TX_CRC_6_port, TX_CRC(5)
                           => TX_CRC_5_port, TX_CRC(4) => TX_CRC_4_port, 
                           TX_CRC(3) => TX_CRC_3_port, TX_CRC(2) => 
                           TX_CRC_2_port, TX_CRC(1) => TX_CRC_1_port, TX_CRC(0)
                           => TX_CRC_0_port);
   U_0 : tx_encode_0 port map( clk => clk, rst => rst, SHIFT_ENABLE_E => 
                           SHIFT_ENABLE_E, d_encode => d_encode, EOP => EOP, 
                           t_bitstuff => t_bitstuff, dp_tx_out => dp_tx_out, 
                           dm_tx_out => dm_tx_out);
   U_2 : tx_shiftreg_0 port map( clk => clk, rst => rst, SHIFT_ENABLE_R => 
                           SHIFT_ENABLE_R, t_bitstuff => t_bitstuff, t_strobe 
                           => t_strobe, send_data(7) => send_data_7_port, 
                           send_data(6) => send_data_6_port, send_data(5) => 
                           send_data_5_port, send_data(4) => send_data_4_port, 
                           send_data(3) => send_data_3_port, send_data(2) => 
                           send_data_2_port, send_data(1) => send_data_1_port, 
                           send_data(0) => send_data_0_port, d_encode => 
                           d_encode);
   U_3 : tx_tcu_0 port map( clk => clk, rst => rst, p_ready => p_ready, 
                           t_bitstuff => t_bitstuff, PRGA_OUT(7) => PRGA_OUT(7)
                           , PRGA_OUT(6) => PRGA_OUT(6), PRGA_OUT(5) => 
                           PRGA_OUT(5), PRGA_OUT(4) => PRGA_OUT(4), PRGA_OUT(3)
                           => PRGA_OUT(3), PRGA_OUT(2) => PRGA_OUT(2), 
                           PRGA_OUT(1) => PRGA_OUT(1), PRGA_OUT(0) => 
                           PRGA_OUT(0), prga_opcode(1) => prga_opcode(1), 
                           prga_opcode(0) => prga_opcode(0), t_crc(15) => 
                           TX_CRC_15_port, t_crc(14) => TX_CRC_14_port, 
                           t_crc(13) => TX_CRC_13_port, t_crc(12) => 
                           TX_CRC_12_port, t_crc(11) => TX_CRC_11_port, 
                           t_crc(10) => TX_CRC_10_port, t_crc(9) => 
                           TX_CRC_9_port, t_crc(8) => TX_CRC_8_port, t_crc(7) 
                           => TX_CRC_7_port, t_crc(6) => TX_CRC_6_port, 
                           t_crc(5) => TX_CRC_5_port, t_crc(4) => TX_CRC_4_port
                           , t_crc(3) => TX_CRC_3_port, t_crc(2) => 
                           TX_CRC_2_port, t_crc(1) => TX_CRC_1_port, t_crc(0) 
                           => TX_CRC_0_port, sending => SENDING_port, EOP => 
                           EOP, next_byte => NEXT_BYTE, send_data(7) => 
                           send_data_7_port, send_data(6) => send_data_6_port, 
                           send_data(5) => send_data_5_port, send_data(4) => 
                           send_data_4_port, send_data(3) => send_data_3_port, 
                           send_data(2) => send_data_2_port, send_data(1) => 
                           send_data_1_port, send_data(0) => send_data_0_port, 
                           t_strobe => t_strobe);
   U_4 : tx_timer_0 port map( CLK => clk, RST => rst, SENDING => SENDING_port, 
                           SHIFT_ENABLE_R => SHIFT_ENABLE_R, SHIFT_ENABLE_E => 
                           SHIFT_ENABLE_E);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity receiver_block_rewire_0 is

   port( CLK, DM1_RX, DP1_RX, RST : in std_logic;  BS_ERROR, CRC_ERROR, 
         EOP_external : out std_logic;  OPCODE : out std_logic_vector (1 downto
         0);  RCV_DATA : out std_logic_vector (7 downto 0);  R_ERROR, W_ENABLE 
         : out std_logic);

end receiver_block_rewire_0;

architecture SYN_struct of receiver_block_rewire_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component rx_timer_0
      port( CLK, RST, D_EDGE, RCVING : in std_logic;  SHIFT_ENABLE : out 
            std_logic);
   end component;
   
   component rx_shift_reg_0
      port( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF : in std_logic;  RCV_DATA 
            : out std_logic_vector (7 downto 0));
   end component;
   
   component rx_rcu_0
      port( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR : in 
            std_logic;  RX_CRC, RX_CHECK_CRC : in std_logic_vector (15 downto 
            0);  RCV_DATA : in std_logic_vector (7 downto 0);  RCVING, W_ENABLE
            , R_ERROR, CRC_ERROR : out std_logic;  OPCODE : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component rx_eopdetect_0
      port( DP1_RX, DM1_RX : in std_logic;  EOP : out std_logic);
   end component;
   
   component rx_edgedetect_0
      port( CLK, RST, DP1_RX : in std_logic;  D_EDGE : out std_logic);
   end component;
   
   component rx_decode_0
      port( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP : in std_logic;  D_ORIG, 
            BITSTUFF, BS_ERROR : out std_logic);
   end component;
   
   component rx_accumulator_0
      port( CLK, RST : in std_logic;  RCV_DATA : in std_logic_vector (7 downto 
            0);  W_ENABLE : in std_logic;  rx_CHECK_CRC : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component rx_CRC_CALC_0
      port( CLK, RST, W_ENABLE : in std_logic;  OPCODE : in std_logic_vector (1
            downto 0);  RCV_DATA : in std_logic_vector (7 downto 0);  RX_CRC : 
            out std_logic_vector (15 downto 0));
   end component;
   
   signal BS_ERROR_port, EOP_external_port, OPCODE_1_port, OPCODE_0_port, n8, 
      RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, RCV_DATA_3_port, 
      RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, n9, RX_CRC_15_port, 
      RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, RX_CRC_11_port, 
      RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, RX_CRC_7_port, 
      RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port, RX_CRC_2_port
      , RX_CRC_1_port, RX_CRC_0_port, rx_CHECK_CRC_15_port, 
      rx_CHECK_CRC_14_port, rx_CHECK_CRC_13_port, rx_CHECK_CRC_12_port, 
      rx_CHECK_CRC_11_port, rx_CHECK_CRC_10_port, rx_CHECK_CRC_9_port, 
      rx_CHECK_CRC_8_port, rx_CHECK_CRC_7_port, rx_CHECK_CRC_6_port, 
      rx_CHECK_CRC_5_port, rx_CHECK_CRC_4_port, rx_CHECK_CRC_3_port, 
      rx_CHECK_CRC_2_port, rx_CHECK_CRC_1_port, rx_CHECK_CRC_0_port, 
      SHIFT_ENABLE, BITSTUFF, D_ORIG, D_EDGE, RCVING, RCV_DATA_7_port, n2, n3, 
      n4, n5, n6 : std_logic;

begin
   BS_ERROR <= BS_ERROR_port;
   EOP_external <= EOP_external_port;
   OPCODE <= ( OPCODE_1_port, OPCODE_0_port );
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   U_2 : rx_CRC_CALC_0 port map( CLK => CLK, RST => RST, W_ENABLE => n4, 
                           OPCODE(1) => OPCODE_1_port, OPCODE(0) => 
                           OPCODE_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, RX_CRC(15) => 
                           RX_CRC_15_port, RX_CRC(14) => RX_CRC_14_port, 
                           RX_CRC(13) => RX_CRC_13_port, RX_CRC(12) => 
                           RX_CRC_12_port, RX_CRC(11) => RX_CRC_11_port, 
                           RX_CRC(10) => RX_CRC_10_port, RX_CRC(9) => 
                           RX_CRC_9_port, RX_CRC(8) => RX_CRC_8_port, RX_CRC(7)
                           => RX_CRC_7_port, RX_CRC(6) => RX_CRC_6_port, 
                           RX_CRC(5) => RX_CRC_5_port, RX_CRC(4) => 
                           RX_CRC_4_port, RX_CRC(3) => RX_CRC_3_port, RX_CRC(2)
                           => RX_CRC_2_port, RX_CRC(1) => RX_CRC_1_port, 
                           RX_CRC(0) => RX_CRC_0_port);
   U_3 : rx_accumulator_0 port map( CLK => CLK, RST => RST, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           W_ENABLE => n4, rx_CHECK_CRC(15) => 
                           rx_CHECK_CRC_15_port, rx_CHECK_CRC(14) => 
                           rx_CHECK_CRC_14_port, rx_CHECK_CRC(13) => 
                           rx_CHECK_CRC_13_port, rx_CHECK_CRC(12) => 
                           rx_CHECK_CRC_12_port, rx_CHECK_CRC(11) => 
                           rx_CHECK_CRC_11_port, rx_CHECK_CRC(10) => 
                           rx_CHECK_CRC_10_port, rx_CHECK_CRC(9) => 
                           rx_CHECK_CRC_9_port, rx_CHECK_CRC(8) => 
                           rx_CHECK_CRC_8_port, rx_CHECK_CRC(7) => 
                           rx_CHECK_CRC_7_port, rx_CHECK_CRC(6) => 
                           rx_CHECK_CRC_6_port, rx_CHECK_CRC(5) => 
                           rx_CHECK_CRC_5_port, rx_CHECK_CRC(4) => 
                           rx_CHECK_CRC_4_port, rx_CHECK_CRC(3) => 
                           rx_CHECK_CRC_3_port, rx_CHECK_CRC(2) => 
                           rx_CHECK_CRC_2_port, rx_CHECK_CRC(1) => 
                           rx_CHECK_CRC_1_port, rx_CHECK_CRC(0) => 
                           rx_CHECK_CRC_0_port);
   U_1 : rx_decode_0 port map( CLK => CLK, RST => RST, DP1_RX => DP1_RX, 
                           SHIFT_ENABLE => n5, EOP => EOP_external_port, D_ORIG
                           => D_ORIG, BITSTUFF => BITSTUFF, BS_ERROR => 
                           BS_ERROR_port);
   U_0 : rx_edgedetect_0 port map( CLK => CLK, RST => RST, DP1_RX => DP1_RX, 
                           D_EDGE => D_EDGE);
   U_4 : rx_eopdetect_0 port map( DP1_RX => DP1_RX, DM1_RX => DM1_RX, EOP => 
                           EOP_external_port);
   U_5 : rx_rcu_0 port map( CLK => CLK, RST => RST, D_EDGE => D_EDGE, EOP => 
                           EOP_external_port, SHIFT_ENABLE => SHIFT_ENABLE, 
                           BITSTUFF => BITSTUFF, BS_ERROR => BS_ERROR_port, 
                           RX_CRC(15) => RX_CRC_15_port, RX_CRC(14) => 
                           RX_CRC_14_port, RX_CRC(13) => RX_CRC_13_port, 
                           RX_CRC(12) => RX_CRC_12_port, RX_CRC(11) => 
                           RX_CRC_11_port, RX_CRC(10) => RX_CRC_10_port, 
                           RX_CRC(9) => RX_CRC_9_port, RX_CRC(8) => 
                           RX_CRC_8_port, RX_CRC(7) => RX_CRC_7_port, RX_CRC(6)
                           => RX_CRC_6_port, RX_CRC(5) => RX_CRC_5_port, 
                           RX_CRC(4) => RX_CRC_4_port, RX_CRC(3) => 
                           RX_CRC_3_port, RX_CRC(2) => RX_CRC_2_port, RX_CRC(1)
                           => RX_CRC_1_port, RX_CRC(0) => RX_CRC_0_port, 
                           RX_CHECK_CRC(15) => rx_CHECK_CRC_15_port, 
                           RX_CHECK_CRC(14) => rx_CHECK_CRC_14_port, 
                           RX_CHECK_CRC(13) => rx_CHECK_CRC_13_port, 
                           RX_CHECK_CRC(12) => rx_CHECK_CRC_12_port, 
                           RX_CHECK_CRC(11) => rx_CHECK_CRC_11_port, 
                           RX_CHECK_CRC(10) => rx_CHECK_CRC_10_port, 
                           RX_CHECK_CRC(9) => rx_CHECK_CRC_9_port, 
                           RX_CHECK_CRC(8) => rx_CHECK_CRC_8_port, 
                           RX_CHECK_CRC(7) => rx_CHECK_CRC_7_port, 
                           RX_CHECK_CRC(6) => rx_CHECK_CRC_6_port, 
                           RX_CHECK_CRC(5) => rx_CHECK_CRC_5_port, 
                           RX_CHECK_CRC(4) => rx_CHECK_CRC_4_port, 
                           RX_CHECK_CRC(3) => rx_CHECK_CRC_3_port, 
                           RX_CHECK_CRC(2) => rx_CHECK_CRC_2_port, 
                           RX_CHECK_CRC(1) => rx_CHECK_CRC_1_port, 
                           RX_CHECK_CRC(0) => rx_CHECK_CRC_0_port, RCV_DATA(7) 
                           => n8, RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) 
                           => RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, RCVING => RCVING, 
                           W_ENABLE => n9, R_ERROR => R_ERROR, CRC_ERROR => 
                           CRC_ERROR, OPCODE(1) => OPCODE_1_port, OPCODE(0) => 
                           OPCODE_0_port);
   U_6 : rx_shift_reg_0 port map( CLK => CLK, RST => RST, SHIFT_ENABLE => n3, 
                           D_ORIG => D_ORIG, BITSTUFF => BITSTUFF, RCV_DATA(7) 
                           => n8, RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) 
                           => RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port);
   U_7 : rx_timer_0 port map( CLK => CLK, RST => RST, D_EDGE => D_EDGE, RCVING 
                           => RCVING, SHIFT_ENABLE => SHIFT_ENABLE);
   U1 : BUFX2 port map( A => n8, Y => RCV_DATA_7_port);
   U2 : INVX1 port map( A => SHIFT_ENABLE, Y => n2);
   U3 : INVX1 port map( A => n2, Y => n3);
   U4 : INVX1 port map( A => n6, Y => n4);
   U5 : BUFX2 port map( A => SHIFT_ENABLE, Y => n5);
   U6 : INVX4 port map( A => n6, Y => W_ENABLE);
   U7 : INVX2 port map( A => n9, Y => n6);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity memoryblock_0 is

   port( CLK, NEXT_BYTE : in std_logic;  RCV_DATA : in std_logic_vector (7 
         downto 0);  RCV_OPCODE : in std_logic_vector (1 downto 0);  RST, 
         W_ENABLE, EOP : in std_logic;  EMPTY, FULL, B_READY : out std_logic;  
         PRGA_IN : out std_logic_vector (7 downto 0);  PRGA_OPCODE : out 
         std_logic_vector (1 downto 0));

end memoryblock_0;

architecture SYN_struct of memoryblock_0 is

   component RFIFO_0
      port( CLK, RST, W_ENABLE, R_ENABLE : in std_logic;  RCV_DATA : in 
            std_logic_vector (7 downto 0);  RCV_OPCODE : in std_logic_vector (1
            downto 0);  DATA : out std_logic_vector (7 downto 0);  OUT_OPCODE :
            out std_logic_vector (1 downto 0);  BYTE_COUNT : out 
            std_logic_vector (4 downto 0);  EMPTY, FULL : out std_logic);
   end component;
   
   component RBUFFER_0
      port( CLK, RST, NEXT_BYTE : in std_logic;  DATA : in std_logic_vector (7 
            downto 0);  OPCODE : in std_logic_vector (1 downto 0);  BYTE_COUNT 
            : in std_logic_vector (4 downto 0);  EOP : in std_logic;  B_READY, 
            R_ENABLE : out std_logic;  PRGA_IN : out std_logic_vector (7 downto
            0);  PRGA_OPCODE : out std_logic_vector (1 downto 0));
   end component;
   
   signal BYTE_COUNT_4_port, BYTE_COUNT_3_port, BYTE_COUNT_2_port, 
      BYTE_COUNT_1_port, BYTE_COUNT_0_port, DATA_7_port, DATA_6_port, 
      DATA_5_port, DATA_4_port, DATA_3_port, DATA_2_port, DATA_1_port, 
      DATA_0_port, OUT_OPCODE_1_port, OUT_OPCODE_0_port, R_ENABLE : std_logic;

begin
   
   U_0 : RBUFFER_0 port map( CLK => CLK, RST => RST, NEXT_BYTE => NEXT_BYTE, 
                           DATA(7) => DATA_7_port, DATA(6) => DATA_6_port, 
                           DATA(5) => DATA_5_port, DATA(4) => DATA_4_port, 
                           DATA(3) => DATA_3_port, DATA(2) => DATA_2_port, 
                           DATA(1) => DATA_1_port, DATA(0) => DATA_0_port, 
                           OPCODE(1) => OUT_OPCODE_1_port, OPCODE(0) => 
                           OUT_OPCODE_0_port, BYTE_COUNT(4) => 
                           BYTE_COUNT_4_port, BYTE_COUNT(3) => 
                           BYTE_COUNT_3_port, BYTE_COUNT(2) => 
                           BYTE_COUNT_2_port, BYTE_COUNT(1) => 
                           BYTE_COUNT_1_port, BYTE_COUNT(0) => 
                           BYTE_COUNT_0_port, EOP => EOP, B_READY => B_READY, 
                           R_ENABLE => R_ENABLE, PRGA_IN(7) => PRGA_IN(7), 
                           PRGA_IN(6) => PRGA_IN(6), PRGA_IN(5) => PRGA_IN(5), 
                           PRGA_IN(4) => PRGA_IN(4), PRGA_IN(3) => PRGA_IN(3), 
                           PRGA_IN(2) => PRGA_IN(2), PRGA_IN(1) => PRGA_IN(1), 
                           PRGA_IN(0) => PRGA_IN(0), PRGA_OPCODE(1) => 
                           PRGA_OPCODE(1), PRGA_OPCODE(0) => PRGA_OPCODE(0));
   U_1 : RFIFO_0 port map( CLK => CLK, RST => RST, W_ENABLE => W_ENABLE, 
                           R_ENABLE => R_ENABLE, RCV_DATA(7) => RCV_DATA(7), 
                           RCV_DATA(6) => RCV_DATA(6), RCV_DATA(5) => 
                           RCV_DATA(5), RCV_DATA(4) => RCV_DATA(4), RCV_DATA(3)
                           => RCV_DATA(3), RCV_DATA(2) => RCV_DATA(2), 
                           RCV_DATA(1) => RCV_DATA(1), RCV_DATA(0) => 
                           RCV_DATA(0), RCV_OPCODE(1) => RCV_OPCODE(1), 
                           RCV_OPCODE(0) => RCV_OPCODE(0), DATA(7) => 
                           DATA_7_port, DATA(6) => DATA_6_port, DATA(5) => 
                           DATA_5_port, DATA(4) => DATA_4_port, DATA(3) => 
                           DATA_3_port, DATA(2) => DATA_2_port, DATA(1) => 
                           DATA_1_port, DATA(0) => DATA_0_port, OUT_OPCODE(1) 
                           => OUT_OPCODE_1_port, OUT_OPCODE(0) => 
                           OUT_OPCODE_0_port, BYTE_COUNT(4) => 
                           BYTE_COUNT_4_port, BYTE_COUNT(3) => 
                           BYTE_COUNT_3_port, BYTE_COUNT(2) => 
                           BYTE_COUNT_2_port, BYTE_COUNT(1) => 
                           BYTE_COUNT_1_port, BYTE_COUNT(0) => 
                           BYTE_COUNT_0_port, EMPTY => EMPTY, FULL => FULL);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity EDBlock_0 is

   port( BYTE : in std_logic_vector (7 downto 0);  BYTE_READY, CLK : in 
         std_logic;  OPCODE : in std_logic_vector (1 downto 0);  RST, SERIAL_IN
         : in std_logic;  DATA_IN : in std_logic_vector (7 downto 0);  
         KEY_ERROR, PARITY_ERROR, PDATA_READY : out std_logic;  PROCESSED_DATA 
         : out std_logic_vector (7 downto 0);  PROG_ERROR, RBUF_FULL, W_ENABLE,
         R_ENABLE : out std_logic;  DATA, ADDR : out std_logic_vector (7 downto
         0));

end EDBlock_0;

architecture SYN_struct of EDBlock_0 is

   component uart_rcv_block_0
      port( CLK, RST, SERIAL_IN : in std_logic;  KEY_ERROR, PROG_ERROR : out 
            std_logic;  PLAINKEY : out std_logic_vector (63 downto 0);  
            RBUF_FULL, PARITY_ERROR : out std_logic);
   end component;
   
   component KSA_0
      port( KEY : in std_logic_vector (63 downto 0);  CLK, RST, KEY_ERROR, 
            BYTE_READY : in std_logic;  BYTE : in std_logic_vector (7 downto 0)
            ;  OPCODE : in std_logic_vector (1 downto 0);  DATA_IN : in 
            std_logic_vector (7 downto 0);  PROCESSED_DATA : out 
            std_logic_vector (7 downto 0);  PDATA_READY, W_ENABLE, R_ENABLE : 
            out std_logic;  ADDR, DATA : out std_logic_vector (7 downto 0));
   end component;
   
   signal KEY_ERROR_port, PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port,
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port : std_logic;

begin
   KEY_ERROR <= KEY_ERROR_port;
   
   U_0 : KSA_0 port map( KEY(63) => PLAINKEY_63_port, KEY(62) => 
                           PLAINKEY_62_port, KEY(61) => PLAINKEY_61_port, 
                           KEY(60) => PLAINKEY_60_port, KEY(59) => 
                           PLAINKEY_59_port, KEY(58) => PLAINKEY_58_port, 
                           KEY(57) => PLAINKEY_57_port, KEY(56) => 
                           PLAINKEY_56_port, KEY(55) => PLAINKEY_55_port, 
                           KEY(54) => PLAINKEY_54_port, KEY(53) => 
                           PLAINKEY_53_port, KEY(52) => PLAINKEY_52_port, 
                           KEY(51) => PLAINKEY_51_port, KEY(50) => 
                           PLAINKEY_50_port, KEY(49) => PLAINKEY_49_port, 
                           KEY(48) => PLAINKEY_48_port, KEY(47) => 
                           PLAINKEY_47_port, KEY(46) => PLAINKEY_46_port, 
                           KEY(45) => PLAINKEY_45_port, KEY(44) => 
                           PLAINKEY_44_port, KEY(43) => PLAINKEY_43_port, 
                           KEY(42) => PLAINKEY_42_port, KEY(41) => 
                           PLAINKEY_41_port, KEY(40) => PLAINKEY_40_port, 
                           KEY(39) => PLAINKEY_39_port, KEY(38) => 
                           PLAINKEY_38_port, KEY(37) => PLAINKEY_37_port, 
                           KEY(36) => PLAINKEY_36_port, KEY(35) => 
                           PLAINKEY_35_port, KEY(34) => PLAINKEY_34_port, 
                           KEY(33) => PLAINKEY_33_port, KEY(32) => 
                           PLAINKEY_32_port, KEY(31) => PLAINKEY_31_port, 
                           KEY(30) => PLAINKEY_30_port, KEY(29) => 
                           PLAINKEY_29_port, KEY(28) => PLAINKEY_28_port, 
                           KEY(27) => PLAINKEY_27_port, KEY(26) => 
                           PLAINKEY_26_port, KEY(25) => PLAINKEY_25_port, 
                           KEY(24) => PLAINKEY_24_port, KEY(23) => 
                           PLAINKEY_23_port, KEY(22) => PLAINKEY_22_port, 
                           KEY(21) => PLAINKEY_21_port, KEY(20) => 
                           PLAINKEY_20_port, KEY(19) => PLAINKEY_19_port, 
                           KEY(18) => PLAINKEY_18_port, KEY(17) => 
                           PLAINKEY_17_port, KEY(16) => PLAINKEY_16_port, 
                           KEY(15) => PLAINKEY_15_port, KEY(14) => 
                           PLAINKEY_14_port, KEY(13) => PLAINKEY_13_port, 
                           KEY(12) => PLAINKEY_12_port, KEY(11) => 
                           PLAINKEY_11_port, KEY(10) => PLAINKEY_10_port, 
                           KEY(9) => PLAINKEY_9_port, KEY(8) => PLAINKEY_8_port
                           , KEY(7) => PLAINKEY_7_port, KEY(6) => 
                           PLAINKEY_6_port, KEY(5) => PLAINKEY_5_port, KEY(4) 
                           => PLAINKEY_4_port, KEY(3) => PLAINKEY_3_port, 
                           KEY(2) => PLAINKEY_2_port, KEY(1) => PLAINKEY_1_port
                           , KEY(0) => PLAINKEY_0_port, CLK => CLK, RST => RST,
                           KEY_ERROR => KEY_ERROR_port, BYTE_READY => 
                           BYTE_READY, BYTE(7) => BYTE(7), BYTE(6) => BYTE(6), 
                           BYTE(5) => BYTE(5), BYTE(4) => BYTE(4), BYTE(3) => 
                           BYTE(3), BYTE(2) => BYTE(2), BYTE(1) => BYTE(1), 
                           BYTE(0) => BYTE(0), OPCODE(1) => OPCODE(1), 
                           OPCODE(0) => OPCODE(0), DATA_IN(7) => DATA_IN(7), 
                           DATA_IN(6) => DATA_IN(6), DATA_IN(5) => DATA_IN(5), 
                           DATA_IN(4) => DATA_IN(4), DATA_IN(3) => DATA_IN(3), 
                           DATA_IN(2) => DATA_IN(2), DATA_IN(1) => DATA_IN(1), 
                           DATA_IN(0) => DATA_IN(0), PROCESSED_DATA(7) => 
                           PROCESSED_DATA(7), PROCESSED_DATA(6) => 
                           PROCESSED_DATA(6), PROCESSED_DATA(5) => 
                           PROCESSED_DATA(5), PROCESSED_DATA(4) => 
                           PROCESSED_DATA(4), PROCESSED_DATA(3) => 
                           PROCESSED_DATA(3), PROCESSED_DATA(2) => 
                           PROCESSED_DATA(2), PROCESSED_DATA(1) => 
                           PROCESSED_DATA(1), PROCESSED_DATA(0) => 
                           PROCESSED_DATA(0), PDATA_READY => PDATA_READY, 
                           W_ENABLE => W_ENABLE, R_ENABLE => R_ENABLE, ADDR(7) 
                           => ADDR(7), ADDR(6) => ADDR(6), ADDR(5) => ADDR(5), 
                           ADDR(4) => ADDR(4), ADDR(3) => ADDR(3), ADDR(2) => 
                           ADDR(2), ADDR(1) => ADDR(1), ADDR(0) => ADDR(0), 
                           DATA(7) => DATA(7), DATA(6) => DATA(6), DATA(5) => 
                           DATA(5), DATA(4) => DATA(4), DATA(3) => DATA(3), 
                           DATA(2) => DATA(2), DATA(1) => DATA(1), DATA(0) => 
                           DATA(0));
   U_1 : uart_rcv_block_0 port map( CLK => CLK, RST => RST, SERIAL_IN => 
                           SERIAL_IN, KEY_ERROR => KEY_ERROR_port, PROG_ERROR 
                           => PROG_ERROR, PLAINKEY(63) => PLAINKEY_63_port, 
                           PLAINKEY(62) => PLAINKEY_62_port, PLAINKEY(61) => 
                           PLAINKEY_61_port, PLAINKEY(60) => PLAINKEY_60_port, 
                           PLAINKEY(59) => PLAINKEY_59_port, PLAINKEY(58) => 
                           PLAINKEY_58_port, PLAINKEY(57) => PLAINKEY_57_port, 
                           PLAINKEY(56) => PLAINKEY_56_port, PLAINKEY(55) => 
                           PLAINKEY_55_port, PLAINKEY(54) => PLAINKEY_54_port, 
                           PLAINKEY(53) => PLAINKEY_53_port, PLAINKEY(52) => 
                           PLAINKEY_52_port, PLAINKEY(51) => PLAINKEY_51_port, 
                           PLAINKEY(50) => PLAINKEY_50_port, PLAINKEY(49) => 
                           PLAINKEY_49_port, PLAINKEY(48) => PLAINKEY_48_port, 
                           PLAINKEY(47) => PLAINKEY_47_port, PLAINKEY(46) => 
                           PLAINKEY_46_port, PLAINKEY(45) => PLAINKEY_45_port, 
                           PLAINKEY(44) => PLAINKEY_44_port, PLAINKEY(43) => 
                           PLAINKEY_43_port, PLAINKEY(42) => PLAINKEY_42_port, 
                           PLAINKEY(41) => PLAINKEY_41_port, PLAINKEY(40) => 
                           PLAINKEY_40_port, PLAINKEY(39) => PLAINKEY_39_port, 
                           PLAINKEY(38) => PLAINKEY_38_port, PLAINKEY(37) => 
                           PLAINKEY_37_port, PLAINKEY(36) => PLAINKEY_36_port, 
                           PLAINKEY(35) => PLAINKEY_35_port, PLAINKEY(34) => 
                           PLAINKEY_34_port, PLAINKEY(33) => PLAINKEY_33_port, 
                           PLAINKEY(32) => PLAINKEY_32_port, PLAINKEY(31) => 
                           PLAINKEY_31_port, PLAINKEY(30) => PLAINKEY_30_port, 
                           PLAINKEY(29) => PLAINKEY_29_port, PLAINKEY(28) => 
                           PLAINKEY_28_port, PLAINKEY(27) => PLAINKEY_27_port, 
                           PLAINKEY(26) => PLAINKEY_26_port, PLAINKEY(25) => 
                           PLAINKEY_25_port, PLAINKEY(24) => PLAINKEY_24_port, 
                           PLAINKEY(23) => PLAINKEY_23_port, PLAINKEY(22) => 
                           PLAINKEY_22_port, PLAINKEY(21) => PLAINKEY_21_port, 
                           PLAINKEY(20) => PLAINKEY_20_port, PLAINKEY(19) => 
                           PLAINKEY_19_port, PLAINKEY(18) => PLAINKEY_18_port, 
                           PLAINKEY(17) => PLAINKEY_17_port, PLAINKEY(16) => 
                           PLAINKEY_16_port, PLAINKEY(15) => PLAINKEY_15_port, 
                           PLAINKEY(14) => PLAINKEY_14_port, PLAINKEY(13) => 
                           PLAINKEY_13_port, PLAINKEY(12) => PLAINKEY_12_port, 
                           PLAINKEY(11) => PLAINKEY_11_port, PLAINKEY(10) => 
                           PLAINKEY_10_port, PLAINKEY(9) => PLAINKEY_9_port, 
                           PLAINKEY(8) => PLAINKEY_8_port, PLAINKEY(7) => 
                           PLAINKEY_7_port, PLAINKEY(6) => PLAINKEY_6_port, 
                           PLAINKEY(5) => PLAINKEY_5_port, PLAINKEY(4) => 
                           PLAINKEY_4_port, PLAINKEY(3) => PLAINKEY_3_port, 
                           PLAINKEY(2) => PLAINKEY_2_port, PLAINKEY(1) => 
                           PLAINKEY_1_port, PLAINKEY(0) => PLAINKEY_0_port, 
                           RBUF_FULL => RBUF_FULL, PARITY_ERROR => PARITY_ERROR
                           );

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RMEDT_REWIRE_0 is

   port( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN : in std_logic;  DATA_IN : in 
         std_logic_vector (7 downto 0);  BS_ERROR, CRC_ERROR, EMPTY, FULL, 
         KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, R_ERROR, SENDING, 
         dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE : out std_logic;  DATA, 
         ADDR : out std_logic_vector (7 downto 0));

end RMEDT_REWIRE_0;

architecture SYN_struct of RMEDT_REWIRE_0 is

   component transmitter_block_0
      port( PRGA_OUT : in std_logic_vector (7 downto 0);  clk, p_ready : in 
            std_logic;  prga_opcode : in std_logic_vector (1 downto 0);  rst : 
            in std_logic;  SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE : out 
            std_logic);
   end component;
   
   component receiver_block_rewire_0
      port( CLK, DM1_RX, DP1_RX, RST : in std_logic;  BS_ERROR, CRC_ERROR, 
            EOP_external : out std_logic;  OPCODE : out std_logic_vector (1 
            downto 0);  RCV_DATA : out std_logic_vector (7 downto 0);  R_ERROR,
            W_ENABLE : out std_logic);
   end component;
   
   component memoryblock_0
      port( CLK, NEXT_BYTE : in std_logic;  RCV_DATA : in std_logic_vector (7 
            downto 0);  RCV_OPCODE : in std_logic_vector (1 downto 0);  RST, 
            W_ENABLE, EOP : in std_logic;  EMPTY, FULL, B_READY : out std_logic
            ;  PRGA_IN : out std_logic_vector (7 downto 0);  PRGA_OPCODE : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component EDBlock_0
      port( BYTE : in std_logic_vector (7 downto 0);  BYTE_READY, CLK : in 
            std_logic;  OPCODE : in std_logic_vector (1 downto 0);  RST, 
            SERIAL_IN : in std_logic;  DATA_IN : in std_logic_vector (7 downto 
            0);  KEY_ERROR, PARITY_ERROR, PDATA_READY : out std_logic;  
            PROCESSED_DATA : out std_logic_vector (7 downto 0);  PROG_ERROR, 
            RBUF_FULL, W_ENABLE, R_ENABLE : out std_logic;  DATA, ADDR : out 
            std_logic_vector (7 downto 0));
   end component;
   
   signal PRGA_IN_7_port, PRGA_IN_6_port, PRGA_IN_5_port, PRGA_IN_4_port, 
      PRGA_IN_3_port, PRGA_IN_2_port, PRGA_IN_1_port, PRGA_IN_0_port, B_READY, 
      PRGA_OPCODE_1_port, PRGA_OPCODE_0_port, PDATA_READY, 
      PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, PROCESSED_DATA_5_port, 
      PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, PROCESSED_DATA_2_port, 
      PROCESSED_DATA_1_port, PROCESSED_DATA_0_port, EOP_external, NEXT_BYTE, 
      RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      OPCODE_1_port, OPCODE_0_port, W_ENABLE : std_logic;

begin
   
   U_0 : EDBlock_0 port map( BYTE(7) => PRGA_IN_7_port, BYTE(6) => 
                           PRGA_IN_6_port, BYTE(5) => PRGA_IN_5_port, BYTE(4) 
                           => PRGA_IN_4_port, BYTE(3) => PRGA_IN_3_port, 
                           BYTE(2) => PRGA_IN_2_port, BYTE(1) => PRGA_IN_1_port
                           , BYTE(0) => PRGA_IN_0_port, BYTE_READY => B_READY, 
                           CLK => CLK, OPCODE(1) => PRGA_OPCODE_1_port, 
                           OPCODE(0) => PRGA_OPCODE_0_port, RST => RST, 
                           SERIAL_IN => SERIAL_IN, DATA_IN(7) => DATA_IN(7), 
                           DATA_IN(6) => DATA_IN(6), DATA_IN(5) => DATA_IN(5), 
                           DATA_IN(4) => DATA_IN(4), DATA_IN(3) => DATA_IN(3), 
                           DATA_IN(2) => DATA_IN(2), DATA_IN(1) => DATA_IN(1), 
                           DATA_IN(0) => DATA_IN(0), KEY_ERROR => KEY_ERROR, 
                           PARITY_ERROR => PARITY_ERROR, PDATA_READY => 
                           PDATA_READY, PROCESSED_DATA(7) => 
                           PROCESSED_DATA_7_port, PROCESSED_DATA(6) => 
                           PROCESSED_DATA_6_port, PROCESSED_DATA(5) => 
                           PROCESSED_DATA_5_port, PROCESSED_DATA(4) => 
                           PROCESSED_DATA_4_port, PROCESSED_DATA(3) => 
                           PROCESSED_DATA_3_port, PROCESSED_DATA(2) => 
                           PROCESSED_DATA_2_port, PROCESSED_DATA(1) => 
                           PROCESSED_DATA_1_port, PROCESSED_DATA(0) => 
                           PROCESSED_DATA_0_port, PROG_ERROR => PROG_ERROR, 
                           RBUF_FULL => RBUF_FULL, W_ENABLE => W_ENABLE_R, 
                           R_ENABLE => R_ENABLE, DATA(7) => DATA(7), DATA(6) =>
                           DATA(6), DATA(5) => DATA(5), DATA(4) => DATA(4), 
                           DATA(3) => DATA(3), DATA(2) => DATA(2), DATA(1) => 
                           DATA(1), DATA(0) => DATA(0), ADDR(7) => ADDR(7), 
                           ADDR(6) => ADDR(6), ADDR(5) => ADDR(5), ADDR(4) => 
                           ADDR(4), ADDR(3) => ADDR(3), ADDR(2) => ADDR(2), 
                           ADDR(1) => ADDR(1), ADDR(0) => ADDR(0));
   U_1 : memoryblock_0 port map( CLK => CLK, NEXT_BYTE => NEXT_BYTE, 
                           RCV_DATA(7) => RCV_DATA_7_port, RCV_DATA(6) => 
                           RCV_DATA_6_port, RCV_DATA(5) => RCV_DATA_5_port, 
                           RCV_DATA(4) => RCV_DATA_4_port, RCV_DATA(3) => 
                           RCV_DATA_3_port, RCV_DATA(2) => RCV_DATA_2_port, 
                           RCV_DATA(1) => RCV_DATA_1_port, RCV_DATA(0) => 
                           RCV_DATA_0_port, RCV_OPCODE(1) => OPCODE_1_port, 
                           RCV_OPCODE(0) => OPCODE_0_port, RST => RST, W_ENABLE
                           => W_ENABLE, EOP => EOP_external, EMPTY => EMPTY, 
                           FULL => FULL, B_READY => B_READY, PRGA_IN(7) => 
                           PRGA_IN_7_port, PRGA_IN(6) => PRGA_IN_6_port, 
                           PRGA_IN(5) => PRGA_IN_5_port, PRGA_IN(4) => 
                           PRGA_IN_4_port, PRGA_IN(3) => PRGA_IN_3_port, 
                           PRGA_IN(2) => PRGA_IN_2_port, PRGA_IN(1) => 
                           PRGA_IN_1_port, PRGA_IN(0) => PRGA_IN_0_port, 
                           PRGA_OPCODE(1) => PRGA_OPCODE_1_port, PRGA_OPCODE(0)
                           => PRGA_OPCODE_0_port);
   U_2 : receiver_block_rewire_0 port map( CLK => CLK, DM1_RX => DM1_RX, DP1_RX
                           => DP1_RX, RST => RST, BS_ERROR => BS_ERROR, 
                           CRC_ERROR => CRC_ERROR, EOP_external => EOP_external
                           , OPCODE(1) => OPCODE_1_port, OPCODE(0) => 
                           OPCODE_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, R_ERROR => R_ERROR, 
                           W_ENABLE => W_ENABLE);
   U_3 : transmitter_block_0 port map( PRGA_OUT(7) => PROCESSED_DATA_7_port, 
                           PRGA_OUT(6) => PROCESSED_DATA_6_port, PRGA_OUT(5) =>
                           PROCESSED_DATA_5_port, PRGA_OUT(4) => 
                           PROCESSED_DATA_4_port, PRGA_OUT(3) => 
                           PROCESSED_DATA_3_port, PRGA_OUT(2) => 
                           PROCESSED_DATA_2_port, PRGA_OUT(1) => 
                           PROCESSED_DATA_1_port, PRGA_OUT(0) => 
                           PROCESSED_DATA_0_port, clk => CLK, p_ready => 
                           PDATA_READY, prga_opcode(1) => PRGA_OPCODE_1_port, 
                           prga_opcode(0) => PRGA_OPCODE_0_port, rst => RST, 
                           SENDING => SENDING, dm_tx_out => dm_tx_out, 
                           dp_tx_out => dp_tx_out, NEXT_BYTE => NEXT_BYTE);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_timer_1 is

   port( CLK, RST, TIMER_TRIG : in std_logic;  STOP_RCVING, SHIFT_STROBE : out 
         std_logic);

end uart_timer_1;

architecture SYN_timerB of uart_timer_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component uart_timer_1_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal state_7_port, state_6_port, state_5_port, state_4_port, state_3_port,
      state_2_port, state_1_port, state_0_port, nextState_7_port, 
      nextState_6_port, nextState_5_port, nextState_4_port, nextState_3_port, 
      nextState_2_port, nextState_1_port, nextState_0_port, N26, N27, N28, N29,
      N30, N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, 
      n14, n15, n16, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n10, n17
      , n19, n20, n21, n22, n23, n24, n25, n26_port, n27_port, n28_port, 
      n29_port, n30_port, n31_port, n32_port, n33_port, n34 : std_logic;

begin
   
   nextState_reg_0_inst : DFFSR port map( D => n71, CLK => CLK, R => n17, S => 
                           n18, Q => nextState_0_port);
   nextState_reg_1_inst : DFFSR port map( D => n70, CLK => CLK, R => n17, S => 
                           n16, Q => nextState_1_port);
   nextState_reg_2_inst : DFFSR port map( D => n69, CLK => CLK, R => n17, S => 
                           n15, Q => nextState_2_port);
   nextState_reg_3_inst : DFFSR port map( D => n68, CLK => CLK, R => n17, S => 
                           n14, Q => nextState_3_port);
   nextState_reg_4_inst : DFFSR port map( D => n67, CLK => CLK, R => n17, S => 
                           n13, Q => nextState_4_port);
   nextState_reg_5_inst : DFFSR port map( D => n66, CLK => CLK, R => n17, S => 
                           n12, Q => nextState_5_port);
   nextState_reg_6_inst : DFFSR port map( D => n65, CLK => CLK, R => n17, S => 
                           n11, Q => nextState_6_port);
   STOP_RCVING_reg : DFFSR port map( D => n72, CLK => CLK, R => n17, S => n9, Q
                           => STOP_RCVING);
   state_reg_7_inst : DFFSR port map( D => nextState_7_port, CLK => CLK, R => 
                           n17, S => n8, Q => state_7_port);
   state_reg_6_inst : DFFSR port map( D => nextState_6_port, CLK => CLK, R => 
                           n17, S => n7, Q => state_6_port);
   state_reg_5_inst : DFFSR port map( D => nextState_5_port, CLK => CLK, R => 
                           n17, S => n6, Q => state_5_port);
   state_reg_4_inst : DFFSR port map( D => nextState_4_port, CLK => CLK, R => 
                           n17, S => n5, Q => state_4_port);
   state_reg_3_inst : DFFSR port map( D => nextState_3_port, CLK => CLK, R => 
                           n17, S => n4, Q => state_3_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n17, S => n3, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n17, S => n2, Q => state_1_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n17, S => n1, Q => state_0_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n18 <= '1';
   U21 : OR2X2 port map( A => state_7_port, B => n50, Y => n49);
   U38 : OAI21X1 port map( A => n20, B => n27_port, C => n35, Y => n64);
   U39 : NAND2X1 port map( A => N33, B => n36, Y => n35);
   U40 : OAI21X1 port map( A => n26_port, B => n20, C => n37, Y => n65);
   U41 : NAND2X1 port map( A => N32, B => n36, Y => n37);
   U42 : OAI21X1 port map( A => n25, B => n20, C => n38, Y => n66);
   U43 : NAND2X1 port map( A => N31, B => n36, Y => n38);
   U44 : OAI21X1 port map( A => n20, B => n24, C => n39, Y => n67);
   U45 : NAND2X1 port map( A => N30, B => n36, Y => n39);
   U46 : OAI21X1 port map( A => n23, B => n20, C => n40, Y => n68);
   U47 : NAND2X1 port map( A => N29, B => n36, Y => n40);
   U48 : OAI21X1 port map( A => n22, B => n20, C => n41, Y => n69);
   U49 : NAND2X1 port map( A => N28, B => n36, Y => n41);
   U50 : OAI21X1 port map( A => n20, B => n21, C => n42, Y => n70);
   U51 : NAND2X1 port map( A => N27, B => n36, Y => n42);
   U52 : OAI21X1 port map( A => n19, B => n20, C => n43, Y => n71);
   U53 : NAND2X1 port map( A => N26, B => n36, Y => n43);
   U54 : NOR2X1 port map( A => n44, B => n72, Y => n36);
   U55 : NOR2X1 port map( A => n72, B => TIMER_TRIG, Y => n44);
   U56 : NOR2X1 port map( A => n45, B => n46, Y => n72);
   U57 : NAND3X1 port map( A => nextState_6_port, B => nextState_5_port, C => 
                           n47, Y => n46);
   U58 : NOR2X1 port map( A => n22, B => n23, Y => n47);
   U59 : NAND3X1 port map( A => nextState_0_port, B => n21, C => n48, Y => n45)
                           ;
   U60 : NOR2X1 port map( A => nextState_7_port, B => nextState_4_port, Y => 
                           n48);
   U61 : NOR2X1 port map( A => state_0_port, B => n49, Y => SHIFT_STROBE);
   U62 : AOI21X1 port map( A => n51, B => n32_port, C => n52, Y => n50);
   U63 : OAI21X1 port map( A => n33_port, B => n53, C => n54, Y => n52);
   U64 : NAND3X1 port map( A => state_6_port, B => state_1_port, C => n55, Y =>
                           n54);
   U65 : AOI21X1 port map( A => n56, B => n57, C => state_3_port, Y => n55);
   U66 : NAND3X1 port map( A => n33_port, B => n31_port, C => state_4_port, Y 
                           => n57);
   U67 : NAND3X1 port map( A => state_2_port, B => n32_port, C => state_5_port,
                           Y => n56);
   U68 : NAND2X1 port map( A => state_4_port, B => n58, Y => n53);
   U69 : OAI21X1 port map( A => state_2_port, B => n28_port, C => n59, Y => n51
                           );
   U70 : NAND3X1 port map( A => state_2_port, B => n29_port, C => n30_port, Y 
                           => n59);
   U71 : OAI22X1 port map( A => state_6_port, B => n61, C => n29_port, D => n60
                           , Y => n58);
   U72 : NAND3X1 port map( A => n34, B => n31_port, C => state_3_port, Y => n60
                           );
   U73 : AOI22X1 port map( A => n62, B => state_1_port, C => n63, D => 
                           state_5_port, Y => n61);
   U74 : XOR2X1 port map( A => n34, B => state_3_port, Y => n63);
   U75 : NOR2X1 port map( A => state_5_port, B => state_3_port, Y => n62);
   add_39 : uart_timer_1_DW01_inc_0 port map( A(7) => nextState_7_port, A(6) =>
                           nextState_6_port, A(5) => nextState_5_port, A(4) => 
                           nextState_4_port, A(3) => nextState_3_port, A(2) => 
                           nextState_2_port, A(1) => nextState_1_port, A(0) => 
                           nextState_0_port, SUM(7) => N33, SUM(6) => N32, 
                           SUM(5) => N31, SUM(4) => N30, SUM(3) => N29, SUM(2) 
                           => N28, SUM(1) => N27, SUM(0) => N26);
   nextState_reg_7_inst : DFFSR port map( D => n64, CLK => CLK, R => n17, S => 
                           n10, Q => nextState_7_port);
   n10 <= '1';
   U19 : INVX2 port map( A => RST, Y => n17);
   U22 : INVX2 port map( A => nextState_0_port, Y => n19);
   U23 : INVX2 port map( A => n44, Y => n20);
   U24 : INVX2 port map( A => nextState_1_port, Y => n21);
   U25 : INVX2 port map( A => nextState_2_port, Y => n22);
   U26 : INVX2 port map( A => nextState_3_port, Y => n23);
   U27 : INVX2 port map( A => nextState_4_port, Y => n24);
   U28 : INVX2 port map( A => nextState_5_port, Y => n25);
   U29 : INVX2 port map( A => nextState_6_port, Y => n26_port);
   U30 : INVX2 port map( A => nextState_7_port, Y => n27_port);
   U31 : INVX2 port map( A => n58, Y => n28_port);
   U32 : INVX2 port map( A => state_6_port, Y => n29_port);
   U33 : INVX2 port map( A => n60, Y => n30_port);
   U34 : INVX2 port map( A => state_5_port, Y => n31_port);
   U35 : INVX2 port map( A => state_4_port, Y => n32_port);
   U36 : INVX2 port map( A => state_2_port, Y => n33_port);
   U37 : INVX2 port map( A => state_1_port, Y => n34);

end SYN_timerB;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity keyreg_1 is

   port( CLK, RST, SBE, OE, RBUF_FULL : in std_logic;  RCV_DATA : in 
         std_logic_vector (7 downto 0);  PLAINKEY : out std_logic_vector (63 
         downto 0);  KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR : out 
         std_logic);

end keyreg_1;

architecture SYN_keyb of keyreg_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component keyreg_1_DW01_add_1
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port, 
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port, CLR_RBUFF_port, state_3_port, state_2_port, state_1_port
      , state_0_port, parityError, keyCount_3_port, keyCount_2_port, 
      keyCount_1_port, keyCount_0_port, address_7_port, address_6_port, 
      address_5_port, address_4_port, address_3_port, address_2_port, 
      address_1_port, address_0_port, currentPlainKey_63_port, 
      currentPlainKey_62_port, currentPlainKey_61_port, currentPlainKey_60_port
      , currentPlainKey_59_port, currentPlainKey_58_port, 
      currentPlainKey_57_port, currentPlainKey_56_port, currentPlainKey_55_port
      , currentPlainKey_54_port, currentPlainKey_53_port, 
      currentPlainKey_52_port, currentPlainKey_51_port, currentPlainKey_50_port
      , currentPlainKey_49_port, currentPlainKey_48_port, 
      currentPlainKey_47_port, currentPlainKey_46_port, currentPlainKey_45_port
      , currentPlainKey_44_port, currentPlainKey_43_port, 
      currentPlainKey_42_port, currentPlainKey_41_port, currentPlainKey_40_port
      , currentPlainKey_39_port, currentPlainKey_38_port, 
      currentPlainKey_37_port, currentPlainKey_36_port, currentPlainKey_35_port
      , currentPlainKey_34_port, currentPlainKey_33_port, 
      currentPlainKey_32_port, currentPlainKey_31_port, currentPlainKey_30_port
      , currentPlainKey_29_port, currentPlainKey_28_port, 
      currentPlainKey_27_port, currentPlainKey_26_port, currentPlainKey_25_port
      , currentPlainKey_24_port, currentPlainKey_23_port, 
      currentPlainKey_22_port, currentPlainKey_21_port, currentPlainKey_20_port
      , currentPlainKey_19_port, currentPlainKey_18_port, 
      currentPlainKey_17_port, currentPlainKey_16_port, currentPlainKey_15_port
      , currentPlainKey_14_port, currentPlainKey_13_port, 
      currentPlainKey_12_port, currentPlainKey_11_port, currentPlainKey_10_port
      , currentPlainKey_9_port, currentPlainKey_8_port, currentPlainKey_7_port,
      currentPlainKey_6_port, currentPlainKey_5_port, currentPlainKey_4_port, 
      currentPlainKey_3_port, currentPlainKey_2_port, currentPlainKey_1_port, 
      currentPlainKey_0_port, parityAccumulator_7_port, 
      parityAccumulator_6_port, parityAccumulator_5_port, 
      parityAccumulator_4_port, parityAccumulator_3_port, 
      parityAccumulator_2_port, parityAccumulator_1_port, 
      parityAccumulator_0_port, nextParityError, N1792, N1793, N1794, N1795, 
      N1796, N1797, N1798, N1799, n3, n12, n13, n15, n18, n22, n24, n26, n28, 
      n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58
      , n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, n80, n82, n84, n86, 
      n88, n90, n92, n94, n96, n98, n100, n102, n104, n106, n108, n110, n112, 
      n114, n116, n118, n120, n122, n124, n126, n128, n130, n132, n134, n136, 
      n138, n140, n142, n144, n146, n148, n1178, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n14
      , n16, n17, n19, n20, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, 
      n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63, n65, n67, n69
      , n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95, n97, 
      n99, n101, n103, n105, n107, n109, n111, n113, n115, n117, n119, n121, 
      n123, n125, n127, n129, n131, n133, n135, n137, n139, n141, n143, n145, 
      n147, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1267, n1268, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
      n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
      n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
      n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
      n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, 
      n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
      n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, 
      n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
      n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
      n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
      n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n_1028 : std_logic;

begin
   PLAINKEY <= ( PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port, 
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port );
   CLR_RBUFF <= CLR_RBUFF_port;
   
   n3 <= '0';
   keyCount_reg_0_inst : DFFPOSX1 port map( D => n1356, CLK => CLK, Q => 
                           keyCount_0_port);
   keyCount_reg_2_inst : DFFPOSX1 port map( D => n1349, CLK => CLK, Q => 
                           keyCount_2_port);
   keyCount_reg_3_inst : DFFPOSX1 port map( D => n1355, CLK => CLK, Q => 
                           keyCount_3_port);
   state_reg_0_inst : DFFSR port map( D => n1353, CLK => CLK, R => n252, S => 
                           n1266, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => n1351, CLK => CLK, R => n252, S => 
                           n1265, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => n1352, CLK => CLK, R => n253, S => 
                           n1264, Q => state_2_port);
   state_reg_3_inst : DFFSR port map( D => n1354, CLK => CLK, R => n252, S => 
                           n1263, Q => state_3_port);
   parityAccumulator_reg_0_inst : DFFPOSX1 port map( D => n1348, CLK => CLK, Q 
                           => parityAccumulator_0_port);
   parityAccumulator_reg_1_inst : DFFPOSX1 port map( D => n1347, CLK => CLK, Q 
                           => parityAccumulator_1_port);
   parityAccumulator_reg_2_inst : DFFPOSX1 port map( D => n1346, CLK => CLK, Q 
                           => parityAccumulator_2_port);
   parityAccumulator_reg_3_inst : DFFPOSX1 port map( D => n1345, CLK => CLK, Q 
                           => parityAccumulator_3_port);
   parityAccumulator_reg_4_inst : DFFPOSX1 port map( D => n1344, CLK => CLK, Q 
                           => parityAccumulator_4_port);
   parityAccumulator_reg_5_inst : DFFPOSX1 port map( D => n1343, CLK => CLK, Q 
                           => parityAccumulator_5_port);
   parityAccumulator_reg_6_inst : DFFPOSX1 port map( D => n1342, CLK => CLK, Q 
                           => parityAccumulator_6_port);
   parityAccumulator_reg_7_inst : DFFPOSX1 port map( D => n1341, CLK => CLK, Q 
                           => parityAccumulator_7_port);
   keyCount_reg_1_inst : DFFPOSX1 port map( D => n1350, CLK => CLK, Q => 
                           keyCount_1_port);
   PARITY_ERROR_reg : DFFSR port map( D => nextParityError, CLK => CLK, R => 
                           n253, S => n1262, Q => PARITY_ERROR);
   parityError_reg : DFFSR port map( D => nextParityError, CLK => CLK, R => 
                           n253, S => n1261, Q => parityError);
   address_reg_7_inst : DFFPOSX1 port map( D => n1340, CLK => CLK, Q => 
                           address_7_port);
   address_reg_6_inst : DFFPOSX1 port map( D => n1339, CLK => CLK, Q => 
                           address_6_port);
   address_reg_5_inst : DFFPOSX1 port map( D => n1338, CLK => CLK, Q => 
                           address_5_port);
   address_reg_4_inst : DFFPOSX1 port map( D => n1337, CLK => CLK, Q => 
                           address_4_port);
   address_reg_3_inst : DFFPOSX1 port map( D => n1336, CLK => CLK, Q => 
                           address_3_port);
   address_reg_2_inst : DFFPOSX1 port map( D => n1335, CLK => CLK, Q => 
                           address_2_port);
   address_reg_1_inst : DFFPOSX1 port map( D => n1334, CLK => CLK, Q => 
                           address_1_port);
   address_reg_0_inst : DFFPOSX1 port map( D => n1333, CLK => CLK, Q => 
                           address_0_port);
   currentPlainKey_reg_63_inst : DFFPOSX1 port map( D => n1269, CLK => CLK, Q 
                           => currentPlainKey_63_port);
   currentPlainKey_reg_62_inst : DFFPOSX1 port map( D => n1270, CLK => CLK, Q 
                           => currentPlainKey_62_port);
   currentPlainKey_reg_61_inst : DFFPOSX1 port map( D => n1271, CLK => CLK, Q 
                           => currentPlainKey_61_port);
   currentPlainKey_reg_60_inst : DFFPOSX1 port map( D => n1272, CLK => CLK, Q 
                           => currentPlainKey_60_port);
   currentPlainKey_reg_59_inst : DFFPOSX1 port map( D => n1273, CLK => CLK, Q 
                           => currentPlainKey_59_port);
   currentPlainKey_reg_58_inst : DFFPOSX1 port map( D => n1274, CLK => CLK, Q 
                           => currentPlainKey_58_port);
   currentPlainKey_reg_57_inst : DFFPOSX1 port map( D => n1275, CLK => CLK, Q 
                           => currentPlainKey_57_port);
   currentPlainKey_reg_56_inst : DFFPOSX1 port map( D => n1276, CLK => CLK, Q 
                           => currentPlainKey_56_port);
   currentPlainKey_reg_55_inst : DFFPOSX1 port map( D => n1277, CLK => CLK, Q 
                           => currentPlainKey_55_port);
   currentPlainKey_reg_54_inst : DFFPOSX1 port map( D => n1278, CLK => CLK, Q 
                           => currentPlainKey_54_port);
   currentPlainKey_reg_53_inst : DFFPOSX1 port map( D => n1279, CLK => CLK, Q 
                           => currentPlainKey_53_port);
   currentPlainKey_reg_52_inst : DFFPOSX1 port map( D => n1280, CLK => CLK, Q 
                           => currentPlainKey_52_port);
   currentPlainKey_reg_51_inst : DFFPOSX1 port map( D => n1281, CLK => CLK, Q 
                           => currentPlainKey_51_port);
   currentPlainKey_reg_50_inst : DFFPOSX1 port map( D => n1282, CLK => CLK, Q 
                           => currentPlainKey_50_port);
   currentPlainKey_reg_49_inst : DFFPOSX1 port map( D => n1283, CLK => CLK, Q 
                           => currentPlainKey_49_port);
   currentPlainKey_reg_48_inst : DFFPOSX1 port map( D => n1284, CLK => CLK, Q 
                           => currentPlainKey_48_port);
   currentPlainKey_reg_47_inst : DFFPOSX1 port map( D => n1285, CLK => CLK, Q 
                           => currentPlainKey_47_port);
   currentPlainKey_reg_46_inst : DFFPOSX1 port map( D => n1286, CLK => CLK, Q 
                           => currentPlainKey_46_port);
   currentPlainKey_reg_45_inst : DFFPOSX1 port map( D => n1287, CLK => CLK, Q 
                           => currentPlainKey_45_port);
   currentPlainKey_reg_44_inst : DFFPOSX1 port map( D => n1288, CLK => CLK, Q 
                           => currentPlainKey_44_port);
   currentPlainKey_reg_43_inst : DFFPOSX1 port map( D => n1289, CLK => CLK, Q 
                           => currentPlainKey_43_port);
   currentPlainKey_reg_42_inst : DFFPOSX1 port map( D => n1290, CLK => CLK, Q 
                           => currentPlainKey_42_port);
   currentPlainKey_reg_41_inst : DFFPOSX1 port map( D => n1291, CLK => CLK, Q 
                           => currentPlainKey_41_port);
   currentPlainKey_reg_40_inst : DFFPOSX1 port map( D => n1292, CLK => CLK, Q 
                           => currentPlainKey_40_port);
   currentPlainKey_reg_39_inst : DFFPOSX1 port map( D => n1293, CLK => CLK, Q 
                           => currentPlainKey_39_port);
   currentPlainKey_reg_38_inst : DFFPOSX1 port map( D => n1294, CLK => CLK, Q 
                           => currentPlainKey_38_port);
   currentPlainKey_reg_37_inst : DFFPOSX1 port map( D => n1295, CLK => CLK, Q 
                           => currentPlainKey_37_port);
   currentPlainKey_reg_36_inst : DFFPOSX1 port map( D => n1296, CLK => CLK, Q 
                           => currentPlainKey_36_port);
   currentPlainKey_reg_35_inst : DFFPOSX1 port map( D => n1297, CLK => CLK, Q 
                           => currentPlainKey_35_port);
   currentPlainKey_reg_34_inst : DFFPOSX1 port map( D => n1298, CLK => CLK, Q 
                           => currentPlainKey_34_port);
   currentPlainKey_reg_33_inst : DFFPOSX1 port map( D => n1299, CLK => CLK, Q 
                           => currentPlainKey_33_port);
   currentPlainKey_reg_32_inst : DFFPOSX1 port map( D => n1300, CLK => CLK, Q 
                           => currentPlainKey_32_port);
   currentPlainKey_reg_31_inst : DFFPOSX1 port map( D => n1301, CLK => CLK, Q 
                           => currentPlainKey_31_port);
   currentPlainKey_reg_30_inst : DFFPOSX1 port map( D => n1302, CLK => CLK, Q 
                           => currentPlainKey_30_port);
   currentPlainKey_reg_29_inst : DFFPOSX1 port map( D => n1303, CLK => CLK, Q 
                           => currentPlainKey_29_port);
   currentPlainKey_reg_28_inst : DFFPOSX1 port map( D => n1304, CLK => CLK, Q 
                           => currentPlainKey_28_port);
   currentPlainKey_reg_27_inst : DFFPOSX1 port map( D => n1305, CLK => CLK, Q 
                           => currentPlainKey_27_port);
   currentPlainKey_reg_26_inst : DFFPOSX1 port map( D => n1306, CLK => CLK, Q 
                           => currentPlainKey_26_port);
   currentPlainKey_reg_25_inst : DFFPOSX1 port map( D => n1307, CLK => CLK, Q 
                           => currentPlainKey_25_port);
   currentPlainKey_reg_24_inst : DFFPOSX1 port map( D => n1308, CLK => CLK, Q 
                           => currentPlainKey_24_port);
   currentPlainKey_reg_23_inst : DFFPOSX1 port map( D => n1309, CLK => CLK, Q 
                           => currentPlainKey_23_port);
   currentPlainKey_reg_22_inst : DFFPOSX1 port map( D => n1310, CLK => CLK, Q 
                           => currentPlainKey_22_port);
   currentPlainKey_reg_21_inst : DFFPOSX1 port map( D => n1311, CLK => CLK, Q 
                           => currentPlainKey_21_port);
   currentPlainKey_reg_20_inst : DFFPOSX1 port map( D => n1312, CLK => CLK, Q 
                           => currentPlainKey_20_port);
   currentPlainKey_reg_19_inst : DFFPOSX1 port map( D => n1313, CLK => CLK, Q 
                           => currentPlainKey_19_port);
   currentPlainKey_reg_18_inst : DFFPOSX1 port map( D => n1314, CLK => CLK, Q 
                           => currentPlainKey_18_port);
   currentPlainKey_reg_17_inst : DFFPOSX1 port map( D => n1315, CLK => CLK, Q 
                           => currentPlainKey_17_port);
   currentPlainKey_reg_16_inst : DFFPOSX1 port map( D => n1316, CLK => CLK, Q 
                           => currentPlainKey_16_port);
   currentPlainKey_reg_15_inst : DFFPOSX1 port map( D => n1317, CLK => CLK, Q 
                           => currentPlainKey_15_port);
   currentPlainKey_reg_14_inst : DFFPOSX1 port map( D => n1318, CLK => CLK, Q 
                           => currentPlainKey_14_port);
   currentPlainKey_reg_13_inst : DFFPOSX1 port map( D => n1319, CLK => CLK, Q 
                           => currentPlainKey_13_port);
   currentPlainKey_reg_12_inst : DFFPOSX1 port map( D => n1320, CLK => CLK, Q 
                           => currentPlainKey_12_port);
   currentPlainKey_reg_11_inst : DFFPOSX1 port map( D => n1321, CLK => CLK, Q 
                           => currentPlainKey_11_port);
   currentPlainKey_reg_10_inst : DFFPOSX1 port map( D => n1322, CLK => CLK, Q 
                           => currentPlainKey_10_port);
   currentPlainKey_reg_9_inst : DFFPOSX1 port map( D => n1323, CLK => CLK, Q =>
                           currentPlainKey_9_port);
   currentPlainKey_reg_8_inst : DFFPOSX1 port map( D => n1324, CLK => CLK, Q =>
                           currentPlainKey_8_port);
   currentPlainKey_reg_7_inst : DFFPOSX1 port map( D => n1325, CLK => CLK, Q =>
                           currentPlainKey_7_port);
   currentPlainKey_reg_6_inst : DFFPOSX1 port map( D => n1326, CLK => CLK, Q =>
                           currentPlainKey_6_port);
   currentPlainKey_reg_5_inst : DFFPOSX1 port map( D => n1327, CLK => CLK, Q =>
                           currentPlainKey_5_port);
   currentPlainKey_reg_4_inst : DFFPOSX1 port map( D => n1328, CLK => CLK, Q =>
                           currentPlainKey_4_port);
   currentPlainKey_reg_3_inst : DFFPOSX1 port map( D => n1329, CLK => CLK, Q =>
                           currentPlainKey_3_port);
   currentPlainKey_reg_2_inst : DFFPOSX1 port map( D => n1330, CLK => CLK, Q =>
                           currentPlainKey_2_port);
   currentPlainKey_reg_1_inst : DFFPOSX1 port map( D => n1331, CLK => CLK, Q =>
                           currentPlainKey_1_port);
   currentPlainKey_reg_0_inst : DFFPOSX1 port map( D => n1332, CLK => CLK, Q =>
                           currentPlainKey_0_port);
   PLAINKEY_reg_63_inst : DFFPOSX1 port map( D => n1260, CLK => CLK, Q => 
                           PLAINKEY_63_port);
   PLAINKEY_reg_62_inst : DFFPOSX1 port map( D => n1259, CLK => CLK, Q => 
                           PLAINKEY_62_port);
   PLAINKEY_reg_61_inst : DFFPOSX1 port map( D => n1258, CLK => CLK, Q => 
                           PLAINKEY_61_port);
   PLAINKEY_reg_60_inst : DFFPOSX1 port map( D => n1257, CLK => CLK, Q => 
                           PLAINKEY_60_port);
   PLAINKEY_reg_59_inst : DFFPOSX1 port map( D => n1256, CLK => CLK, Q => 
                           PLAINKEY_59_port);
   PLAINKEY_reg_58_inst : DFFPOSX1 port map( D => n1255, CLK => CLK, Q => 
                           PLAINKEY_58_port);
   PLAINKEY_reg_57_inst : DFFPOSX1 port map( D => n1254, CLK => CLK, Q => 
                           PLAINKEY_57_port);
   PLAINKEY_reg_56_inst : DFFPOSX1 port map( D => n1253, CLK => CLK, Q => 
                           PLAINKEY_56_port);
   PLAINKEY_reg_55_inst : DFFPOSX1 port map( D => n1252, CLK => CLK, Q => 
                           PLAINKEY_55_port);
   PLAINKEY_reg_54_inst : DFFPOSX1 port map( D => n1251, CLK => CLK, Q => 
                           PLAINKEY_54_port);
   PLAINKEY_reg_53_inst : DFFPOSX1 port map( D => n1250, CLK => CLK, Q => 
                           PLAINKEY_53_port);
   PLAINKEY_reg_52_inst : DFFPOSX1 port map( D => n1249, CLK => CLK, Q => 
                           PLAINKEY_52_port);
   PLAINKEY_reg_51_inst : DFFPOSX1 port map( D => n1248, CLK => CLK, Q => 
                           PLAINKEY_51_port);
   PLAINKEY_reg_50_inst : DFFPOSX1 port map( D => n1247, CLK => CLK, Q => 
                           PLAINKEY_50_port);
   PLAINKEY_reg_49_inst : DFFPOSX1 port map( D => n1246, CLK => CLK, Q => 
                           PLAINKEY_49_port);
   PLAINKEY_reg_48_inst : DFFPOSX1 port map( D => n1245, CLK => CLK, Q => 
                           PLAINKEY_48_port);
   PLAINKEY_reg_47_inst : DFFPOSX1 port map( D => n1244, CLK => CLK, Q => 
                           PLAINKEY_47_port);
   PLAINKEY_reg_46_inst : DFFPOSX1 port map( D => n1243, CLK => CLK, Q => 
                           PLAINKEY_46_port);
   PLAINKEY_reg_45_inst : DFFPOSX1 port map( D => n1242, CLK => CLK, Q => 
                           PLAINKEY_45_port);
   PLAINKEY_reg_44_inst : DFFPOSX1 port map( D => n1241, CLK => CLK, Q => 
                           PLAINKEY_44_port);
   PLAINKEY_reg_43_inst : DFFPOSX1 port map( D => n1240, CLK => CLK, Q => 
                           PLAINKEY_43_port);
   PLAINKEY_reg_42_inst : DFFPOSX1 port map( D => n1239, CLK => CLK, Q => 
                           PLAINKEY_42_port);
   PLAINKEY_reg_41_inst : DFFPOSX1 port map( D => n1238, CLK => CLK, Q => 
                           PLAINKEY_41_port);
   PLAINKEY_reg_40_inst : DFFPOSX1 port map( D => n1237, CLK => CLK, Q => 
                           PLAINKEY_40_port);
   PLAINKEY_reg_39_inst : DFFPOSX1 port map( D => n1236, CLK => CLK, Q => 
                           PLAINKEY_39_port);
   PLAINKEY_reg_38_inst : DFFPOSX1 port map( D => n1235, CLK => CLK, Q => 
                           PLAINKEY_38_port);
   PLAINKEY_reg_37_inst : DFFPOSX1 port map( D => n1234, CLK => CLK, Q => 
                           PLAINKEY_37_port);
   PLAINKEY_reg_36_inst : DFFPOSX1 port map( D => n1233, CLK => CLK, Q => 
                           PLAINKEY_36_port);
   PLAINKEY_reg_35_inst : DFFPOSX1 port map( D => n1232, CLK => CLK, Q => 
                           PLAINKEY_35_port);
   PLAINKEY_reg_34_inst : DFFPOSX1 port map( D => n1231, CLK => CLK, Q => 
                           PLAINKEY_34_port);
   PLAINKEY_reg_33_inst : DFFPOSX1 port map( D => n1230, CLK => CLK, Q => 
                           PLAINKEY_33_port);
   PLAINKEY_reg_32_inst : DFFPOSX1 port map( D => n1229, CLK => CLK, Q => 
                           PLAINKEY_32_port);
   PLAINKEY_reg_31_inst : DFFPOSX1 port map( D => n1228, CLK => CLK, Q => 
                           PLAINKEY_31_port);
   PLAINKEY_reg_30_inst : DFFPOSX1 port map( D => n1227, CLK => CLK, Q => 
                           PLAINKEY_30_port);
   PLAINKEY_reg_29_inst : DFFPOSX1 port map( D => n1226, CLK => CLK, Q => 
                           PLAINKEY_29_port);
   PLAINKEY_reg_28_inst : DFFPOSX1 port map( D => n1225, CLK => CLK, Q => 
                           PLAINKEY_28_port);
   PLAINKEY_reg_27_inst : DFFPOSX1 port map( D => n1224, CLK => CLK, Q => 
                           PLAINKEY_27_port);
   PLAINKEY_reg_26_inst : DFFPOSX1 port map( D => n1223, CLK => CLK, Q => 
                           PLAINKEY_26_port);
   PLAINKEY_reg_25_inst : DFFPOSX1 port map( D => n1222, CLK => CLK, Q => 
                           PLAINKEY_25_port);
   PLAINKEY_reg_24_inst : DFFPOSX1 port map( D => n1221, CLK => CLK, Q => 
                           PLAINKEY_24_port);
   PLAINKEY_reg_23_inst : DFFPOSX1 port map( D => n1220, CLK => CLK, Q => 
                           PLAINKEY_23_port);
   PLAINKEY_reg_22_inst : DFFPOSX1 port map( D => n1219, CLK => CLK, Q => 
                           PLAINKEY_22_port);
   PLAINKEY_reg_21_inst : DFFPOSX1 port map( D => n1218, CLK => CLK, Q => 
                           PLAINKEY_21_port);
   PLAINKEY_reg_20_inst : DFFPOSX1 port map( D => n1217, CLK => CLK, Q => 
                           PLAINKEY_20_port);
   PLAINKEY_reg_19_inst : DFFPOSX1 port map( D => n1216, CLK => CLK, Q => 
                           PLAINKEY_19_port);
   PLAINKEY_reg_18_inst : DFFPOSX1 port map( D => n1215, CLK => CLK, Q => 
                           PLAINKEY_18_port);
   PLAINKEY_reg_17_inst : DFFPOSX1 port map( D => n1214, CLK => CLK, Q => 
                           PLAINKEY_17_port);
   PLAINKEY_reg_16_inst : DFFPOSX1 port map( D => n1213, CLK => CLK, Q => 
                           PLAINKEY_16_port);
   PLAINKEY_reg_15_inst : DFFPOSX1 port map( D => n1212, CLK => CLK, Q => 
                           PLAINKEY_15_port);
   PLAINKEY_reg_14_inst : DFFPOSX1 port map( D => n1211, CLK => CLK, Q => 
                           PLAINKEY_14_port);
   PLAINKEY_reg_13_inst : DFFPOSX1 port map( D => n1210, CLK => CLK, Q => 
                           PLAINKEY_13_port);
   PLAINKEY_reg_12_inst : DFFPOSX1 port map( D => n1209, CLK => CLK, Q => 
                           PLAINKEY_12_port);
   PLAINKEY_reg_11_inst : DFFPOSX1 port map( D => n1208, CLK => CLK, Q => 
                           PLAINKEY_11_port);
   PLAINKEY_reg_10_inst : DFFPOSX1 port map( D => n1207, CLK => CLK, Q => 
                           PLAINKEY_10_port);
   PLAINKEY_reg_9_inst : DFFPOSX1 port map( D => n1206, CLK => CLK, Q => 
                           PLAINKEY_9_port);
   PLAINKEY_reg_8_inst : DFFPOSX1 port map( D => n1205, CLK => CLK, Q => 
                           PLAINKEY_8_port);
   PLAINKEY_reg_7_inst : DFFPOSX1 port map( D => n1204, CLK => CLK, Q => 
                           PLAINKEY_7_port);
   PLAINKEY_reg_6_inst : DFFPOSX1 port map( D => n1203, CLK => CLK, Q => 
                           PLAINKEY_6_port);
   PLAINKEY_reg_5_inst : DFFPOSX1 port map( D => n1202, CLK => CLK, Q => 
                           PLAINKEY_5_port);
   PLAINKEY_reg_4_inst : DFFPOSX1 port map( D => n1201, CLK => CLK, Q => 
                           PLAINKEY_4_port);
   PLAINKEY_reg_3_inst : DFFPOSX1 port map( D => n1200, CLK => CLK, Q => 
                           PLAINKEY_3_port);
   PLAINKEY_reg_2_inst : DFFPOSX1 port map( D => n1199, CLK => CLK, Q => 
                           PLAINKEY_2_port);
   PLAINKEY_reg_1_inst : DFFPOSX1 port map( D => n1198, CLK => CLK, Q => 
                           PLAINKEY_1_port);
   PLAINKEY_reg_0_inst : DFFPOSX1 port map( D => n1197, CLK => CLK, Q => 
                           PLAINKEY_0_port);
   U9 : NAND3X1 port map( A => parityAccumulator_7_port, B => 
                           parityAccumulator_6_port, C => n15, Y => n13);
   U10 : NOR2X1 port map( A => n1627, B => n1628, Y => n15);
   U11 : NAND3X1 port map( A => parityAccumulator_3_port, B => 
                           parityAccumulator_2_port, C => n18, Y => n12);
   U12 : NOR2X1 port map( A => n1623, B => n1624, Y => n18);
   U13 : OAI21X1 port map( A => n239, B => n1694, C => n22, Y => n1197);
   U14 : NAND2X1 port map( A => PLAINKEY_0_port, B => n244, Y => n22);
   U15 : OAI21X1 port map( A => n239, B => n1693, C => n24, Y => n1198);
   U16 : NAND2X1 port map( A => PLAINKEY_1_port, B => n247, Y => n24);
   U17 : OAI21X1 port map( A => n239, B => n1692, C => n26, Y => n1199);
   U18 : NAND2X1 port map( A => PLAINKEY_2_port, B => n247, Y => n26);
   U19 : OAI21X1 port map( A => n239, B => n1691, C => n28, Y => n1200);
   U20 : NAND2X1 port map( A => PLAINKEY_3_port, B => n247, Y => n28);
   U21 : OAI21X1 port map( A => n239, B => n1690, C => n30, Y => n1201);
   U22 : NAND2X1 port map( A => PLAINKEY_4_port, B => n247, Y => n30);
   U24 : OAI21X1 port map( A => n239, B => n1689, C => n32, Y => n1202);
   U25 : NAND2X1 port map( A => PLAINKEY_5_port, B => n247, Y => n32);
   U27 : OAI21X1 port map( A => n239, B => n1688, C => n34, Y => n1203);
   U28 : NAND2X1 port map( A => PLAINKEY_6_port, B => n247, Y => n34);
   U30 : OAI21X1 port map( A => n239, B => n1687, C => n36, Y => n1204);
   U31 : NAND2X1 port map( A => PLAINKEY_7_port, B => n247, Y => n36);
   U33 : OAI21X1 port map( A => n239, B => n1686, C => n38, Y => n1205);
   U34 : NAND2X1 port map( A => PLAINKEY_8_port, B => n247, Y => n38);
   U36 : OAI21X1 port map( A => n240, B => n1685, C => n40, Y => n1206);
   U37 : NAND2X1 port map( A => PLAINKEY_9_port, B => n247, Y => n40);
   U39 : OAI21X1 port map( A => n240, B => n1684, C => n42, Y => n1207);
   U40 : NAND2X1 port map( A => PLAINKEY_10_port, B => n247, Y => n42);
   U42 : OAI21X1 port map( A => n240, B => n1683, C => n44, Y => n1208);
   U43 : NAND2X1 port map( A => PLAINKEY_11_port, B => n246, Y => n44);
   U45 : OAI21X1 port map( A => n240, B => n1682, C => n46, Y => n1209);
   U46 : NAND2X1 port map( A => PLAINKEY_12_port, B => n246, Y => n46);
   U48 : OAI21X1 port map( A => n240, B => n1681, C => n48, Y => n1210);
   U49 : NAND2X1 port map( A => PLAINKEY_13_port, B => n246, Y => n48);
   U51 : OAI21X1 port map( A => n240, B => n1680, C => n50, Y => n1211);
   U52 : NAND2X1 port map( A => PLAINKEY_14_port, B => n246, Y => n50);
   U54 : OAI21X1 port map( A => n240, B => n1679, C => n52, Y => n1212);
   U55 : NAND2X1 port map( A => PLAINKEY_15_port, B => n246, Y => n52);
   U57 : OAI21X1 port map( A => n241, B => n1678, C => n54, Y => n1213);
   U58 : NAND2X1 port map( A => PLAINKEY_16_port, B => n246, Y => n54);
   U60 : OAI21X1 port map( A => n241, B => n1677, C => n56, Y => n1214);
   U61 : NAND2X1 port map( A => PLAINKEY_17_port, B => n246, Y => n56);
   U63 : OAI21X1 port map( A => n241, B => n1676, C => n58, Y => n1215);
   U64 : NAND2X1 port map( A => PLAINKEY_18_port, B => n246, Y => n58);
   U66 : OAI21X1 port map( A => n241, B => n1675, C => n60, Y => n1216);
   U67 : NAND2X1 port map( A => PLAINKEY_19_port, B => n246, Y => n60);
   U69 : OAI21X1 port map( A => n241, B => n1674, C => n62, Y => n1217);
   U70 : NAND2X1 port map( A => PLAINKEY_20_port, B => n246, Y => n62);
   U72 : OAI21X1 port map( A => n241, B => n1673, C => n64, Y => n1218);
   U73 : NAND2X1 port map( A => PLAINKEY_21_port, B => n246, Y => n64);
   U75 : OAI21X1 port map( A => n241, B => n1672, C => n66, Y => n1219);
   U76 : NAND2X1 port map( A => PLAINKEY_22_port, B => n246, Y => n66);
   U78 : OAI21X1 port map( A => n242, B => n1671, C => n68, Y => n1220);
   U79 : NAND2X1 port map( A => PLAINKEY_23_port, B => n246, Y => n68);
   U81 : OAI21X1 port map( A => n241, B => n1670, C => n70, Y => n1221);
   U82 : NAND2X1 port map( A => PLAINKEY_24_port, B => n246, Y => n70);
   U84 : OAI21X1 port map( A => n240, B => n1669, C => n72, Y => n1222);
   U85 : NAND2X1 port map( A => PLAINKEY_25_port, B => n246, Y => n72);
   U87 : OAI21X1 port map( A => n242, B => n1668, C => n74, Y => n1223);
   U88 : NAND2X1 port map( A => PLAINKEY_26_port, B => n246, Y => n74);
   U90 : OAI21X1 port map( A => n242, B => n1667, C => n76, Y => n1224);
   U91 : NAND2X1 port map( A => PLAINKEY_27_port, B => n246, Y => n76);
   U93 : OAI21X1 port map( A => n241, B => n1666, C => n78, Y => n1225);
   U94 : NAND2X1 port map( A => PLAINKEY_28_port, B => n246, Y => n78);
   U96 : OAI21X1 port map( A => n242, B => n1665, C => n80, Y => n1226);
   U97 : NAND2X1 port map( A => PLAINKEY_29_port, B => n245, Y => n80);
   U99 : OAI21X1 port map( A => n242, B => n1664, C => n82, Y => n1227);
   U100 : NAND2X1 port map( A => PLAINKEY_30_port, B => n245, Y => n82);
   U102 : OAI21X1 port map( A => n243, B => n1663, C => n84, Y => n1228);
   U103 : NAND2X1 port map( A => PLAINKEY_31_port, B => n245, Y => n84);
   U105 : OAI21X1 port map( A => n243, B => n1662, C => n86, Y => n1229);
   U106 : NAND2X1 port map( A => PLAINKEY_32_port, B => n245, Y => n86);
   U108 : OAI21X1 port map( A => n242, B => n1661, C => n88, Y => n1230);
   U109 : NAND2X1 port map( A => PLAINKEY_33_port, B => n245, Y => n88);
   U111 : OAI21X1 port map( A => n243, B => n1660, C => n90, Y => n1231);
   U112 : NAND2X1 port map( A => PLAINKEY_34_port, B => n245, Y => n90);
   U114 : OAI21X1 port map( A => n242, B => n1659, C => n92, Y => n1232);
   U115 : NAND2X1 port map( A => PLAINKEY_35_port, B => n245, Y => n92);
   U117 : OAI21X1 port map( A => n242, B => n1658, C => n94, Y => n1233);
   U118 : NAND2X1 port map( A => PLAINKEY_36_port, B => n245, Y => n94);
   U120 : OAI21X1 port map( A => n243, B => n1657, C => n96, Y => n1234);
   U121 : NAND2X1 port map( A => PLAINKEY_37_port, B => n245, Y => n96);
   U123 : OAI21X1 port map( A => n243, B => n1656, C => n98, Y => n1235);
   U124 : NAND2X1 port map( A => PLAINKEY_38_port, B => n245, Y => n98);
   U126 : OAI21X1 port map( A => n243, B => n1655, C => n100, Y => n1236);
   U127 : NAND2X1 port map( A => PLAINKEY_39_port, B => n245, Y => n100);
   U129 : OAI21X1 port map( A => n243, B => n1654, C => n102, Y => n1237);
   U130 : NAND2X1 port map( A => PLAINKEY_40_port, B => n245, Y => n102);
   U132 : OAI21X1 port map( A => n243, B => n1653, C => n104, Y => n1238);
   U133 : NAND2X1 port map( A => PLAINKEY_41_port, B => n245, Y => n104);
   U135 : OAI21X1 port map( A => n242, B => n1652, C => n106, Y => n1239);
   U136 : NAND2X1 port map( A => PLAINKEY_42_port, B => n245, Y => n106);
   U138 : OAI21X1 port map( A => n243, B => n1651, C => n108, Y => n1240);
   U139 : NAND2X1 port map( A => PLAINKEY_43_port, B => n245, Y => n108);
   U141 : OAI21X1 port map( A => n243, B => n1650, C => n110, Y => n1241);
   U142 : NAND2X1 port map( A => PLAINKEY_44_port, B => n244, Y => n110);
   U144 : OAI21X1 port map( A => n243, B => n1649, C => n112, Y => n1242);
   U145 : NAND2X1 port map( A => PLAINKEY_45_port, B => n244, Y => n112);
   U147 : OAI21X1 port map( A => n243, B => n1648, C => n114, Y => n1243);
   U148 : NAND2X1 port map( A => PLAINKEY_46_port, B => n245, Y => n114);
   U150 : OAI21X1 port map( A => n240, B => n1647, C => n116, Y => n1244);
   U151 : NAND2X1 port map( A => PLAINKEY_47_port, B => n244, Y => n116);
   U153 : OAI21X1 port map( A => n242, B => n1646, C => n118, Y => n1245);
   U154 : NAND2X1 port map( A => PLAINKEY_48_port, B => n244, Y => n118);
   U156 : OAI21X1 port map( A => n242, B => n1645, C => n120, Y => n1246);
   U157 : NAND2X1 port map( A => PLAINKEY_49_port, B => n244, Y => n120);
   U159 : OAI21X1 port map( A => n242, B => n1644, C => n122, Y => n1247);
   U160 : NAND2X1 port map( A => PLAINKEY_50_port, B => n244, Y => n122);
   U162 : OAI21X1 port map( A => n241, B => n1643, C => n124, Y => n1248);
   U163 : NAND2X1 port map( A => PLAINKEY_51_port, B => n244, Y => n124);
   U165 : OAI21X1 port map( A => n242, B => n1642, C => n126, Y => n1249);
   U166 : NAND2X1 port map( A => PLAINKEY_52_port, B => n244, Y => n126);
   U168 : OAI21X1 port map( A => n241, B => n1641, C => n128, Y => n1250);
   U169 : NAND2X1 port map( A => PLAINKEY_53_port, B => n244, Y => n128);
   U171 : OAI21X1 port map( A => n241, B => n1640, C => n130, Y => n1251);
   U172 : NAND2X1 port map( A => PLAINKEY_54_port, B => n244, Y => n130);
   U174 : OAI21X1 port map( A => n240, B => n1639, C => n132, Y => n1252);
   U175 : NAND2X1 port map( A => PLAINKEY_55_port, B => n245, Y => n132);
   U177 : OAI21X1 port map( A => n241, B => n1638, C => n134, Y => n1253);
   U178 : NAND2X1 port map( A => PLAINKEY_56_port, B => n244, Y => n134);
   U180 : OAI21X1 port map( A => n240, B => n1637, C => n136, Y => n1254);
   U181 : NAND2X1 port map( A => PLAINKEY_57_port, B => n244, Y => n136);
   U183 : OAI21X1 port map( A => n240, B => n1636, C => n138, Y => n1255);
   U184 : NAND2X1 port map( A => PLAINKEY_58_port, B => n244, Y => n138);
   U186 : OAI21X1 port map( A => n240, B => n1635, C => n140, Y => n1256);
   U187 : NAND2X1 port map( A => PLAINKEY_59_port, B => n244, Y => n140);
   U188 : OAI21X1 port map( A => n239, B => n1634, C => n142, Y => n1257);
   U189 : NAND2X1 port map( A => PLAINKEY_60_port, B => n244, Y => n142);
   U191 : OAI21X1 port map( A => n239, B => n1633, C => n144, Y => n1258);
   U192 : NAND2X1 port map( A => PLAINKEY_61_port, B => n244, Y => n144);
   U194 : OAI21X1 port map( A => n239, B => n1620, C => n146, Y => n1259);
   U195 : NAND2X1 port map( A => PLAINKEY_62_port, B => n244, Y => n146);
   U196 : OAI21X1 port map( A => n239, B => n1632, C => n148, Y => n1260);
   U197 : NAND2X1 port map( A => PLAINKEY_63_port, B => n245, Y => n148);
   U1305 : NAND2X1 port map( A => n1584, B => n1695, Y => n1178);
   n1261 <= '1';
   n1262 <= '1';
   n1263 <= '1';
   n1264 <= '1';
   n1265 <= '1';
   n1266 <= '1';
   r577 : keyreg_1_DW01_add_1 port map( A(7) => parityAccumulator_7_port, A(6) 
                           => parityAccumulator_6_port, A(5) => 
                           parityAccumulator_5_port, A(4) => 
                           parityAccumulator_4_port, A(3) => 
                           parityAccumulator_3_port, A(2) => 
                           parityAccumulator_2_port, A(1) => 
                           parityAccumulator_1_port, A(0) => 
                           parityAccumulator_0_port, B(7) => RCV_DATA(7), B(6) 
                           => RCV_DATA(6), B(5) => RCV_DATA(5), B(4) => 
                           RCV_DATA(4), B(3) => RCV_DATA(3), B(2) => n236, B(1)
                           => n190, B(0) => n189, CI => n3, SUM(7) => N1799, 
                           SUM(6) => N1798, SUM(5) => N1797, SUM(4) => N1796, 
                           SUM(3) => N1795, SUM(2) => N1794, SUM(1) => N1793, 
                           SUM(0) => N1792, CO => n_1028);
   U3 : INVX2 port map( A => n191, Y => n193);
   U4 : BUFX2 port map( A => n1503, Y => n211);
   U5 : INVX4 port map( A => n31, Y => n143);
   U7 : INVX2 port map( A => n835, Y => n1080);
   U8 : BUFX2 port map( A => RCV_DATA(1), Y => n190);
   U23 : INVX4 port map( A => n67, Y => n113);
   U26 : INVX2 port map( A => RCV_DATA(1), Y => n220);
   U29 : AND2X2 port map( A => n270, B => n682, Y => n1);
   U32 : INVX1 port map( A => n167, Y => n168);
   U35 : INVX1 port map( A => n163, Y => n164);
   U38 : INVX2 port map( A => n73, Y => n1118);
   U41 : INVX2 port map( A => n81, Y => n85);
   U44 : INVX2 port map( A => n169, Y => n170);
   U47 : INVX2 port map( A => n1400, Y => n169);
   U50 : AND2X2 port map( A => n1080, B => n125, Y => n2);
   U53 : INVX1 port map( A => n1130, Y => n4);
   U56 : INVX1 port map( A => n894, Y => n5);
   U59 : INVX1 port map( A => n628, Y => n6);
   U62 : INVX1 port map( A => n1573, Y => n7);
   U65 : INVX2 port map( A => n160, Y => n1573);
   U68 : BUFX2 port map( A => n1394, Y => n8);
   U71 : INVX2 port map( A => n256, Y => n9);
   U74 : BUFX4 port map( A => state_2_port, Y => n159);
   U77 : INVX2 port map( A => n397, Y => n10);
   U80 : NAND2X1 port map( A => n156, B => n150, Y => n11);
   U83 : BUFX2 port map( A => n1600, Y => n14);
   U86 : BUFX2 port map( A => n1511, Y => n16);
   U89 : OR2X2 port map( A => n139, B => n1574, Y => n17);
   U92 : OR2X1 port map( A => n139, B => n1574, Y => n1599);
   U95 : OR2X2 port map( A => n159, B => n1573, Y => n139);
   U98 : BUFX2 port map( A => n1503, Y => n19);
   U101 : BUFX2 port map( A => n1503, Y => n20);
   U104 : NAND2X1 port map( A => RCV_DATA(6), B => n223, Y => n21);
   U107 : BUFX4 port map( A => n1527, Y => n223);
   U110 : INVX2 port map( A => n378, Y => n348);
   U113 : NAND3X1 port map( A => n1553, B => n1593, C => n267, Y => n23);
   U116 : OR2X2 port map( A => n1400, B => n191, Y => n450);
   U119 : INVX4 port map( A => address_3_port, Y => n191);
   U122 : INVX2 port map( A => n1420, Y => n25);
   U125 : NOR2X1 port map( A => address_6_port, B => address_7_port, Y => n27);
   U128 : NOR2X1 port map( A => address_6_port, B => address_7_port, Y => n29);
   U131 : AND2X2 port map( A => n266, B => n1600, Y => n267);
   U134 : OR2X2 port map( A => n835, B => n192, Y => n31);
   U137 : AND2X2 port map( A => n935, B => n1007, Y => n33);
   U140 : INVX1 port map( A => n33, Y => n987);
   U143 : AND2X2 port map( A => n902, B => n975, Y => n35);
   U146 : INVX1 port map( A => n35, Y => n955);
   U149 : AND2X2 port map( A => n438, B => n510, Y => n37);
   U152 : INVX1 port map( A => n37, Y => n490);
   U155 : INVX1 port map( A => n477, Y => n496);
   U158 : AND2X2 port map( A => n372, B => n444, Y => n39);
   U161 : INVX1 port map( A => n39, Y => n424);
   U164 : AND2X1 port map( A => n1599, B => n1578, Y => n41);
   U167 : AND2X2 port map( A => n271, B => n286, Y => n43);
   U170 : INVX1 port map( A => n43, Y => n1081);
   U173 : NAND3X1 port map( A => n1553, B => n11, C => n267, Y => n45);
   U176 : INVX2 port map( A => n1548, Y => n47);
   U179 : AND2X2 port map( A => n769, B => n844, Y => n49);
   U182 : INVX1 port map( A => n49, Y => n823);
   U185 : INVX4 port map( A => n379, Y => n51);
   U190 : BUFX2 port map( A => n161, Y => n235);
   U193 : AND2X2 port map( A => n107, B => n109, Y => n53);
   U198 : AND2X2 port map( A => n111, B => n1405, Y => n55);
   U199 : INVX1 port map( A => n55, Y => n1447);
   U200 : AND2X2 port map( A => n1033, B => n1110, Y => n57);
   U201 : INVX1 port map( A => n57, Y => n1089);
   U202 : AND2X2 port map( A => n504, B => n578, Y => n59);
   U203 : INVX1 port map( A => n59, Y => n557);
   U204 : INVX2 port map( A => n1151, Y => n61);
   U205 : INVX1 port map( A => n61, Y => n63);
   U206 : INVX4 port map( A => n152, Y => n166);
   U207 : BUFX4 port map( A => n1503, Y => n213);
   U208 : INVX1 port map( A => n447, Y => n65);
   U209 : INVX4 port map( A => n69, Y => n135);
   U210 : OR2X2 port map( A => n1514, B => n192, Y => n67);
   U211 : INVX2 port map( A => n1514, Y => n1495);
   U212 : OR2X2 port map( A => n268, B => n45, Y => n69);
   U213 : INVX1 port map( A => n369, Y => n107);
   U214 : INVX1 port map( A => n1398, Y => n1399);
   U215 : INVX4 port map( A => n332, Y => n415);
   U216 : AND2X2 port map( A => n1067, B => n1145, Y => n71);
   U217 : INVX1 port map( A => n71, Y => n1124);
   U218 : AND2X2 port map( A => n189, B => n1420, Y => n73);
   U219 : INVX1 port map( A => n1371, Y => n1394);
   U220 : AND2X2 port map( A => n803, B => n876, Y => n75);
   U221 : INVX1 port map( A => n75, Y => n856);
   U222 : AND2X2 port map( A => n537, B => n610, Y => n77);
   U223 : INVX1 port map( A => n77, Y => n590);
   U224 : AND2X2 port map( A => n1365, B => n1383, Y => n79);
   U225 : INVX1 port map( A => n79, Y => n1427);
   U226 : INVX4 port map( A => n1438, Y => n1504);
   U227 : INVX4 port map( A => n372, Y => n447);
   U228 : MUX2X1 port map( B => n208, A => n1430, S => n1380, Y => n1432);
   U229 : INVX2 port map( A => state_1_port, Y => n81);
   U230 : INVX1 port map( A => n81, Y => n83);
   U231 : NAND2X1 port map( A => n306, B => n135, Y => n87);
   U232 : INVX4 port map( A => n87, Y => n162);
   U233 : INVX1 port map( A => n204, Y => n199);
   U234 : OR2X2 port map( A => n1545, B => n1580, Y => n1546);
   U235 : INVX2 port map( A => n1545, Y => n1542);
   U236 : INVX4 port map( A => n1116, Y => n1420);
   U237 : AND2X2 port map( A => n202, B => n348, Y => n303);
   U238 : INVX4 port map( A => n1458, Y => n1528);
   U239 : INVX1 port map( A => n17, Y => n1549);
   U240 : INVX8 port map( A => n200, Y => n198);
   U241 : AND2X2 port map( A => n154, B => address_0_port, Y => n152);
   U242 : AND2X2 port map( A => n154, B => n283, Y => n89);
   U243 : INVX2 port map( A => n89, Y => n1185);
   U244 : AND2X2 port map( A => n838, B => n908, Y => n91);
   U245 : INVX1 port map( A => n91, Y => n888);
   U246 : INVX1 port map( A => n1545, Y => n1544);
   U247 : BUFX4 port map( A => n162, Y => n103);
   U248 : INVX4 port map( A => n119, Y => n195);
   U249 : INVX4 port map( A => n119, Y => n196);
   U250 : AND2X2 port map( A => n89, B => n193, Y => n93);
   U251 : INVX2 port map( A => n93, Y => n1513);
   U252 : BUFX2 port map( A => n1608, Y => n158);
   U253 : BUFX4 port map( A => n1608, Y => n157);
   U254 : BUFX4 port map( A => n1527, Y => n222);
   U255 : BUFX4 port map( A => n1527, Y => n225);
   U256 : AND2X2 port map( A => n83, B => n159, Y => n153);
   U257 : INVX4 port map( A => n322, Y => n1503);
   U258 : INVX1 port map( A => n911, Y => n95);
   U259 : INVX1 port map( A => n85, Y => n259);
   U260 : AND2X2 port map( A => n1104, B => n1179, Y => n97);
   U261 : INVX1 port map( A => n97, Y => n1158);
   U262 : AND2X2 port map( A => n572, B => n642, Y => n99);
   U263 : INVX1 port map( A => n99, Y => n622);
   U264 : INVX1 port map( A => n364, Y => n382);
   U265 : INVX1 port map( A => n14, Y => n1587);
   U266 : OR2X2 port map( A => n370, B => n369, Y => n117);
   U267 : NAND2X1 port map( A => n147, B => n260, Y => n101);
   U268 : BUFX2 port map( A => n162, Y => n105);
   U269 : BUFX4 port map( A => n1503, Y => n212);
   U270 : AND2X1 port map( A => n41, B => n302, Y => n109);
   U271 : INVX2 port map( A => n1, Y => n165);
   U272 : AND2X1 port map( A => n151, B => n1101, Y => n141);
   U273 : INVX4 port map( A => RCV_DATA(2), Y => n238);
   U274 : INVX2 port map( A => n249, Y => n242);
   U275 : INVX2 port map( A => n249, Y => n241);
   U276 : INVX2 port map( A => n248, Y => n240);
   U277 : INVX2 port map( A => n248, Y => n239);
   U278 : INVX2 port map( A => n250, Y => n243);
   U279 : INVX2 port map( A => n251, Y => n244);
   U280 : INVX2 port map( A => n251, Y => n245);
   U281 : INVX2 port map( A => n252, Y => n246);
   U282 : INVX2 port map( A => n250, Y => n247);
   U283 : BUFX2 port map( A => n1510, Y => n219);
   U284 : AND2X2 port map( A => n1399, B => n223, Y => n111);
   U285 : BUFX2 port map( A => n255, Y => n250);
   U286 : BUFX2 port map( A => n254, Y => n251);
   U287 : BUFX2 port map( A => n255, Y => n249);
   U288 : BUFX2 port map( A => n255, Y => n248);
   U289 : BUFX2 port map( A => n254, Y => n252);
   U290 : BUFX2 port map( A => n254, Y => n253);
   U291 : INVX2 port map( A => n275, Y => n360);
   U292 : INVX2 port map( A => n117, Y => n205);
   U293 : INVX2 port map( A => n117, Y => n206);
   U294 : AND2X2 port map( A => n125, B => n1495, Y => n115);
   U295 : INVX2 port map( A => n117, Y => n207);
   U296 : INVX2 port map( A => RST, Y => n254);
   U297 : INVX2 port map( A => RST, Y => n255);
   U298 : BUFX2 port map( A => n162, Y => n209);
   U299 : BUFX2 port map( A => n162, Y => n210);
   U300 : AND2X2 port map( A => n367, B => n135, Y => n119);
   U301 : AND2X2 port map( A => n1420, B => n193, Y => n121);
   U302 : AND2X2 port map( A => n61, B => n193, Y => n123);
   U303 : AND2X2 port map( A => n167, B => n193, Y => n125);
   U304 : AND2X2 port map( A => n163, B => n193, Y => n127);
   U305 : INVX2 port map( A => RCV_DATA(1), Y => n221);
   U306 : AND2X2 port map( A => n550, B => n1101, Y => n129);
   U307 : AND2X2 port map( A => n193, B => n43, Y => n131);
   U308 : AND2X2 port map( A => n152, B => n193, Y => n133);
   U309 : INVX2 port map( A => n171, Y => n172);
   U310 : INVX2 port map( A => n171, Y => n173);
   U311 : AND2X2 port map( A => n284, B => n121, Y => n137);
   U312 : INVX2 port map( A => n141, Y => n186);
   U313 : INVX2 port map( A => n141, Y => n187);
   U314 : BUFX2 port map( A => n1503, Y => n214);
   U315 : INVX2 port map( A => n238, Y => n236);
   U316 : INVX2 port map( A => n533, Y => n171);
   U317 : AND2X2 port map( A => n816, B => n1101, Y => n145);
   U318 : AND2X2 port map( A => n159, B => n81, Y => n147);
   U319 : INVX2 port map( A => n174, Y => n175);
   U320 : INVX2 port map( A => n174, Y => n176);
   U321 : INVX2 port map( A => n180, Y => n181);
   U322 : INVX2 port map( A => n180, Y => n182);
   U323 : INVX2 port map( A => n177, Y => n178);
   U324 : INVX2 port map( A => n183, Y => n184);
   U325 : INVX2 port map( A => n177, Y => n179);
   U326 : INVX2 port map( A => n183, Y => n185);
   U327 : INVX2 port map( A => n238, Y => n237);
   U328 : NOR2X1 port map( A => n160, B => n194, Y => n149);
   U329 : AND2X2 port map( A => n194, B => n1573, Y => n150);
   U330 : INVX2 port map( A => n191, Y => n192);
   U331 : INVX2 port map( A => n1476, Y => n167);
   U332 : INVX2 port map( A => n1440, Y => n163);
   U333 : INVX2 port map( A => n665, Y => n174);
   U334 : INVX2 port map( A => n931, Y => n180);
   U335 : INVX2 port map( A => n799, Y => n177);
   U336 : INVX2 port map( A => n1063, Y => n183);
   U337 : AND2X2 port map( A => address_4_port, B => address_5_port, Y => n151)
                           ;
   U338 : INVX4 port map( A => n188, Y => n189);
   U339 : INVX2 port map( A => RCV_DATA(0), Y => n188);
   U340 : AND2X2 port map( A => address_1_port, B => address_2_port, Y => n154)
                           ;
   U341 : NOR2X1 port map( A => address_6_port, B => address_7_port, Y => n155)
                           ;
   U342 : NOR2X1 port map( A => n85, B => n159, Y => n156);
   U343 : BUFX4 port map( A => state_0_port, Y => n194);
   U344 : BUFX4 port map( A => state_3_port, Y => n160);
   U345 : INVX4 port map( A => n333, Y => n1527);
   U346 : BUFX2 port map( A => n53, Y => n204);
   U347 : BUFX2 port map( A => n53, Y => n203);
   U348 : BUFX2 port map( A => n53, Y => n201);
   U349 : AND2X2 port map( A => RCV_DATA(7), B => n223, Y => n161);
   U350 : INVX1 port map( A => n161, Y => n379);
   U351 : INVX2 port map( A => n162, Y => n1439);
   U352 : INVX1 port map( A => n1593, Y => n1548);
   U353 : MUX2X1 port map( B => n1439, A => n307, S => n275, Y => n308);
   U354 : INVX4 port map( A => n298, Y => n550);
   U355 : INVX4 port map( A => n569, Y => n816);
   U356 : INVX8 port map( A => n202, Y => n197);
   U357 : BUFX4 port map( A => n53, Y => n200);
   U358 : BUFX4 port map( A => n53, Y => n202);
   U359 : BUFX4 port map( A => n162, Y => n208);
   U360 : BUFX4 port map( A => n1510, Y => n215);
   U361 : BUFX4 port map( A => n1510, Y => n216);
   U362 : BUFX4 port map( A => n1510, Y => n217);
   U363 : BUFX4 port map( A => n1510, Y => n218);
   U364 : BUFX4 port map( A => n1527, Y => n224);
   U365 : INVX8 port map( A => n228, Y => n226);
   U366 : INVX8 port map( A => n228, Y => n227);
   U367 : BUFX4 port map( A => n1529, Y => n228);
   U368 : BUFX4 port map( A => n21, Y => n229);
   U369 : BUFX4 port map( A => n21, Y => n230);
   U370 : BUFX4 port map( A => n161, Y => n231);
   U371 : BUFX4 port map( A => n161, Y => n232);
   U372 : BUFX4 port map( A => n161, Y => n233);
   U373 : BUFX4 port map( A => n161, Y => n234);
   U374 : NOR2X1 port map( A => n160, B => n194, Y => n257);
   U375 : INVX2 port map( A => n159, Y => n256);
   U376 : NAND3X1 port map( A => n257, B => n85, C => n256, Y => n1608);
   U377 : NOR2X1 port map( A => n160, B => n259, Y => n258);
   U378 : NAND3X1 port map( A => n9, B => n194, C => n258, Y => n1578);
   U379 : NAND2X1 port map( A => n158, B => n1578, Y => CLR_RBUFF_port);
   U380 : NOR2X1 port map( A => n160, B => n194, Y => n260);
   U381 : NAND2X1 port map( A => n147, B => n260, Y => n1553);
   U382 : INVX2 port map( A => n101, Y => PROG_ERROR);
   U383 : NAND2X1 port map( A => n153, B => n260, Y => n1597);
   U384 : NAND2X1 port map( A => n1597, B => n1553, Y => n264);
   U385 : INVX2 port map( A => n194, Y => n261);
   U386 : NAND2X1 port map( A => n156, B => n261, Y => n1598);
   U387 : NOR2X1 port map( A => n160, B => n159, Y => n262);
   U388 : NAND3X1 port map( A => n85, B => n194, C => n262, Y => n1600);
   U389 : OAI21X1 port map( A => n7, B => n1598, C => n1600, Y => n263);
   U390 : NOR3X1 port map( A => n264, B => CLR_RBUFF_port, C => n263, Y => 
                           n1535);
   U391 : OR2X2 port map( A => n83, B => n194, Y => n1574);
   U392 : NAND2X1 port map( A => n150, B => n147, Y => n1605);
   U393 : INVX2 port map( A => n1605, Y => n1583);
   U394 : NAND2X1 port map( A => n156, B => n150, Y => n1593);
   U395 : AOI21X1 port map( A => n1583, B => parityError, C => n1548, Y => n265
                           );
   U396 : NAND3X1 port map( A => n1535, B => n17, C => n265, Y => KEY_ERROR);
   U397 : INVX2 port map( A => currentPlainKey_63_port, Y => n1632);
   U398 : INVX2 port map( A => currentPlainKey_62_port, Y => n1620);
   U399 : INVX2 port map( A => currentPlainKey_3_port, Y => n1691);
   U400 : INVX2 port map( A => currentPlainKey_2_port, Y => n1692);
   U401 : INVX2 port map( A => currentPlainKey_1_port, Y => n1693);
   U402 : INVX2 port map( A => currentPlainKey_0_port, Y => n1694);
   U403 : INVX2 port map( A => parityAccumulator_4_port, Y => n1627);
   U404 : INVX2 port map( A => parityAccumulator_5_port, Y => n1628);
   U405 : NAND2X1 port map( A => n1599, B => n1578, Y => n268);
   U406 : AOI21X1 port map( A => n149, B => n153, C => n243, Y => n266);
   U407 : NAND3X1 port map( A => n1593, B => n1553, C => n267, Y => n369);
   U408 : NAND2X1 port map( A => n135, B => n1605, Y => n1510);
   U409 : NAND2X1 port map( A => n219, B => currentPlainKey_0_port, Y => n292);
   U410 : NAND3X1 port map( A => address_6_port, B => address_7_port, C => n151
                           , Y => n288);
   U411 : INVX2 port map( A => n288, Y => n284);
   U412 : INVX2 port map( A => address_0_port, Y => n283);
   U413 : INVX2 port map( A => address_1_port, Y => n287);
   U414 : NAND3X1 port map( A => address_2_port, B => n283, C => n287, Y => 
                           n1151);
   U415 : NAND2X1 port map( A => n284, B => n123, Y => n269);
   U416 : INVX2 port map( A => n269, Y => n344);
   U417 : INVX2 port map( A => RCV_DATA(4), Y => n305);
   U418 : NAND2X1 port map( A => n344, B => n305, Y => n282);
   U419 : NAND2X1 port map( A => n284, B => n93, Y => n378);
   U420 : INVX2 port map( A => address_2_port, Y => n286);
   U421 : NAND3X1 port map( A => address_0_port, B => address_1_port, C => n286
                           , Y => n1440);
   U422 : NAND2X1 port map( A => n284, B => n127, Y => n294);
   U423 : NAND2X1 port map( A => n294, B => n269, Y => n296);
   U424 : AOI21X1 port map( A => n348, B => n236, C => n296, Y => n278);
   U425 : NOR2X1 port map( A => address_4_port, B => n192, Y => n270);
   U426 : INVX2 port map( A => address_5_port, Y => n682);
   U427 : INVX2 port map( A => n165, Y => n314);
   U428 : NOR2X1 port map( A => address_1_port, B => address_0_port, Y => n271)
                           ;
   U429 : NAND2X1 port map( A => n314, B => n43, Y => n272);
   U430 : NAND2X1 port map( A => n189, B => n43, Y => n1083);
   U431 : INVX2 port map( A => n1083, Y => n1378);
   U432 : AOI22X1 port map( A => n272, B => currentPlainKey_0_port, C => n314, 
                           D => n1378, Y => n274);
   U433 : NAND2X1 port map( A => n284, B => n133, Y => n331);
   U434 : NAND2X1 port map( A => n378, B => n331, Y => n364);
   U435 : INVX2 port map( A => n331, Y => n397);
   U436 : NAND2X1 port map( A => n397, B => n190, Y => n273);
   U437 : OAI21X1 port map( A => n274, B => n364, C => n273, Y => n276);
   U438 : NAND3X1 port map( A => address_0_port, B => address_2_port, C => n287
                           , Y => n1476);
   U439 : NAND2X1 port map( A => n284, B => n125, Y => n275);
   U440 : MUX2X1 port map( B => n276, A => RCV_DATA(3), S => n360, Y => n277);
   U441 : NAND2X1 port map( A => n278, B => n277, Y => n281);
   U442 : INVX2 port map( A => n294, Y => n327);
   U443 : OR2X2 port map( A => n23, B => n158, Y => n333);
   U444 : INVX2 port map( A => n158, Y => n1596);
   U445 : NAND2X1 port map( A => n1596, B => RCV_DATA(5), Y => n279);
   U446 : OR2X2 port map( A => n369, B => n279, Y => n322);
   U447 : OAI21X1 port map( A => n327, B => n333, C => n322, Y => n280);
   U448 : NAND3X1 port map( A => n282, B => n281, C => n280, Y => n285);
   U449 : NAND2X1 port map( A => RCV_DATA(6), B => n223, Y => n1529);
   U450 : NAND3X1 port map( A => address_1_port, B => n283, C => n286, Y => 
                           n1116);
   U451 : MUX2X1 port map( B => n285, A => n229, S => n137, Y => n290);
   U452 : NAND3X1 port map( A => address_0_port, B => n287, C => n286, Y => 
                           n1400);
   U453 : NOR2X1 port map( A => n450, B => n288, Y => n289);
   U454 : MUX2X1 port map( B => n290, A => n232, S => n289, Y => n291);
   U455 : NAND2X1 port map( A => n292, B => n291, Y => n1332);
   U456 : NAND2X1 port map( A => n219, B => currentPlainKey_1_port, Y => n313);
   U457 : INVX2 port map( A => RCV_DATA(6), Y => n293);
   U458 : NOR2X1 port map( A => n294, B => n293, Y => n295);
   U459 : AOI22X1 port map( A => n344, B => n214, C => n295, D => n222, Y => 
                           n310);
   U460 : INVX2 port map( A => n296, Y => n324);
   U461 : NAND2X1 port map( A => n189, B => n169, Y => n1402);
   U462 : OAI21X1 port map( A => n170, B => n165, C => currentPlainKey_1_port, 
                           Y => n297);
   U463 : OAI21X1 port map( A => n1402, B => n165, C => n297, Y => n299);
   U464 : INVX2 port map( A => address_4_port, Y => n948);
   U465 : NAND3X1 port map( A => n27, B => n948, C => n682, Y => n298);
   U466 : INVX2 port map( A => n192, Y => n1101);
   U467 : NAND2X1 port map( A => n129, B => n43, Y => n332);
   U468 : MUX2X1 port map( B => n299, A => n190, S => n415, Y => n301);
   U469 : NAND2X1 port map( A => n397, B => n236, Y => n300);
   U470 : OAI21X1 port map( A => n364, B => n301, C => n300, Y => n304);
   U471 : INVX2 port map( A => RCV_DATA(3), Y => n1520);
   U472 : NOR2X1 port map( A => n1520, B => n157, Y => n302);
   U473 : AOI21X1 port map( A => n222, B => n304, C => n303, Y => n307);
   U474 : NOR2X1 port map( A => n305, B => n157, Y => n306);
   U475 : NAND2X1 port map( A => n324, B => n308, Y => n309);
   U476 : NAND2X1 port map( A => n310, B => n309, Y => n311);
   U477 : MUX2X1 port map( B => n311, A => n234, S => n137, Y => n312);
   U478 : NAND2X1 port map( A => n312, B => n313, Y => n1331);
   U479 : NOR2X1 port map( A => n1439, B => n378, Y => n326);
   U480 : NAND2X1 port map( A => n314, B => n1420, Y => n315);
   U481 : AOI22X1 port map( A => n315, B => currentPlainKey_2_port, C => n314, 
                           D => n73, Y => n317);
   U482 : NAND2X1 port map( A => n129, B => n169, Y => n411);
   U483 : NAND2X1 port map( A => n332, B => n411, Y => n391);
   U484 : INVX2 port map( A => n411, Y => n430);
   U485 : NAND2X1 port map( A => n430, B => n190, Y => n316);
   U486 : OAI21X1 port map( A => n317, B => n391, C => n316, Y => n319);
   U487 : NOR2X1 port map( A => n238, B => n332, Y => n318);
   U488 : AOI21X1 port map( A => n319, B => n10, C => n318, Y => n320);
   U489 : OAI22X1 port map( A => n320, B => n333, C => n197, D => n10, Y => 
                           n321);
   U490 : NAND2X1 port map( A => n321, B => n378, Y => n323);
   U491 : MUX2X1 port map( B => n323, A => n322, S => n360, Y => n325);
   U492 : OAI21X1 port map( A => n326, B => n325, C => n324, Y => n330);
   U493 : NAND2X1 port map( A => n344, B => n227, Y => n329);
   U494 : AOI22X1 port map( A => n327, B => n231, C => n219, D => 
                           currentPlainKey_2_port, Y => n328);
   U495 : NAND3X1 port map( A => n330, B => n329, C => n328, Y => n1330);
   U496 : NAND2X1 port map( A => n219, B => currentPlainKey_3_port, Y => n347);
   U497 : NOR2X1 port map( A => n1439, B => n10, Y => n342);
   U498 : NAND2X1 port map( A => n189, B => n163, Y => n1135);
   U499 : OAI21X1 port map( A => n164, B => n165, C => currentPlainKey_3_port, 
                           Y => n334);
   U500 : OAI21X1 port map( A => n1135, B => n165, C => n334, Y => n335);
   U501 : NAND2X1 port map( A => n129, B => n1420, Y => n372);
   U502 : MUX2X1 port map( B => n335, A => n190, S => n447, Y => n337);
   U503 : NAND2X1 port map( A => n430, B => n237, Y => n336);
   U504 : OAI21X1 port map( A => n337, B => n391, C => n336, Y => n338);
   U505 : AOI22X1 port map( A => n415, B => n203, C => n338, D => n225, Y => 
                           n340);
   U506 : NAND2X1 port map( A => n348, B => n211, Y => n339);
   U507 : OAI21X1 port map( A => n340, B => n364, C => n339, Y => n341);
   U508 : NOR2X1 port map( A => n342, B => n341, Y => n343);
   U509 : MUX2X1 port map( B => n343, A => n229, S => n360, Y => n345);
   U510 : MUX2X1 port map( B => n345, A => n233, S => n344, Y => n346);
   U511 : NAND2X1 port map( A => n347, B => n346, Y => n1329);
   U512 : AOI22X1 port map( A => n348, B => n227, C => currentPlainKey_4_port, 
                           D => n219, Y => n363);
   U513 : NAND2X1 port map( A => n129, B => n163, Y => n444);
   U514 : NAND2X1 port map( A => n189, B => n61, Y => n1455);
   U515 : OAI21X1 port map( A => n63, B => n165, C => currentPlainKey_4_port, Y
                           => n349);
   U516 : OAI21X1 port map( A => n1455, B => n165, C => n349, Y => n351);
   U517 : NOR2X1 port map( A => n221, B => n444, Y => n350);
   U518 : AOI21X1 port map( A => n39, B => n351, C => n350, Y => n353);
   U519 : NAND2X1 port map( A => n447, B => n237, Y => n352);
   U520 : OAI21X1 port map( A => n430, B => n353, C => n352, Y => n354);
   U521 : NAND2X1 port map( A => n222, B => n354, Y => n356);
   U522 : NAND2X1 port map( A => n430, B => n201, Y => n355);
   U523 : AOI21X1 port map( A => n356, B => n355, C => n364, Y => n357);
   U524 : MUX2X1 port map( B => n357, A => n208, S => n415, Y => n359);
   U525 : NAND2X1 port map( A => n397, B => n20, Y => n358);
   U526 : NAND2X1 port map( A => n359, B => n358, Y => n361);
   U527 : MUX2X1 port map( B => n361, A => n51, S => n360, Y => n362);
   U528 : NAND2X1 port map( A => n362, B => n363, Y => n1328);
   U529 : NAND2X1 port map( A => n430, B => n210, Y => n377);
   U530 : NAND2X1 port map( A => n189, B => n167, Y => n1478);
   U531 : OAI21X1 port map( A => n168, B => n165, C => currentPlainKey_5_port, 
                           Y => n365);
   U532 : OAI21X1 port map( A => n1478, B => n165, C => n365, Y => n366);
   U533 : NAND3X1 port map( A => n39, B => n222, C => n366, Y => n368);
   U534 : NOR2X1 port map( A => n220, B => n157, Y => n367);
   U535 : NAND2X1 port map( A => n129, B => n61, Y => n405);
   U536 : INVX2 port map( A => n405, Y => n481);
   U537 : MUX2X1 port map( B => n368, A => n195, S => n481, Y => n374);
   U538 : INVX2 port map( A => n444, Y => n463);
   U539 : NAND2X1 port map( A => n1596, B => n237, Y => n370);
   U540 : NAND2X1 port map( A => n463, B => n205, Y => n371);
   U541 : OAI21X1 port map( A => n199, B => n65, C => n371, Y => n373);
   U542 : INVX2 port map( A => n391, Y => n414);
   U543 : OAI21X1 port map( A => n374, B => n373, C => n414, Y => n376);
   U544 : NAND2X1 port map( A => n415, B => n212, Y => n375);
   U545 : NAND3X1 port map( A => n377, B => n376, C => n375, Y => n381);
   U546 : NOR2X1 port map( A => n379, B => n378, Y => n380);
   U547 : AOI21X1 port map( A => n382, B => n381, C => n380, Y => n384);
   U548 : AOI22X1 port map( A => n397, B => n226, C => currentPlainKey_5_port, 
                           D => n219, Y => n383);
   U549 : NAND2X1 port map( A => n384, B => n383, Y => n1327);
   U550 : AOI22X1 port map( A => n415, B => n226, C => currentPlainKey_6_port, 
                           D => n219, Y => n400);
   U551 : NAND2X1 port map( A => n129, B => n167, Y => n477);
   U552 : NAND2X1 port map( A => n405, B => n477, Y => n457);
   U553 : INVX2 port map( A => n457, Y => n480);
   U554 : NAND2X1 port map( A => n189, B => n89, Y => n1490);
   U555 : OAI21X1 port map( A => n1185, B => n165, C => currentPlainKey_6_port,
                           Y => n385);
   U556 : OAI21X1 port map( A => n1490, B => n165, C => n385, Y => n387);
   U557 : NOR2X1 port map( A => n220, B => n477, Y => n386);
   U558 : AOI21X1 port map( A => n480, B => n387, C => n386, Y => n389);
   U559 : NAND2X1 port map( A => n481, B => n237, Y => n388);
   U560 : OAI21X1 port map( A => n463, B => n389, C => n388, Y => n390);
   U561 : NAND2X1 port map( A => n222, B => n390, Y => n393);
   U562 : NAND2X1 port map( A => n463, B => n200, Y => n392);
   U563 : AOI21X1 port map( A => n393, B => n392, C => n391, Y => n394);
   U564 : MUX2X1 port map( B => n394, A => n209, S => n447, Y => n396);
   U565 : NAND2X1 port map( A => n430, B => n214, Y => n395);
   U566 : NAND2X1 port map( A => n396, B => n395, Y => n398);
   U567 : MUX2X1 port map( B => n398, A => n234, S => n397, Y => n399);
   U568 : NAND2X1 port map( A => n400, B => n399, Y => n1326);
   U569 : NAND2X1 port map( A => n463, B => n210, Y => n410);
   U570 : NAND2X1 port map( A => n189, B => n152, Y => n1361);
   U571 : OAI21X1 port map( A => n166, B => n165, C => currentPlainKey_7_port, 
                           Y => n401);
   U572 : OAI21X1 port map( A => n1361, B => n165, C => n401, Y => n402);
   U573 : NAND3X1 port map( A => n480, B => n225, C => n402, Y => n403);
   U574 : NAND2X1 port map( A => n129, B => n89, Y => n438);
   U575 : INVX2 port map( A => n438, Y => n513);
   U576 : MUX2X1 port map( B => n403, A => n195, S => n513, Y => n407);
   U577 : NAND2X1 port map( A => n496, B => n205, Y => n404);
   U578 : OAI21X1 port map( A => n198, B => n405, C => n404, Y => n406);
   U579 : OAI21X1 port map( A => n407, B => n406, C => n39, Y => n409);
   U580 : NAND2X1 port map( A => n447, B => n20, Y => n408);
   U581 : NAND3X1 port map( A => n410, B => n409, C => n408, Y => n413);
   U582 : NOR2X1 port map( A => n230, B => n411, Y => n412);
   U583 : AOI21X1 port map( A => n414, B => n413, C => n412, Y => n417);
   U584 : AOI22X1 port map( A => n415, B => n235, C => currentPlainKey_7_port, 
                           D => n219, Y => n416);
   U585 : NAND2X1 port map( A => n417, B => n416, Y => n1325);
   U586 : AOI22X1 port map( A => n447, B => n227, C => currentPlainKey_8_port, 
                           D => n219, Y => n433);
   U587 : NAND2X1 port map( A => n129, B => n152, Y => n510);
   U588 : NAND3X1 port map( A => n192, B => n948, C => n682, Y => n533);
   U589 : OAI21X1 port map( A => n1081, B => n172, C => currentPlainKey_8_port,
                           Y => n418);
   U590 : OAI21X1 port map( A => n1083, B => n173, C => n418, Y => n420);
   U591 : NOR2X1 port map( A => n220, B => n510, Y => n419);
   U592 : AOI21X1 port map( A => n37, B => n420, C => n419, Y => n422);
   U593 : NAND2X1 port map( A => n513, B => n237, Y => n421);
   U594 : OAI21X1 port map( A => n496, B => n422, C => n421, Y => n423);
   U595 : NAND2X1 port map( A => n222, B => n423, Y => n426);
   U596 : NAND2X1 port map( A => n496, B => n201, Y => n425);
   U597 : AOI21X1 port map( A => n426, B => n425, C => n424, Y => n427);
   U598 : MUX2X1 port map( B => n427, A => n210, S => n481, Y => n429);
   U599 : NAND2X1 port map( A => n463, B => n20, Y => n428);
   U600 : NAND2X1 port map( A => n429, B => n428, Y => n431);
   U601 : MUX2X1 port map( B => n431, A => n233, S => n430, Y => n432);
   U602 : NAND2X1 port map( A => n433, B => n432, Y => n1324);
   U603 : NAND2X1 port map( A => n496, B => n105, Y => n443);
   U604 : OAI21X1 port map( A => n170, B => n172, C => currentPlainKey_9_port, 
                           Y => n434);
   U605 : OAI21X1 port map( A => n1402, B => n173, C => n434, Y => n435);
   U606 : NAND3X1 port map( A => n37, B => n224, C => n435, Y => n436);
   U607 : NAND2X1 port map( A => n550, B => n131, Y => n471);
   U608 : INVX2 port map( A => n471, Y => n547);
   U609 : MUX2X1 port map( B => n436, A => n196, S => n547, Y => n440);
   U610 : INVX2 port map( A => n510, Y => n528);
   U611 : NAND2X1 port map( A => n528, B => n205, Y => n437);
   U612 : OAI21X1 port map( A => n198, B => n438, C => n437, Y => n439);
   U613 : OAI21X1 port map( A => n440, B => n439, C => n480, Y => n442);
   U614 : NAND2X1 port map( A => n481, B => n212, Y => n441);
   U615 : NAND3X1 port map( A => n443, B => n442, C => n441, Y => n446);
   U616 : NOR2X1 port map( A => n230, B => n444, Y => n445);
   U617 : AOI21X1 port map( A => n39, B => n446, C => n445, Y => n449);
   U618 : AOI22X1 port map( A => n447, B => n235, C => currentPlainKey_9_port, 
                           D => n218, Y => n448);
   U619 : NAND2X1 port map( A => n449, B => n448, Y => n1323);
   U620 : AOI22X1 port map( A => n481, B => n227, C => currentPlainKey_10_port,
                           D => n219, Y => n466);
   U621 : INVX2 port map( A => n450, Y => n1422);
   U622 : NAND2X1 port map( A => n550, B => n1422, Y => n543);
   U623 : NAND2X1 port map( A => n471, B => n543, Y => n522);
   U624 : INVX2 port map( A => n522, Y => n546);
   U625 : OAI21X1 port map( A => n25, B => n172, C => currentPlainKey_10_port, 
                           Y => n451);
   U626 : OAI21X1 port map( A => n1118, B => n173, C => n451, Y => n453);
   U627 : NOR2X1 port map( A => n220, B => n543, Y => n452);
   U628 : AOI21X1 port map( A => n546, B => n453, C => n452, Y => n455);
   U629 : NAND2X1 port map( A => n547, B => n237, Y => n454);
   U630 : OAI21X1 port map( A => n528, B => n455, C => n454, Y => n456);
   U631 : NAND2X1 port map( A => n224, B => n456, Y => n459);
   U632 : NAND2X1 port map( A => n528, B => n200, Y => n458);
   U633 : AOI21X1 port map( A => n459, B => n458, C => n457, Y => n460);
   U634 : MUX2X1 port map( B => n460, A => n210, S => n513, Y => n462);
   U635 : NAND2X1 port map( A => n496, B => n19, Y => n461);
   U636 : NAND2X1 port map( A => n462, B => n461, Y => n464);
   U637 : MUX2X1 port map( B => n464, A => n232, S => n463, Y => n465);
   U638 : NAND2X1 port map( A => n466, B => n465, Y => n1322);
   U639 : NAND2X1 port map( A => n528, B => n209, Y => n476);
   U640 : OAI21X1 port map( A => n164, B => n172, C => currentPlainKey_11_port,
                           Y => n467);
   U641 : OAI21X1 port map( A => n1135, B => n173, C => n467, Y => n468);
   U642 : NAND3X1 port map( A => n546, B => n222, C => n468, Y => n469);
   U643 : NAND2X1 port map( A => n550, B => n121, Y => n504);
   U644 : INVX2 port map( A => n504, Y => n581);
   U645 : MUX2X1 port map( B => n469, A => n196, S => n581, Y => n473);
   U646 : INVX2 port map( A => n543, Y => n563);
   U647 : NAND2X1 port map( A => n563, B => n205, Y => n470);
   U648 : OAI21X1 port map( A => n198, B => n471, C => n470, Y => n472);
   U649 : OAI21X1 port map( A => n473, B => n472, C => n37, Y => n475);
   U650 : NAND2X1 port map( A => n513, B => n212, Y => n474);
   U651 : NAND3X1 port map( A => n476, B => n475, C => n474, Y => n479);
   U652 : NOR2X1 port map( A => n230, B => n477, Y => n478);
   U653 : AOI21X1 port map( A => n480, B => n479, C => n478, Y => n483);
   U654 : AOI22X1 port map( A => n481, B => n234, C => currentPlainKey_11_port,
                           D => n218, Y => n482);
   U655 : NAND2X1 port map( A => n483, B => n482, Y => n1321);
   U656 : AOI22X1 port map( A => n513, B => n227, C => currentPlainKey_12_port,
                           D => n218, Y => n499);
   U657 : NAND2X1 port map( A => n550, B => n127, Y => n578);
   U658 : OAI21X1 port map( A => n63, B => n172, C => currentPlainKey_12_port, 
                           Y => n484);
   U659 : OAI21X1 port map( A => n1455, B => n173, C => n484, Y => n486);
   U660 : NOR2X1 port map( A => n220, B => n578, Y => n485);
   U661 : AOI21X1 port map( A => n59, B => n486, C => n485, Y => n488);
   U662 : NAND2X1 port map( A => n581, B => n237, Y => n487);
   U663 : OAI21X1 port map( A => n563, B => n488, C => n487, Y => n489);
   U664 : NAND2X1 port map( A => n224, B => n489, Y => n492);
   U665 : NAND2X1 port map( A => n563, B => n200, Y => n491);
   U666 : AOI21X1 port map( A => n492, B => n491, C => n490, Y => n493);
   U667 : MUX2X1 port map( B => n493, A => n208, S => n547, Y => n495);
   U668 : NAND2X1 port map( A => n528, B => n19, Y => n494);
   U669 : NAND2X1 port map( A => n495, B => n494, Y => n497);
   U670 : MUX2X1 port map( B => n497, A => n51, S => n496, Y => n498);
   U671 : NAND2X1 port map( A => n499, B => n498, Y => n1320);
   U672 : NAND2X1 port map( A => n563, B => n103, Y => n509);
   U673 : OAI21X1 port map( A => n168, B => n172, C => currentPlainKey_13_port,
                           Y => n500);
   U674 : OAI21X1 port map( A => n1478, B => n173, C => n500, Y => n501);
   U675 : NAND3X1 port map( A => n59, B => n225, C => n501, Y => n502);
   U676 : NAND2X1 port map( A => n550, B => n123, Y => n537);
   U677 : INVX2 port map( A => n537, Y => n613);
   U678 : MUX2X1 port map( B => n502, A => n196, S => n613, Y => n506);
   U679 : INVX2 port map( A => n578, Y => n596);
   U680 : NAND2X1 port map( A => n596, B => n205, Y => n503);
   U681 : OAI21X1 port map( A => n198, B => n504, C => n503, Y => n505);
   U682 : OAI21X1 port map( A => n506, B => n505, C => n546, Y => n508);
   U683 : NAND2X1 port map( A => n547, B => n214, Y => n507);
   U684 : NAND3X1 port map( A => n509, B => n508, C => n507, Y => n512);
   U685 : NOR2X1 port map( A => n229, B => n510, Y => n511);
   U686 : AOI21X1 port map( A => n37, B => n512, C => n511, Y => n515);
   U687 : AOI22X1 port map( A => n513, B => n233, C => currentPlainKey_13_port,
                           D => n218, Y => n514);
   U688 : NAND2X1 port map( A => n515, B => n514, Y => n1319);
   U689 : AOI22X1 port map( A => n547, B => n227, C => currentPlainKey_14_port,
                           D => n218, Y => n531);
   U690 : NAND2X1 port map( A => n550, B => n125, Y => n610);
   U691 : OAI21X1 port map( A => n1185, B => n172, C => currentPlainKey_14_port
                           , Y => n516);
   U692 : OAI21X1 port map( A => n1490, B => n173, C => n516, Y => n518);
   U693 : NOR2X1 port map( A => n220, B => n610, Y => n517);
   U694 : AOI21X1 port map( A => n77, B => n518, C => n517, Y => n520);
   U695 : NAND2X1 port map( A => n613, B => n237, Y => n519);
   U696 : OAI21X1 port map( A => n596, B => n520, C => n519, Y => n521);
   U697 : NAND2X1 port map( A => n225, B => n521, Y => n524);
   U698 : NAND2X1 port map( A => n596, B => n201, Y => n523);
   U699 : AOI21X1 port map( A => n524, B => n523, C => n522, Y => n525);
   U700 : MUX2X1 port map( B => n525, A => n208, S => n581, Y => n527);
   U701 : NAND2X1 port map( A => n563, B => n214, Y => n526);
   U702 : NAND2X1 port map( A => n527, B => n526, Y => n529);
   U703 : MUX2X1 port map( B => n529, A => n234, S => n528, Y => n530);
   U704 : NAND2X1 port map( A => n531, B => n530, Y => n1318);
   U705 : NAND2X1 port map( A => n596, B => n209, Y => n542);
   U706 : OAI21X1 port map( A => n166, B => n172, C => currentPlainKey_15_port,
                           Y => n532);
   U707 : OAI21X1 port map( A => n1361, B => n173, C => n532, Y => n534);
   U708 : NAND3X1 port map( A => n77, B => n225, C => n534, Y => n535);
   U709 : NAND2X1 port map( A => n550, B => n93, Y => n572);
   U710 : INVX2 port map( A => n572, Y => n645);
   U711 : MUX2X1 port map( B => n535, A => n195, S => n645, Y => n539);
   U712 : INVX2 port map( A => n610, Y => n628);
   U713 : NAND2X1 port map( A => n628, B => n205, Y => n536);
   U714 : OAI21X1 port map( A => n198, B => n537, C => n536, Y => n538);
   U715 : OAI21X1 port map( A => n539, B => n538, C => n59, Y => n541);
   U716 : NAND2X1 port map( A => n581, B => n19, Y => n540);
   U717 : NAND3X1 port map( A => n542, B => n541, C => n540, Y => n545);
   U718 : NOR2X1 port map( A => n229, B => n543, Y => n544);
   U719 : AOI21X1 port map( A => n546, B => n545, C => n544, Y => n549);
   U720 : AOI22X1 port map( A => n547, B => n231, C => currentPlainKey_15_port,
                           D => n218, Y => n548);
   U721 : NAND2X1 port map( A => n549, B => n548, Y => n1317);
   U722 : AOI22X1 port map( A => n581, B => n227, C => currentPlainKey_16_port,
                           D => n218, Y => n566);
   U723 : NAND2X1 port map( A => n550, B => n133, Y => n642);
   U724 : NAND3X1 port map( A => address_4_port, B => n1101, C => n682, Y => 
                           n665);
   U725 : OAI21X1 port map( A => n1081, B => n175, C => currentPlainKey_16_port
                           , Y => n551);
   U726 : OAI21X1 port map( A => n1083, B => n176, C => n551, Y => n553);
   U727 : NOR2X1 port map( A => n220, B => n642, Y => n552);
   U728 : AOI21X1 port map( A => n99, B => n553, C => n552, Y => n555);
   U729 : NAND2X1 port map( A => n645, B => n237, Y => n554);
   U730 : OAI21X1 port map( A => n628, B => n555, C => n554, Y => n556);
   U731 : NAND2X1 port map( A => n225, B => n556, Y => n559);
   U732 : NAND2X1 port map( A => n628, B => n204, Y => n558);
   U733 : AOI21X1 port map( A => n559, B => n558, C => n557, Y => n560);
   U734 : MUX2X1 port map( B => n560, A => n105, S => n613, Y => n562);
   U735 : NAND2X1 port map( A => n596, B => n213, Y => n561);
   U736 : NAND2X1 port map( A => n562, B => n561, Y => n564);
   U737 : MUX2X1 port map( B => n564, A => n232, S => n563, Y => n565);
   U738 : NAND2X1 port map( A => n566, B => n565, Y => n1316);
   U739 : NAND2X1 port map( A => n628, B => n105, Y => n577);
   U740 : OAI21X1 port map( A => n170, B => n175, C => currentPlainKey_17_port,
                           Y => n567);
   U741 : OAI21X1 port map( A => n1402, B => n176, C => n567, Y => n568);
   U742 : NAND3X1 port map( A => n99, B => n222, C => n568, Y => n570);
   U743 : NAND3X1 port map( A => n155, B => address_4_port, C => n682, Y => 
                           n569);
   U744 : NAND2X1 port map( A => n145, B => n43, Y => n604);
   U745 : INVX2 port map( A => n604, Y => n679);
   U746 : MUX2X1 port map( B => n570, A => n196, S => n679, Y => n574);
   U747 : INVX2 port map( A => n642, Y => n660);
   U748 : NAND2X1 port map( A => n660, B => n205, Y => n571);
   U749 : OAI21X1 port map( A => n198, B => n572, C => n571, Y => n573);
   U750 : OAI21X1 port map( A => n574, B => n573, C => n77, Y => n576);
   U751 : NAND2X1 port map( A => n613, B => n20, Y => n575);
   U752 : NAND3X1 port map( A => n577, B => n576, C => n575, Y => n580);
   U753 : NOR2X1 port map( A => n229, B => n578, Y => n579);
   U754 : AOI21X1 port map( A => n59, B => n580, C => n579, Y => n583);
   U755 : AOI22X1 port map( A => n581, B => n231, C => currentPlainKey_17_port,
                           D => n218, Y => n582);
   U756 : NAND2X1 port map( A => n583, B => n582, Y => n1315);
   U757 : AOI22X1 port map( A => n613, B => n227, C => currentPlainKey_18_port,
                           D => n218, Y => n599);
   U758 : NAND2X1 port map( A => n145, B => n169, Y => n675);
   U759 : NAND2X1 port map( A => n604, B => n675, Y => n654);
   U760 : INVX2 port map( A => n654, Y => n678);
   U761 : OAI21X1 port map( A => n25, B => n175, C => currentPlainKey_18_port, 
                           Y => n584);
   U762 : OAI21X1 port map( A => n1118, B => n176, C => n584, Y => n586);
   U763 : NOR2X1 port map( A => n220, B => n675, Y => n585);
   U764 : AOI21X1 port map( A => n678, B => n586, C => n585, Y => n588);
   U765 : NAND2X1 port map( A => n679, B => n237, Y => n587);
   U766 : OAI21X1 port map( A => n660, B => n588, C => n587, Y => n589);
   U767 : NAND2X1 port map( A => n224, B => n589, Y => n592);
   U768 : NAND2X1 port map( A => n660, B => n204, Y => n591);
   U769 : AOI21X1 port map( A => n592, B => n591, C => n590, Y => n593);
   U770 : MUX2X1 port map( B => n593, A => n209, S => n645, Y => n595);
   U771 : NAND2X1 port map( A => n628, B => n213, Y => n594);
   U772 : NAND2X1 port map( A => n595, B => n594, Y => n597);
   U773 : MUX2X1 port map( B => n597, A => n51, S => n596, Y => n598);
   U774 : NAND2X1 port map( A => n599, B => n598, Y => n1314);
   U775 : NAND2X1 port map( A => n660, B => n103, Y => n609);
   U776 : OAI21X1 port map( A => n164, B => n175, C => currentPlainKey_19_port,
                           Y => n600);
   U777 : OAI21X1 port map( A => n1135, B => n176, C => n600, Y => n601);
   U778 : NAND3X1 port map( A => n678, B => n224, C => n601, Y => n602);
   U779 : NAND2X1 port map( A => n145, B => n1420, Y => n636);
   U780 : INVX2 port map( A => n636, Y => n713);
   U781 : MUX2X1 port map( B => n602, A => n195, S => n713, Y => n606);
   U782 : INVX2 port map( A => n675, Y => n695);
   U783 : NAND2X1 port map( A => n695, B => n205, Y => n603);
   U784 : OAI21X1 port map( A => n198, B => n604, C => n603, Y => n605);
   U785 : OAI21X1 port map( A => n606, B => n605, C => n99, Y => n608);
   U786 : NAND2X1 port map( A => n645, B => n213, Y => n607);
   U787 : NAND3X1 port map( A => n609, B => n608, C => n607, Y => n612);
   U788 : NOR2X1 port map( A => n230, B => n6, Y => n611);
   U789 : AOI21X1 port map( A => n77, B => n612, C => n611, Y => n615);
   U790 : AOI22X1 port map( A => n613, B => n235, C => currentPlainKey_19_port,
                           D => n218, Y => n614);
   U791 : NAND2X1 port map( A => n615, B => n614, Y => n1313);
   U792 : AOI22X1 port map( A => n645, B => n227, C => currentPlainKey_20_port,
                           D => n218, Y => n631);
   U793 : NAND2X1 port map( A => n145, B => n163, Y => n709);
   U794 : NAND2X1 port map( A => n636, B => n709, Y => n689);
   U795 : INVX2 port map( A => n689, Y => n712);
   U796 : OAI21X1 port map( A => n63, B => n175, C => currentPlainKey_20_port, 
                           Y => n616);
   U797 : OAI21X1 port map( A => n1455, B => n176, C => n616, Y => n618);
   U798 : NOR2X1 port map( A => n220, B => n709, Y => n617);
   U799 : AOI21X1 port map( A => n712, B => n618, C => n617, Y => n620);
   U800 : NAND2X1 port map( A => n713, B => n236, Y => n619);
   U801 : OAI21X1 port map( A => n695, B => n620, C => n619, Y => n621);
   U802 : NAND2X1 port map( A => n224, B => n621, Y => n624);
   U803 : NAND2X1 port map( A => n695, B => n201, Y => n623);
   U804 : AOI21X1 port map( A => n624, B => n623, C => n622, Y => n625);
   U805 : MUX2X1 port map( B => n625, A => n103, S => n679, Y => n627);
   U806 : NAND2X1 port map( A => n660, B => n19, Y => n626);
   U807 : NAND2X1 port map( A => n627, B => n626, Y => n629);
   U808 : MUX2X1 port map( B => n629, A => n234, S => n628, Y => n630);
   U809 : NAND2X1 port map( A => n631, B => n630, Y => n1312);
   U810 : NAND2X1 port map( A => n695, B => n208, Y => n641);
   U811 : OAI21X1 port map( A => n168, B => n175, C => currentPlainKey_21_port,
                           Y => n632);
   U812 : OAI21X1 port map( A => n1478, B => n176, C => n632, Y => n633);
   U813 : NAND3X1 port map( A => n712, B => n225, C => n633, Y => n634);
   U814 : NAND2X1 port map( A => n145, B => n61, Y => n669);
   U815 : INVX2 port map( A => n669, Y => n746);
   U816 : MUX2X1 port map( B => n634, A => n195, S => n746, Y => n638);
   U817 : INVX2 port map( A => n709, Y => n728);
   U818 : NAND2X1 port map( A => n728, B => n205, Y => n635);
   U819 : OAI21X1 port map( A => n198, B => n636, C => n635, Y => n637);
   U820 : OAI21X1 port map( A => n638, B => n637, C => n678, Y => n640);
   U821 : NAND2X1 port map( A => n679, B => n212, Y => n639);
   U822 : NAND3X1 port map( A => n641, B => n640, C => n639, Y => n644);
   U823 : NOR2X1 port map( A => n229, B => n642, Y => n643);
   U824 : AOI21X1 port map( A => n99, B => n644, C => n643, Y => n647);
   U825 : AOI22X1 port map( A => n645, B => n234, C => currentPlainKey_21_port,
                           D => n218, Y => n646);
   U826 : NAND2X1 port map( A => n647, B => n646, Y => n1311);
   U827 : AOI22X1 port map( A => n679, B => n227, C => currentPlainKey_22_port,
                           D => n218, Y => n663);
   U828 : NAND2X1 port map( A => n145, B => n167, Y => n742);
   U829 : NAND2X1 port map( A => n669, B => n742, Y => n722);
   U830 : INVX2 port map( A => n722, Y => n745);
   U831 : OAI21X1 port map( A => n1185, B => n175, C => currentPlainKey_22_port
                           , Y => n648);
   U832 : OAI21X1 port map( A => n1490, B => n176, C => n648, Y => n650);
   U833 : NOR2X1 port map( A => n221, B => n742, Y => n649);
   U834 : AOI21X1 port map( A => n745, B => n650, C => n649, Y => n652);
   U835 : NAND2X1 port map( A => n746, B => n236, Y => n651);
   U836 : OAI21X1 port map( A => n728, B => n652, C => n651, Y => n653);
   U837 : NAND2X1 port map( A => n224, B => n653, Y => n656);
   U838 : NAND2X1 port map( A => n728, B => n200, Y => n655);
   U839 : AOI21X1 port map( A => n656, B => n655, C => n654, Y => n657);
   U840 : MUX2X1 port map( B => n657, A => n103, S => n713, Y => n659);
   U841 : NAND2X1 port map( A => n695, B => n19, Y => n658);
   U842 : NAND2X1 port map( A => n659, B => n658, Y => n661);
   U843 : MUX2X1 port map( B => n661, A => n233, S => n660, Y => n662);
   U844 : NAND2X1 port map( A => n663, B => n662, Y => n1310);
   U845 : NAND2X1 port map( A => n728, B => n208, Y => n674);
   U846 : OAI21X1 port map( A => n166, B => n175, C => currentPlainKey_23_port,
                           Y => n664);
   U847 : OAI21X1 port map( A => n1361, B => n176, C => n664, Y => n666);
   U848 : NAND3X1 port map( A => n745, B => n225, C => n666, Y => n667);
   U849 : NAND2X1 port map( A => n145, B => n89, Y => n703);
   U850 : INVX2 port map( A => n703, Y => n779);
   U851 : MUX2X1 port map( B => n667, A => n195, S => n779, Y => n671);
   U852 : INVX2 port map( A => n742, Y => n761);
   U853 : NAND2X1 port map( A => n761, B => n205, Y => n668);
   U854 : OAI21X1 port map( A => n198, B => n669, C => n668, Y => n670);
   U855 : OAI21X1 port map( A => n671, B => n670, C => n712, Y => n673);
   U856 : NAND2X1 port map( A => n713, B => n213, Y => n672);
   U857 : NAND3X1 port map( A => n674, B => n673, C => n672, Y => n677);
   U858 : NOR2X1 port map( A => n229, B => n675, Y => n676);
   U859 : AOI21X1 port map( A => n678, B => n677, C => n676, Y => n681);
   U860 : AOI22X1 port map( A => n679, B => n233, C => currentPlainKey_23_port,
                           D => n217, Y => n680);
   U861 : NAND2X1 port map( A => n681, B => n680, Y => n1309);
   U862 : AOI22X1 port map( A => n713, B => n227, C => currentPlainKey_24_port,
                           D => n217, Y => n698);
   U863 : NAND2X1 port map( A => n145, B => n152, Y => n775);
   U864 : NAND2X1 port map( A => n703, B => n775, Y => n755);
   U865 : INVX2 port map( A => n755, Y => n778);
   U866 : NAND3X1 port map( A => n192, B => address_4_port, C => n682, Y => 
                           n799);
   U867 : OAI21X1 port map( A => n1081, B => n178, C => currentPlainKey_24_port
                           , Y => n683);
   U868 : OAI21X1 port map( A => n1083, B => n179, C => n683, Y => n685);
   U869 : NOR2X1 port map( A => n221, B => n775, Y => n684);
   U870 : AOI21X1 port map( A => n778, B => n685, C => n684, Y => n687);
   U871 : NAND2X1 port map( A => n779, B => n236, Y => n686);
   U872 : OAI21X1 port map( A => n761, B => n687, C => n686, Y => n688);
   U873 : NAND2X1 port map( A => n225, B => n688, Y => n691);
   U874 : NAND2X1 port map( A => n761, B => n203, Y => n690);
   U875 : AOI21X1 port map( A => n691, B => n690, C => n689, Y => n692);
   U876 : MUX2X1 port map( B => n692, A => n105, S => n746, Y => n694);
   U877 : NAND2X1 port map( A => n728, B => n214, Y => n693);
   U878 : NAND2X1 port map( A => n694, B => n693, Y => n696);
   U879 : MUX2X1 port map( B => n696, A => n51, S => n695, Y => n697);
   U880 : NAND2X1 port map( A => n698, B => n697, Y => n1308);
   U881 : NAND2X1 port map( A => n761, B => n208, Y => n708);
   U882 : OAI21X1 port map( A => n170, B => n178, C => currentPlainKey_25_port,
                           Y => n699);
   U883 : OAI21X1 port map( A => n1402, B => n179, C => n699, Y => n700);
   U884 : NAND3X1 port map( A => n778, B => n222, C => n700, Y => n701);
   U885 : NAND2X1 port map( A => n816, B => n131, Y => n736);
   U886 : INVX2 port map( A => n736, Y => n813);
   U887 : MUX2X1 port map( B => n701, A => n195, S => n813, Y => n705);
   U888 : INVX2 port map( A => n775, Y => n794);
   U889 : NAND2X1 port map( A => n794, B => n205, Y => n702);
   U890 : OAI21X1 port map( A => n198, B => n703, C => n702, Y => n704);
   U891 : OAI21X1 port map( A => n705, B => n704, C => n745, Y => n707);
   U892 : NAND2X1 port map( A => n746, B => n213, Y => n706);
   U893 : NAND3X1 port map( A => n708, B => n707, C => n706, Y => n711);
   U894 : NOR2X1 port map( A => n229, B => n709, Y => n710);
   U895 : AOI21X1 port map( A => n712, B => n711, C => n710, Y => n715);
   U896 : AOI22X1 port map( A => n713, B => n235, C => currentPlainKey_25_port,
                           D => n217, Y => n714);
   U897 : NAND2X1 port map( A => n715, B => n714, Y => n1307);
   U898 : AOI22X1 port map( A => n746, B => n227, C => currentPlainKey_26_port,
                           D => n217, Y => n731);
   U899 : NAND2X1 port map( A => n816, B => n1422, Y => n809);
   U900 : NAND2X1 port map( A => n736, B => n809, Y => n788);
   U901 : INVX2 port map( A => n788, Y => n812);
   U902 : OAI21X1 port map( A => n25, B => n178, C => currentPlainKey_26_port, 
                           Y => n716);
   U903 : OAI21X1 port map( A => n1118, B => n179, C => n716, Y => n718);
   U904 : NOR2X1 port map( A => n221, B => n809, Y => n717);
   U905 : AOI21X1 port map( A => n812, B => n718, C => n717, Y => n720);
   U906 : NAND2X1 port map( A => n813, B => n236, Y => n719);
   U907 : OAI21X1 port map( A => n794, B => n720, C => n719, Y => n721);
   U908 : NAND2X1 port map( A => n225, B => n721, Y => n724);
   U909 : NAND2X1 port map( A => n794, B => n204, Y => n723);
   U910 : AOI21X1 port map( A => n724, B => n723, C => n722, Y => n725);
   U911 : MUX2X1 port map( B => n725, A => n105, S => n779, Y => n727);
   U912 : NAND2X1 port map( A => n761, B => n213, Y => n726);
   U913 : NAND2X1 port map( A => n727, B => n726, Y => n729);
   U914 : MUX2X1 port map( B => n729, A => n232, S => n728, Y => n730);
   U915 : NAND2X1 port map( A => n731, B => n730, Y => n1306);
   U916 : NAND2X1 port map( A => n794, B => n208, Y => n741);
   U917 : OAI21X1 port map( A => n164, B => n178, C => currentPlainKey_27_port,
                           Y => n732);
   U918 : OAI21X1 port map( A => n1135, B => n179, C => n732, Y => n733);
   U919 : NAND3X1 port map( A => n812, B => n222, C => n733, Y => n734);
   U920 : NAND2X1 port map( A => n816, B => n121, Y => n769);
   U921 : INVX2 port map( A => n769, Y => n847);
   U922 : MUX2X1 port map( B => n734, A => n195, S => n847, Y => n738);
   U923 : INVX2 port map( A => n809, Y => n829);
   U924 : NAND2X1 port map( A => n829, B => n205, Y => n735);
   U925 : OAI21X1 port map( A => n198, B => n736, C => n735, Y => n737);
   U926 : OAI21X1 port map( A => n738, B => n737, C => n778, Y => n740);
   U927 : NAND2X1 port map( A => n779, B => n212, Y => n739);
   U928 : NAND3X1 port map( A => n741, B => n740, C => n739, Y => n744);
   U929 : NOR2X1 port map( A => n229, B => n742, Y => n743);
   U930 : AOI21X1 port map( A => n745, B => n744, C => n743, Y => n748);
   U931 : AOI22X1 port map( A => n746, B => n232, C => currentPlainKey_27_port,
                           D => n217, Y => n747);
   U932 : NAND2X1 port map( A => n748, B => n747, Y => n1305);
   U933 : AOI22X1 port map( A => n779, B => n227, C => currentPlainKey_28_port,
                           D => n217, Y => n764);
   U934 : NAND2X1 port map( A => n816, B => n127, Y => n844);
   U935 : OAI21X1 port map( A => n63, B => n178, C => currentPlainKey_28_port, 
                           Y => n749);
   U936 : OAI21X1 port map( A => n1455, B => n179, C => n749, Y => n751);
   U937 : NOR2X1 port map( A => n221, B => n844, Y => n750);
   U938 : AOI21X1 port map( A => n49, B => n751, C => n750, Y => n753);
   U939 : NAND2X1 port map( A => n847, B => n236, Y => n752);
   U940 : OAI21X1 port map( A => n829, B => n753, C => n752, Y => n754);
   U941 : NAND2X1 port map( A => n224, B => n754, Y => n757);
   U942 : NAND2X1 port map( A => n829, B => n201, Y => n756);
   U943 : AOI21X1 port map( A => n757, B => n756, C => n755, Y => n758);
   U944 : MUX2X1 port map( B => n758, A => n103, S => n813, Y => n760);
   U945 : NAND2X1 port map( A => n794, B => n20, Y => n759);
   U946 : NAND2X1 port map( A => n760, B => n759, Y => n762);
   U947 : MUX2X1 port map( B => n762, A => n234, S => n761, Y => n763);
   U948 : NAND2X1 port map( A => n764, B => n763, Y => n1304);
   U949 : NAND2X1 port map( A => n829, B => n208, Y => n774);
   U950 : OAI21X1 port map( A => n168, B => n178, C => currentPlainKey_29_port,
                           Y => n765);
   U951 : OAI21X1 port map( A => n1478, B => n179, C => n765, Y => n766);
   U952 : NAND3X1 port map( A => n49, B => n224, C => n766, Y => n767);
   U953 : NAND2X1 port map( A => n816, B => n123, Y => n803);
   U954 : INVX2 port map( A => n803, Y => n879);
   U955 : MUX2X1 port map( B => n767, A => n196, S => n879, Y => n771);
   U956 : INVX2 port map( A => n844, Y => n862);
   U957 : NAND2X1 port map( A => n862, B => n206, Y => n768);
   U958 : OAI21X1 port map( A => n198, B => n769, C => n768, Y => n770);
   U959 : OAI21X1 port map( A => n771, B => n770, C => n812, Y => n773);
   U960 : NAND2X1 port map( A => n813, B => n19, Y => n772);
   U961 : NAND3X1 port map( A => n774, B => n773, C => n772, Y => n777);
   U962 : NOR2X1 port map( A => n230, B => n775, Y => n776);
   U963 : AOI21X1 port map( A => n778, B => n777, C => n776, Y => n781);
   U964 : AOI22X1 port map( A => n779, B => n234, C => currentPlainKey_29_port,
                           D => n217, Y => n780);
   U965 : NAND2X1 port map( A => n781, B => n780, Y => n1303);
   U966 : AOI22X1 port map( A => n813, B => n227, C => currentPlainKey_30_port,
                           D => n217, Y => n797);
   U967 : NAND2X1 port map( A => n816, B => n125, Y => n876);
   U968 : OAI21X1 port map( A => n1185, B => n178, C => currentPlainKey_30_port
                           , Y => n782);
   U969 : OAI21X1 port map( A => n1490, B => n179, C => n782, Y => n784);
   U970 : NOR2X1 port map( A => n221, B => n876, Y => n783);
   U971 : AOI21X1 port map( A => n75, B => n784, C => n783, Y => n786);
   U972 : NAND2X1 port map( A => n879, B => n236, Y => n785);
   U973 : OAI21X1 port map( A => n862, B => n786, C => n785, Y => n787);
   U974 : NAND2X1 port map( A => n224, B => n787, Y => n790);
   U975 : NAND2X1 port map( A => n862, B => n200, Y => n789);
   U976 : AOI21X1 port map( A => n790, B => n789, C => n788, Y => n791);
   U977 : MUX2X1 port map( B => n791, A => n208, S => n847, Y => n793);
   U978 : NAND2X1 port map( A => n829, B => n212, Y => n792);
   U979 : NAND2X1 port map( A => n793, B => n792, Y => n795);
   U980 : MUX2X1 port map( B => n795, A => n232, S => n794, Y => n796);
   U981 : NAND2X1 port map( A => n797, B => n796, Y => n1302);
   U982 : NAND2X1 port map( A => n862, B => n210, Y => n808);
   U983 : OAI21X1 port map( A => n166, B => n178, C => currentPlainKey_31_port,
                           Y => n798);
   U984 : OAI21X1 port map( A => n1361, B => n179, C => n798, Y => n800);
   U985 : NAND3X1 port map( A => n75, B => n222, C => n800, Y => n801);
   U986 : NAND2X1 port map( A => n816, B => n93, Y => n838);
   U987 : INVX2 port map( A => n838, Y => n911);
   U988 : MUX2X1 port map( B => n801, A => n196, S => n911, Y => n805);
   U989 : INVX2 port map( A => n876, Y => n894);
   U990 : NAND2X1 port map( A => n894, B => n206, Y => n802);
   U991 : OAI21X1 port map( A => n197, B => n803, C => n802, Y => n804);
   U992 : OAI21X1 port map( A => n805, B => n804, C => n49, Y => n807);
   U993 : NAND2X1 port map( A => n847, B => n212, Y => n806);
   U994 : NAND3X1 port map( A => n808, B => n807, C => n806, Y => n811);
   U995 : NOR2X1 port map( A => n229, B => n809, Y => n810);
   U996 : AOI21X1 port map( A => n812, B => n811, C => n810, Y => n815);
   U997 : AOI22X1 port map( A => n813, B => n232, C => currentPlainKey_31_port,
                           D => n217, Y => n814);
   U998 : NAND2X1 port map( A => n815, B => n814, Y => n1301);
   U999 : AOI22X1 port map( A => n847, B => n227, C => currentPlainKey_32_port,
                           D => n217, Y => n832);
   U1000 : NAND2X1 port map( A => n816, B => n133, Y => n908);
   U1001 : NAND3X1 port map( A => address_5_port, B => n1101, C => n948, Y => 
                           n931);
   U1002 : OAI21X1 port map( A => n1081, B => n181, C => 
                           currentPlainKey_32_port, Y => n817);
   U1003 : OAI21X1 port map( A => n1083, B => n182, C => n817, Y => n819);
   U1004 : NOR2X1 port map( A => n221, B => n908, Y => n818);
   U1005 : AOI21X1 port map( A => n91, B => n819, C => n818, Y => n821);
   U1006 : NAND2X1 port map( A => n911, B => n236, Y => n820);
   U1007 : OAI21X1 port map( A => n821, B => n894, C => n820, Y => n822);
   U1008 : NAND2X1 port map( A => n225, B => n822, Y => n825);
   U1009 : NAND2X1 port map( A => n894, B => n203, Y => n824);
   U1010 : AOI21X1 port map( A => n825, B => n824, C => n823, Y => n826);
   U1011 : MUX2X1 port map( B => n826, A => n103, S => n879, Y => n828);
   U1012 : NAND2X1 port map( A => n862, B => n213, Y => n827);
   U1013 : NAND2X1 port map( A => n828, B => n827, Y => n830);
   U1014 : MUX2X1 port map( B => n830, A => n234, S => n829, Y => n831);
   U1015 : NAND2X1 port map( A => n832, B => n831, Y => n1300);
   U1016 : NAND2X1 port map( A => n894, B => n105, Y => n843);
   U1017 : OAI21X1 port map( A => n170, B => n181, C => currentPlainKey_33_port
                           , Y => n833);
   U1018 : OAI21X1 port map( A => n1402, B => n182, C => n833, Y => n834);
   U1019 : NAND3X1 port map( A => n91, B => n224, C => n834, Y => n836);
   U1020 : NAND3X1 port map( A => n29, B => address_5_port, C => n948, Y => 
                           n835);
   U1021 : NAND2X1 port map( A => n143, B => n43, Y => n870);
   U1022 : INVX2 port map( A => n870, Y => n945);
   U1023 : MUX2X1 port map( B => n836, A => n196, S => n945, Y => n840);
   U1024 : INVX2 port map( A => n908, Y => n926);
   U1025 : NAND2X1 port map( A => n926, B => n206, Y => n837);
   U1026 : OAI21X1 port map( A => n197, B => n95, C => n837, Y => n839);
   U1027 : OAI21X1 port map( A => n840, B => n839, C => n75, Y => n842);
   U1028 : NAND2X1 port map( A => n879, B => n213, Y => n841);
   U1029 : NAND3X1 port map( A => n843, B => n842, C => n841, Y => n846);
   U1030 : NOR2X1 port map( A => n230, B => n844, Y => n845);
   U1031 : AOI21X1 port map( A => n49, B => n846, C => n845, Y => n849);
   U1032 : AOI22X1 port map( A => n847, B => n233, C => currentPlainKey_33_port
                           , D => n217, Y => n848);
   U1033 : NAND2X1 port map( A => n849, B => n848, Y => n1299);
   U1034 : AOI22X1 port map( A => n879, B => n226, C => currentPlainKey_34_port
                           , D => n217, Y => n865);
   U1035 : NAND2X1 port map( A => n143, B => n169, Y => n941);
   U1036 : NAND2X1 port map( A => n870, B => n941, Y => n920);
   U1037 : INVX2 port map( A => n920, Y => n944);
   U1038 : OAI21X1 port map( A => n25, B => n181, C => currentPlainKey_34_port,
                           Y => n850);
   U1039 : OAI21X1 port map( A => n1118, B => n182, C => n850, Y => n852);
   U1040 : NOR2X1 port map( A => n221, B => n941, Y => n851);
   U1041 : AOI21X1 port map( A => n944, B => n852, C => n851, Y => n854);
   U1042 : NAND2X1 port map( A => n945, B => n236, Y => n853);
   U1043 : OAI21X1 port map( A => n926, B => n854, C => n853, Y => n855);
   U1044 : NAND2X1 port map( A => n222, B => n855, Y => n858);
   U1045 : NAND2X1 port map( A => n926, B => n203, Y => n857);
   U1046 : AOI21X1 port map( A => n858, B => n857, C => n856, Y => n859);
   U1047 : MUX2X1 port map( B => n859, A => n105, S => n911, Y => n861);
   U1048 : NAND2X1 port map( A => n894, B => n212, Y => n860);
   U1049 : NAND2X1 port map( A => n861, B => n860, Y => n863);
   U1050 : MUX2X1 port map( B => n863, A => n233, S => n862, Y => n864);
   U1051 : NAND2X1 port map( A => n865, B => n864, Y => n1298);
   U1052 : NAND2X1 port map( A => n926, B => n105, Y => n875);
   U1053 : OAI21X1 port map( A => n164, B => n181, C => currentPlainKey_35_port
                           , Y => n866);
   U1054 : OAI21X1 port map( A => n1135, B => n182, C => n866, Y => n867);
   U1055 : NAND3X1 port map( A => n944, B => n224, C => n867, Y => n868);
   U1056 : NAND2X1 port map( A => n143, B => n1420, Y => n902);
   U1057 : INVX2 port map( A => n902, Y => n978);
   U1058 : MUX2X1 port map( B => n868, A => n195, S => n978, Y => n872);
   U1059 : INVX2 port map( A => n941, Y => n961);
   U1060 : NAND2X1 port map( A => n961, B => n206, Y => n869);
   U1061 : OAI21X1 port map( A => n197, B => n870, C => n869, Y => n871);
   U1062 : OAI21X1 port map( A => n872, B => n871, C => n91, Y => n874);
   U1063 : NAND2X1 port map( A => n911, B => n20, Y => n873);
   U1064 : NAND3X1 port map( A => n875, B => n874, C => n873, Y => n878);
   U1065 : NOR2X1 port map( A => n230, B => n5, Y => n877);
   U1066 : AOI21X1 port map( A => n75, B => n878, C => n877, Y => n881);
   U1067 : AOI22X1 port map( A => n879, B => n233, C => currentPlainKey_35_port
                           , D => n216, Y => n880);
   U1068 : NAND2X1 port map( A => n881, B => n880, Y => n1297);
   U1069 : AOI22X1 port map( A => n911, B => n226, C => currentPlainKey_36_port
                           , D => n216, Y => n897);
   U1070 : NAND2X1 port map( A => n143, B => n163, Y => n975);
   U1071 : OAI21X1 port map( A => n63, B => n181, C => currentPlainKey_36_port,
                           Y => n882);
   U1072 : OAI21X1 port map( A => n1455, B => n182, C => n882, Y => n884);
   U1073 : NOR2X1 port map( A => n221, B => n975, Y => n883);
   U1074 : AOI21X1 port map( A => n35, B => n884, C => n883, Y => n886);
   U1075 : NAND2X1 port map( A => n978, B => n236, Y => n885);
   U1076 : OAI21X1 port map( A => n961, B => n886, C => n885, Y => n887);
   U1077 : NAND2X1 port map( A => n224, B => n887, Y => n890);
   U1078 : NAND2X1 port map( A => n961, B => n200, Y => n889);
   U1079 : AOI21X1 port map( A => n890, B => n889, C => n888, Y => n891);
   U1080 : MUX2X1 port map( B => n891, A => n208, S => n945, Y => n893);
   U1081 : NAND2X1 port map( A => n926, B => n213, Y => n892);
   U1082 : NAND2X1 port map( A => n893, B => n892, Y => n895);
   U1083 : MUX2X1 port map( B => n895, A => n234, S => n894, Y => n896);
   U1084 : NAND2X1 port map( A => n897, B => n896, Y => n1296);
   U1085 : NAND2X1 port map( A => n961, B => n162, Y => n907);
   U1086 : OAI21X1 port map( A => n168, B => n181, C => currentPlainKey_37_port
                           , Y => n898);
   U1087 : OAI21X1 port map( A => n1478, B => n182, C => n898, Y => n899);
   U1088 : NAND3X1 port map( A => n35, B => n222, C => n899, Y => n900);
   U1089 : NAND2X1 port map( A => n143, B => n61, Y => n935);
   U1090 : INVX2 port map( A => n935, Y => n1010);
   U1091 : MUX2X1 port map( B => n900, A => n195, S => n1010, Y => n904);
   U1092 : INVX2 port map( A => n975, Y => n993);
   U1093 : NAND2X1 port map( A => n993, B => n206, Y => n901);
   U1094 : OAI21X1 port map( A => n197, B => n902, C => n901, Y => n903);
   U1095 : OAI21X1 port map( A => n904, B => n903, C => n944, Y => n906);
   U1096 : NAND2X1 port map( A => n945, B => n20, Y => n905);
   U1097 : NAND3X1 port map( A => n907, B => n906, C => n905, Y => n910);
   U1098 : NOR2X1 port map( A => n230, B => n908, Y => n909);
   U1099 : AOI21X1 port map( A => n91, B => n910, C => n909, Y => n913);
   U1100 : AOI22X1 port map( A => n911, B => n235, C => currentPlainKey_37_port
                           , D => n216, Y => n912);
   U1101 : NAND2X1 port map( A => n913, B => n912, Y => n1295);
   U1102 : AOI22X1 port map( A => n945, B => n226, C => currentPlainKey_38_port
                           , D => n216, Y => n929);
   U1103 : NAND2X1 port map( A => n143, B => n167, Y => n1007);
   U1104 : OAI21X1 port map( A => n1185, B => n181, C => 
                           currentPlainKey_38_port, Y => n914);
   U1105 : OAI21X1 port map( A => n1490, B => n182, C => n914, Y => n916);
   U1106 : NOR2X1 port map( A => n221, B => n1007, Y => n915);
   U1107 : AOI21X1 port map( A => n33, B => n916, C => n915, Y => n918);
   U1108 : NAND2X1 port map( A => n1010, B => n236, Y => n917);
   U1109 : OAI21X1 port map( A => n993, B => n918, C => n917, Y => n919);
   U1110 : NAND2X1 port map( A => n224, B => n919, Y => n922);
   U1111 : NAND2X1 port map( A => n993, B => n200, Y => n921);
   U1112 : AOI21X1 port map( A => n922, B => n921, C => n920, Y => n923);
   U1113 : MUX2X1 port map( B => n923, A => n210, S => n978, Y => n925);
   U1114 : NAND2X1 port map( A => n961, B => n212, Y => n924);
   U1115 : NAND2X1 port map( A => n925, B => n924, Y => n927);
   U1116 : MUX2X1 port map( B => n927, A => n232, S => n926, Y => n928);
   U1117 : NAND2X1 port map( A => n929, B => n928, Y => n1294);
   U1118 : NAND2X1 port map( A => n993, B => n208, Y => n940);
   U1119 : OAI21X1 port map( A => n166, B => n181, C => currentPlainKey_39_port
                           , Y => n930);
   U1120 : OAI21X1 port map( A => n1361, B => n182, C => n930, Y => n932);
   U1121 : NAND3X1 port map( A => n33, B => n225, C => n932, Y => n933);
   U1122 : NAND2X1 port map( A => n143, B => n89, Y => n969);
   U1123 : INVX2 port map( A => n969, Y => n1043);
   U1124 : MUX2X1 port map( B => n933, A => n195, S => n1043, Y => n937);
   U1125 : INVX2 port map( A => n1007, Y => n1025);
   U1126 : NAND2X1 port map( A => n1025, B => n206, Y => n934);
   U1127 : OAI21X1 port map( A => n197, B => n935, C => n934, Y => n936);
   U1128 : OAI21X1 port map( A => n937, B => n936, C => n35, Y => n939);
   U1129 : NAND2X1 port map( A => n978, B => n213, Y => n938);
   U1130 : NAND3X1 port map( A => n940, B => n939, C => n938, Y => n943);
   U1131 : NOR2X1 port map( A => n230, B => n941, Y => n942);
   U1132 : AOI21X1 port map( A => n944, B => n943, C => n942, Y => n947);
   U1133 : AOI22X1 port map( A => n945, B => n232, C => currentPlainKey_39_port
                           , D => n216, Y => n946);
   U1134 : NAND2X1 port map( A => n947, B => n946, Y => n1293);
   U1135 : AOI22X1 port map( A => n978, B => n226, C => currentPlainKey_40_port
                           , D => n216, Y => n964);
   U1136 : NAND2X1 port map( A => n143, B => n152, Y => n1039);
   U1137 : NAND2X1 port map( A => n969, B => n1039, Y => n1019);
   U1138 : INVX2 port map( A => n1019, Y => n1042);
   U1139 : NAND3X1 port map( A => n192, B => address_5_port, C => n948, Y => 
                           n1063);
   U1140 : OAI21X1 port map( A => n1081, B => n184, C => 
                           currentPlainKey_40_port, Y => n949);
   U1141 : OAI21X1 port map( A => n1083, B => n185, C => n949, Y => n951);
   U1142 : NOR2X1 port map( A => n221, B => n1039, Y => n950);
   U1143 : AOI21X1 port map( A => n1042, B => n951, C => n950, Y => n953);
   U1144 : NAND2X1 port map( A => n1043, B => n236, Y => n952);
   U1145 : OAI21X1 port map( A => n1025, B => n953, C => n952, Y => n954);
   U1146 : NAND2X1 port map( A => n225, B => n954, Y => n957);
   U1147 : NAND2X1 port map( A => n1025, B => n201, Y => n956);
   U1148 : AOI21X1 port map( A => n957, B => n956, C => n955, Y => n958);
   U1149 : MUX2X1 port map( B => n958, A => n209, S => n1010, Y => n960);
   U1150 : NAND2X1 port map( A => n993, B => n212, Y => n959);
   U1151 : NAND2X1 port map( A => n960, B => n959, Y => n962);
   U1152 : MUX2X1 port map( B => n962, A => n234, S => n961, Y => n963);
   U1153 : NAND2X1 port map( A => n964, B => n963, Y => n1292);
   U1154 : NAND2X1 port map( A => n1025, B => n209, Y => n974);
   U1155 : OAI21X1 port map( A => n170, B => n184, C => currentPlainKey_41_port
                           , Y => n965);
   U1156 : OAI21X1 port map( A => n1402, B => n185, C => n965, Y => n966);
   U1157 : NAND3X1 port map( A => n1042, B => n225, C => n966, Y => n967);
   U1158 : NAND2X1 port map( A => n1080, B => n131, Y => n1001);
   U1159 : INVX2 port map( A => n1001, Y => n1077);
   U1160 : MUX2X1 port map( B => n967, A => n196, S => n1077, Y => n971);
   U1161 : INVX2 port map( A => n1039, Y => n1058);
   U1162 : NAND2X1 port map( A => n1058, B => n206, Y => n968);
   U1163 : OAI21X1 port map( A => n197, B => n969, C => n968, Y => n970);
   U1164 : OAI21X1 port map( A => n971, B => n970, C => n33, Y => n973);
   U1165 : NAND2X1 port map( A => n1010, B => n212, Y => n972);
   U1166 : NAND3X1 port map( A => n974, B => n973, C => n972, Y => n977);
   U1167 : NOR2X1 port map( A => n229, B => n975, Y => n976);
   U1168 : AOI21X1 port map( A => n35, B => n977, C => n976, Y => n980);
   U1169 : AOI22X1 port map( A => n978, B => n234, C => currentPlainKey_41_port
                           , D => n216, Y => n979);
   U1170 : NAND2X1 port map( A => n980, B => n979, Y => n1291);
   U1171 : AOI22X1 port map( A => n1010, B => n226, C => 
                           currentPlainKey_42_port, D => n216, Y => n996);
   U1172 : NAND2X1 port map( A => n1080, B => n1422, Y => n1073);
   U1173 : NAND2X1 port map( A => n1001, B => n1073, Y => n1052);
   U1174 : INVX2 port map( A => n1052, Y => n1076);
   U1175 : OAI21X1 port map( A => n25, B => n184, C => currentPlainKey_42_port,
                           Y => n981);
   U1176 : OAI21X1 port map( A => n1118, B => n185, C => n981, Y => n983);
   U1177 : NOR2X1 port map( A => n221, B => n1073, Y => n982);
   U1178 : AOI21X1 port map( A => n1076, B => n983, C => n982, Y => n985);
   U1179 : NAND2X1 port map( A => n1077, B => n236, Y => n984);
   U1180 : OAI21X1 port map( A => n1058, B => n985, C => n984, Y => n986);
   U1181 : NAND2X1 port map( A => n222, B => n986, Y => n989);
   U1182 : NAND2X1 port map( A => n1058, B => n202, Y => n988);
   U1183 : AOI21X1 port map( A => n989, B => n988, C => n987, Y => n990);
   U1184 : MUX2X1 port map( B => n990, A => n208, S => n1043, Y => n992);
   U1185 : NAND2X1 port map( A => n1025, B => n212, Y => n991);
   U1186 : NAND2X1 port map( A => n992, B => n991, Y => n994);
   U1187 : MUX2X1 port map( B => n994, A => n51, S => n993, Y => n995);
   U1188 : NAND2X1 port map( A => n996, B => n995, Y => n1290);
   U1189 : NAND2X1 port map( A => n1058, B => n210, Y => n1006);
   U1190 : OAI21X1 port map( A => n164, B => n184, C => currentPlainKey_43_port
                           , Y => n997);
   U1191 : OAI21X1 port map( A => n1135, B => n185, C => n997, Y => n998);
   U1192 : NAND3X1 port map( A => n1076, B => n225, C => n998, Y => n999);
   U1193 : NAND2X1 port map( A => n1080, B => n121, Y => n1033);
   U1194 : INVX2 port map( A => n1033, Y => n1113);
   U1195 : MUX2X1 port map( B => n999, A => n195, S => n1113, Y => n1003);
   U1196 : INVX2 port map( A => n1073, Y => n1095);
   U1197 : NAND2X1 port map( A => n1095, B => n206, Y => n1000);
   U1198 : OAI21X1 port map( A => n198, B => n1001, C => n1000, Y => n1002);
   U1199 : OAI21X1 port map( A => n1003, B => n1002, C => n1042, Y => n1005);
   U1200 : NAND2X1 port map( A => n1043, B => n212, Y => n1004);
   U1201 : NAND3X1 port map( A => n1006, B => n1005, C => n1004, Y => n1009);
   U1202 : NOR2X1 port map( A => n230, B => n1007, Y => n1008);
   U1203 : AOI21X1 port map( A => n33, B => n1009, C => n1008, Y => n1012);
   U1204 : AOI22X1 port map( A => n1010, B => n234, C => 
                           currentPlainKey_43_port, D => n216, Y => n1011);
   U1205 : NAND2X1 port map( A => n1012, B => n1011, Y => n1289);
   U1206 : AOI22X1 port map( A => n1043, B => n226, C => 
                           currentPlainKey_44_port, D => n216, Y => n1028);
   U1207 : NAND2X1 port map( A => n1080, B => n127, Y => n1110);
   U1208 : OAI21X1 port map( A => n63, B => n184, C => currentPlainKey_44_port,
                           Y => n1013);
   U1209 : OAI21X1 port map( A => n1455, B => n185, C => n1013, Y => n1015);
   U1210 : NOR2X1 port map( A => n221, B => n1110, Y => n1014);
   U1211 : AOI21X1 port map( A => n57, B => n1015, C => n1014, Y => n1017);
   U1212 : NAND2X1 port map( A => n1113, B => n236, Y => n1016);
   U1213 : OAI21X1 port map( A => n1095, B => n1017, C => n1016, Y => n1018);
   U1214 : NAND2X1 port map( A => n224, B => n1018, Y => n1021);
   U1215 : NAND2X1 port map( A => n1095, B => n203, Y => n1020);
   U1216 : AOI21X1 port map( A => n1021, B => n1020, C => n1019, Y => n1022);
   U1217 : MUX2X1 port map( B => n1022, A => n208, S => n1077, Y => n1024);
   U1218 : NAND2X1 port map( A => n1058, B => n20, Y => n1023);
   U1219 : NAND2X1 port map( A => n1024, B => n1023, Y => n1026);
   U1220 : MUX2X1 port map( B => n1026, A => n233, S => n1025, Y => n1027);
   U1221 : NAND2X1 port map( A => n1028, B => n1027, Y => n1288);
   U1222 : NAND2X1 port map( A => n1095, B => n162, Y => n1038);
   U1223 : OAI21X1 port map( A => n168, B => n184, C => currentPlainKey_45_port
                           , Y => n1029);
   U1224 : OAI21X1 port map( A => n1478, B => n185, C => n1029, Y => n1030);
   U1225 : NAND3X1 port map( A => n57, B => n224, C => n1030, Y => n1031);
   U1226 : NAND2X1 port map( A => n1080, B => n123, Y => n1067);
   U1227 : INVX2 port map( A => n1067, Y => n1148);
   U1228 : MUX2X1 port map( B => n1031, A => n195, S => n1148, Y => n1035);
   U1229 : INVX2 port map( A => n1110, Y => n1130);
   U1230 : NAND2X1 port map( A => n1130, B => n206, Y => n1032);
   U1231 : OAI21X1 port map( A => n197, B => n1033, C => n1032, Y => n1034);
   U1232 : OAI21X1 port map( A => n1035, B => n1034, C => n1076, Y => n1037);
   U1233 : NAND2X1 port map( A => n1077, B => n212, Y => n1036);
   U1234 : NAND3X1 port map( A => n1038, B => n1037, C => n1036, Y => n1041);
   U1235 : NOR2X1 port map( A => n229, B => n1039, Y => n1040);
   U1236 : AOI21X1 port map( A => n1042, B => n1041, C => n1040, Y => n1045);
   U1237 : AOI22X1 port map( A => n1043, B => n232, C => 
                           currentPlainKey_45_port, D => n216, Y => n1044);
   U1238 : NAND2X1 port map( A => n1045, B => n1044, Y => n1287);
   U1239 : AOI22X1 port map( A => n1077, B => n226, C => 
                           currentPlainKey_46_port, D => n216, Y => n1061);
   U1240 : NAND2X1 port map( A => n1080, B => n125, Y => n1145);
   U1241 : OAI21X1 port map( A => n1185, B => n184, C => 
                           currentPlainKey_46_port, Y => n1046);
   U1242 : OAI21X1 port map( A => n1490, B => n185, C => n1046, Y => n1048);
   U1243 : NOR2X1 port map( A => n221, B => n1145, Y => n1047);
   U1244 : AOI21X1 port map( A => n71, B => n1048, C => n1047, Y => n1050);
   U1245 : NAND2X1 port map( A => n1148, B => n236, Y => n1049);
   U1246 : OAI21X1 port map( A => n1130, B => n1050, C => n1049, Y => n1051);
   U1247 : NAND2X1 port map( A => n225, B => n1051, Y => n1054);
   U1248 : NAND2X1 port map( A => n1130, B => n204, Y => n1053);
   U1249 : AOI21X1 port map( A => n1054, B => n1053, C => n1052, Y => n1055);
   U1250 : MUX2X1 port map( B => n1055, A => n103, S => n1113, Y => n1057);
   U1251 : NAND2X1 port map( A => n1095, B => n213, Y => n1056);
   U1252 : NAND2X1 port map( A => n1057, B => n1056, Y => n1059);
   U1253 : MUX2X1 port map( B => n1059, A => n233, S => n1058, Y => n1060);
   U1254 : NAND2X1 port map( A => n1061, B => n1060, Y => n1286);
   U1255 : NAND2X1 port map( A => n1130, B => n209, Y => n1072);
   U1256 : OAI21X1 port map( A => n166, B => n184, C => currentPlainKey_47_port
                           , Y => n1062);
   U1257 : OAI21X1 port map( A => n1361, B => n185, C => n1062, Y => n1064);
   U1258 : NAND3X1 port map( A => n71, B => n224, C => n1064, Y => n1065);
   U1259 : NAND2X1 port map( A => n1080, B => n93, Y => n1104);
   U1260 : INVX2 port map( A => n1104, Y => n1182);
   U1261 : MUX2X1 port map( B => n1065, A => n196, S => n1182, Y => n1069);
   U1262 : NAND2X1 port map( A => n2, B => n206, Y => n1066);
   U1263 : OAI21X1 port map( A => n197, B => n1067, C => n1066, Y => n1068);
   U1264 : OAI21X1 port map( A => n1069, B => n1068, C => n57, Y => n1071);
   U1265 : NAND2X1 port map( A => n1113, B => n213, Y => n1070);
   U1266 : NAND3X1 port map( A => n1072, B => n1071, C => n1070, Y => n1075);
   U1267 : NOR2X1 port map( A => n230, B => n1073, Y => n1074);
   U1268 : AOI21X1 port map( A => n1076, B => n1075, C => n1074, Y => n1079);
   U1269 : AOI22X1 port map( A => n1077, B => n235, C => 
                           currentPlainKey_47_port, D => n217, Y => n1078);
   U1270 : NAND2X1 port map( A => n1079, B => n1078, Y => n1285);
   U1271 : AOI22X1 port map( A => n1113, B => n226, C => 
                           currentPlainKey_48_port, D => n216, Y => n1098);
   U1272 : NAND2X1 port map( A => n1080, B => n133, Y => n1179);
   U1273 : OAI21X1 port map( A => n1081, B => n186, C => 
                           currentPlainKey_48_port, Y => n1082);
   U1274 : OAI21X1 port map( A => n1083, B => n187, C => n1082, Y => n1085);
   U1275 : NOR2X1 port map( A => n221, B => n1179, Y => n1084);
   U1276 : AOI21X1 port map( A => n97, B => n1085, C => n1084, Y => n1087);
   U1277 : NAND2X1 port map( A => n1182, B => n236, Y => n1086);
   U1278 : OAI21X1 port map( A => n2, B => n1087, C => n1086, Y => n1088);
   U1279 : NAND2X1 port map( A => n222, B => n1088, Y => n1091);
   U1280 : NAND2X1 port map( A => n2, B => n200, Y => n1090);
   U1281 : AOI21X1 port map( A => n1091, B => n1090, C => n1089, Y => n1092);
   U1282 : MUX2X1 port map( B => n1092, A => n210, S => n1148, Y => n1094);
   U1283 : NAND2X1 port map( A => n1130, B => n212, Y => n1093);
   U1284 : NAND2X1 port map( A => n1094, B => n1093, Y => n1096);
   U1285 : MUX2X1 port map( B => n1096, A => n232, S => n1095, Y => n1097);
   U1286 : NAND2X1 port map( A => n1098, B => n1097, Y => n1284);
   U1287 : NAND2X1 port map( A => n2, B => n208, Y => n1109);
   U1288 : OAI21X1 port map( A => n170, B => n186, C => currentPlainKey_49_port
                           , Y => n1099);
   U1289 : OAI21X1 port map( A => n1402, B => n187, C => n1099, Y => n1100);
   U1290 : NAND3X1 port map( A => n97, B => n224, C => n1100, Y => n1102);
   U1291 : NAND2X1 port map( A => n27, B => n151, Y => n1514);
   U1292 : NAND2X1 port map( A => n113, B => n43, Y => n1139);
   U1293 : INVX2 port map( A => n1139, Y => n1375);
   U1294 : MUX2X1 port map( B => n1102, A => n196, S => n1375, Y => n1106);
   U1295 : INVX2 port map( A => n1179, Y => n1268);
   U1296 : NAND2X1 port map( A => n1268, B => n206, Y => n1103);
   U1297 : OAI21X1 port map( A => n197, B => n1104, C => n1103, Y => n1105);
   U1298 : OAI21X1 port map( A => n1106, B => n1105, C => n71, Y => n1108);
   U1299 : NAND2X1 port map( A => n1148, B => n20, Y => n1107);
   U1300 : NAND3X1 port map( A => n1109, B => n1108, C => n1107, Y => n1112);
   U1301 : NOR2X1 port map( A => n229, B => n4, Y => n1111);
   U1302 : AOI21X1 port map( A => n57, B => n1112, C => n1111, Y => n1115);
   U1303 : AOI22X1 port map( A => n1113, B => n232, C => 
                           currentPlainKey_49_port, D => n215, Y => n1114);
   U1304 : NAND2X1 port map( A => n1115, B => n1114, Y => n1283);
   U1306 : AOI22X1 port map( A => n1148, B => n226, C => 
                           currentPlainKey_50_port, D => n215, Y => n1133);
   U1307 : NAND2X1 port map( A => n113, B => n169, Y => n1371);
   U1308 : NAND2X1 port map( A => n1139, B => n1371, Y => n1192);
   U1309 : INVX2 port map( A => n1192, Y => n1374);
   U1310 : OAI21X1 port map( A => n25, B => n186, C => currentPlainKey_50_port,
                           Y => n1117);
   U1311 : OAI21X1 port map( A => n1118, B => n187, C => n1117, Y => n1120);
   U1312 : NOR2X1 port map( A => n220, B => n1371, Y => n1119);
   U1313 : AOI21X1 port map( A => n1374, B => n1120, C => n1119, Y => n1122);
   U1314 : NAND2X1 port map( A => n1375, B => n236, Y => n1121);
   U1315 : OAI21X1 port map( A => n1268, B => n1122, C => n1121, Y => n1123);
   U1316 : NAND2X1 port map( A => n222, B => n1123, Y => n1126);
   U1317 : NAND2X1 port map( A => n1268, B => n204, Y => n1125);
   U1318 : AOI21X1 port map( A => n1126, B => n1125, C => n1124, Y => n1127);
   U1319 : MUX2X1 port map( B => n1127, A => n209, S => n1182, Y => n1129);
   U1320 : NAND2X1 port map( A => n2, B => n214, Y => n1128);
   U1321 : NAND2X1 port map( A => n1129, B => n1128, Y => n1131);
   U1322 : MUX2X1 port map( B => n1131, A => n51, S => n1130, Y => n1132);
   U1323 : NAND2X1 port map( A => n1133, B => n1132, Y => n1282);
   U1324 : NAND2X1 port map( A => n1268, B => n209, Y => n1144);
   U1325 : OAI21X1 port map( A => n164, B => n186, C => currentPlainKey_51_port
                           , Y => n1134);
   U1326 : OAI21X1 port map( A => n187, B => n1135, C => n1134, Y => n1136);
   U1327 : NAND3X1 port map( A => n1374, B => n222, C => n1136, Y => n1137);
   U1328 : NAND2X1 port map( A => n113, B => n1420, Y => n1172);
   U1329 : INVX2 port map( A => n1172, Y => n1416);
   U1330 : MUX2X1 port map( B => n1137, A => n196, S => n1416, Y => n1141);
   U1331 : NAND2X1 port map( A => n1394, B => n206, Y => n1138);
   U1332 : OAI21X1 port map( A => n197, B => n1139, C => n1138, Y => n1140);
   U1333 : OAI21X1 port map( A => n1141, B => n1140, C => n97, Y => n1143);
   U1334 : NAND2X1 port map( A => n1182, B => n213, Y => n1142);
   U1335 : NAND3X1 port map( A => n1144, B => n1143, C => n1142, Y => n1147);
   U1336 : NOR2X1 port map( A => n230, B => n1145, Y => n1146);
   U1337 : AOI21X1 port map( A => n71, B => n1147, C => n1146, Y => n1150);
   U1338 : AOI22X1 port map( A => n1148, B => n231, C => 
                           currentPlainKey_51_port, D => n215, Y => n1149);
   U1339 : NAND2X1 port map( A => n1150, B => n1149, Y => n1281);
   U1340 : AOI22X1 port map( A => n1182, B => n227, C => 
                           currentPlainKey_52_port, D => n215, Y => n1166);
   U1341 : NAND2X1 port map( A => n113, B => n163, Y => n1170);
   U1342 : NAND2X1 port map( A => n1172, B => n1170, Y => n1388);
   U1343 : INVX2 port map( A => n1388, Y => n1412);
   U1344 : OAI21X1 port map( A => n63, B => n187, C => currentPlainKey_52_port,
                           Y => n1152);
   U1345 : OAI21X1 port map( A => n1455, B => n186, C => n1152, Y => n1154);
   U1346 : NOR2X1 port map( A => n220, B => n1170, Y => n1153);
   U1347 : AOI21X1 port map( A => n1412, B => n1154, C => n1153, Y => n1156);
   U1348 : NAND2X1 port map( A => n1416, B => n236, Y => n1155);
   U1349 : OAI21X1 port map( A => n1394, B => n1156, C => n1155, Y => n1157);
   U1350 : NAND2X1 port map( A => n225, B => n1157, Y => n1160);
   U1351 : NAND2X1 port map( A => n1394, B => n203, Y => n1159);
   U1358 : AOI21X1 port map( A => n1160, B => n1159, C => n1158, Y => n1161);
   U1359 : MUX2X1 port map( B => n1161, A => n208, S => n1375, Y => n1163);
   U1360 : NAND2X1 port map( A => n1268, B => n19, Y => n1162);
   U1361 : NAND2X1 port map( A => n1163, B => n1162, Y => n1164);
   U1362 : MUX2X1 port map( B => n1164, A => n233, S => n2, Y => n1165);
   U1363 : NAND2X1 port map( A => n1166, B => n1165, Y => n1280);
   U1364 : NAND2X1 port map( A => n1394, B => n105, Y => n1177);
   U1365 : OAI21X1 port map( A => n168, B => n187, C => currentPlainKey_53_port
                           , Y => n1167);
   U1366 : OAI21X1 port map( A => n1478, B => n186, C => n1167, Y => n1168);
   U1367 : NAND3X1 port map( A => n1412, B => n224, C => n1168, Y => n1169);
   U1368 : NAND2X1 port map( A => n113, B => n61, Y => n1365);
   U1369 : INVX2 port map( A => n1365, Y => n1451);
   U1370 : MUX2X1 port map( B => n1169, A => n196, S => n1451, Y => n1174);
   U1371 : INVX2 port map( A => n1170, Y => n1433);
   U1372 : NAND2X1 port map( A => n1433, B => n207, Y => n1171);
   U1373 : OAI21X1 port map( A => n197, B => n1172, C => n1171, Y => n1173);
   U1374 : OAI21X1 port map( A => n1174, B => n1173, C => n1374, Y => n1176);
   U1375 : NAND2X1 port map( A => n1375, B => n213, Y => n1175);
   U1376 : NAND3X1 port map( A => n1177, B => n1176, C => n1175, Y => n1181);
   U1377 : NOR2X1 port map( A => n230, B => n1179, Y => n1180);
   U1378 : AOI21X1 port map( A => n97, B => n1181, C => n1180, Y => n1184);
   U1379 : AOI22X1 port map( A => n1182, B => n231, C => 
                           currentPlainKey_53_port, D => n215, Y => n1183);
   U1380 : NAND2X1 port map( A => n1184, B => n1183, Y => n1279);
   U1381 : AOI22X1 port map( A => n1375, B => n226, C => 
                           currentPlainKey_54_port, D => n215, Y => n1359);
   U1382 : NAND2X1 port map( A => n113, B => n167, Y => n1383);
   U1383 : OAI21X1 port map( A => n1185, B => n187, C => 
                           currentPlainKey_54_port, Y => n1186);
   U1384 : OAI21X1 port map( A => n186, B => n1490, C => n1186, Y => n1188);
   U1385 : NOR2X1 port map( A => n220, B => n1383, Y => n1187);
   U1386 : AOI21X1 port map( A => n79, B => n1188, C => n1187, Y => n1190);
   U1387 : NAND2X1 port map( A => n1451, B => n236, Y => n1189);
   U1388 : OAI21X1 port map( A => n1433, B => n1190, C => n1189, Y => n1191);
   U1389 : NAND2X1 port map( A => n222, B => n1191, Y => n1194);
   U1390 : NAND2X1 port map( A => n1433, B => n200, Y => n1193);
   U1391 : AOI21X1 port map( A => n1194, B => n1193, C => n1192, Y => n1195);
   U1392 : MUX2X1 port map( B => n1195, A => n103, S => n1416, Y => n1267);
   U1393 : NAND2X1 port map( A => n1394, B => n214, Y => n1196);
   U1394 : NAND2X1 port map( A => n1267, B => n1196, Y => n1357);
   U1395 : MUX2X1 port map( B => n1357, A => n232, S => n1268, Y => n1358);
   U1396 : NAND2X1 port map( A => n1359, B => n1358, Y => n1278);
   U1397 : NAND2X1 port map( A => n1433, B => n210, Y => n1370);
   U1398 : OAI21X1 port map( A => n166, B => n186, C => currentPlainKey_55_port
                           , Y => n1360);
   U1399 : OAI21X1 port map( A => n187, B => n1361, C => n1360, Y => n1362);
   U1400 : NAND3X1 port map( A => n79, B => n222, C => n1362, Y => n1363);
   U1401 : NAND2X1 port map( A => n113, B => n89, Y => n1380);
   U1402 : INVX2 port map( A => n1380, Y => n1486);
   U1403 : MUX2X1 port map( B => n1363, A => n196, S => n1486, Y => n1367);
   U1404 : INVX2 port map( A => n1383, Y => n1468);
   U1405 : NAND2X1 port map( A => n207, B => n1468, Y => n1364);
   U1406 : OAI21X1 port map( A => n1365, B => n197, C => n1364, Y => n1366);
   U1407 : OAI21X1 port map( A => n1367, B => n1366, C => n1412, Y => n1369);
   U1408 : NAND2X1 port map( A => n1416, B => n214, Y => n1368);
   U1409 : NAND3X1 port map( A => n1370, B => n1369, C => n1368, Y => n1373);
   U1410 : NOR2X1 port map( A => n229, B => n1371, Y => n1372);
   U1411 : AOI21X1 port map( A => n1374, B => n1373, C => n1372, Y => n1377);
   U1412 : AOI22X1 port map( A => n1375, B => n231, C => 
                           currentPlainKey_55_port, D => n215, Y => n1376);
   U1413 : NAND2X1 port map( A => n1377, B => n1376, Y => n1277);
   U1414 : AOI22X1 port map( A => n1416, B => n226, C => 
                           currentPlainKey_56_port, D => n215, Y => n1397);
   U1415 : NAND2X1 port map( A => n1486, B => n236, Y => n1386);
   U1416 : NAND2X1 port map( A => n193, B => n151, Y => n1511);
   U1417 : INVX2 port map( A => n1511, Y => n1491);
   U1418 : NAND2X1 port map( A => n1491, B => n43, Y => n1379);
   U1419 : AOI22X1 port map( A => currentPlainKey_56_port, B => n1379, C => 
                           n1378, D => n1491, Y => n1382);
   U1420 : NAND2X1 port map( A => n113, B => n152, Y => n1438);
   U1421 : NAND2X1 port map( A => n1380, B => n1438, Y => n1398);
   U1422 : NAND2X1 port map( A => n1504, B => n190, Y => n1381);
   U1423 : OAI21X1 port map( A => n1382, B => n1398, C => n1381, Y => n1384);
   U1424 : NAND2X1 port map( A => n1384, B => n1383, Y => n1385);
   U1425 : NAND2X1 port map( A => n1386, B => n1385, Y => n1387);
   U1426 : NAND2X1 port map( A => n225, B => n1387, Y => n1390);
   U1427 : NAND2X1 port map( A => n203, B => n1468, Y => n1389);
   U1428 : AOI21X1 port map( A => n1390, B => n1389, C => n1388, Y => n1391);
   U1429 : MUX2X1 port map( B => n1391, A => n103, S => n1451, Y => n1393);
   U1430 : NAND2X1 port map( A => n1433, B => n212, Y => n1392);
   U1431 : NAND2X1 port map( A => n1393, B => n1392, Y => n1395);
   U1432 : MUX2X1 port map( B => n1395, A => n51, S => n8, Y => n1396);
   U1433 : NAND2X1 port map( A => n1396, B => n1397, Y => n1276);
   U1434 : NAND2X1 port map( A => n1433, B => n226, Y => n1419);
   U1435 : NAND2X1 port map( A => n1495, B => n131, Y => n1405);
   U1436 : OAI21X1 port map( A => n170, B => n16, C => currentPlainKey_57_port,
                           Y => n1401);
   U1437 : OAI21X1 port map( A => n16, B => n1402, C => n1401, Y => n1403);
   U1438 : NAND2X1 port map( A => n55, B => n1403, Y => n1404);
   U1439 : NAND2X1 port map( A => n1468, B => n162, Y => n1409);
   U1440 : NAND2X1 port map( A => n1451, B => n211, Y => n1410);
   U1441 : NAND3X1 port map( A => n1404, B => n1409, C => n1410, Y => n1415);
   U1442 : NAND2X1 port map( A => n207, B => n1504, Y => n1408);
   U1443 : INVX2 port map( A => n1405, Y => n1531);
   U1444 : NAND2X1 port map( A => n1531, B => n111, Y => n1446);
   U1445 : INVX2 port map( A => n1446, Y => n1485);
   U1446 : NAND2X1 port map( A => n1485, B => n190, Y => n1407);
   U1447 : NAND2X1 port map( A => n201, B => n1486, Y => n1406);
   U1448 : NAND3X1 port map( A => n1408, B => n1407, C => n1406, Y => n1414);
   U1449 : NAND3X1 port map( A => n1410, B => n1409, C => n1427, Y => n1411);
   U1450 : AND2X2 port map( A => n1412, B => n1411, Y => n1413);
   U1451 : OAI21X1 port map( A => n1415, B => n1414, C => n1413, Y => n1418);
   U1452 : AOI22X1 port map( A => n1416, B => n231, C => 
                           currentPlainKey_57_port, D => n215, Y => n1417);
   U1453 : NAND3X1 port map( A => n1419, B => n1418, C => n1417, Y => n1275);
   U1454 : AOI22X1 port map( A => n1451, B => n226, C => 
                           currentPlainKey_58_port, D => n215, Y => n1436);
   U1455 : NAND2X1 port map( A => n204, B => n1504, Y => n1429);
   U1456 : NAND2X1 port map( A => n1420, B => n1491, Y => n1421);
   U1457 : AOI22X1 port map( A => currentPlainKey_58_port, B => n1421, C => n73
                           , D => n1491, Y => n1423);
   U1458 : NAND2X1 port map( A => n1422, B => n1495, Y => n1458);
   U1459 : MUX2X1 port map( B => n1423, A => n220, S => n1528, Y => n1424);
   U1460 : NAND2X1 port map( A => n1424, B => n1438, Y => n1425);
   U1461 : MUX2X1 port map( B => n1425, A => n238, S => n1531, Y => n1426);
   U1462 : NAND2X1 port map( A => n225, B => n1426, Y => n1428);
   U1463 : AOI21X1 port map( A => n1429, B => n1428, C => n1427, Y => n1430);
   U1464 : NAND2X1 port map( A => n1468, B => n213, Y => n1431);
   U1465 : NAND2X1 port map( A => n1432, B => n1431, Y => n1434);
   U1466 : MUX2X1 port map( B => n1434, A => n234, S => n1433, Y => n1435);
   U1467 : NAND2X1 port map( A => n1435, B => n1436, Y => n1274);
   U1468 : NAND2X1 port map( A => n1468, B => n226, Y => n1454);
   U1469 : NAND2X1 port map( A => n1486, B => n213, Y => n1437);
   U1470 : OAI21X1 port map( A => n1439, B => n1438, C => n1437, Y => n1450);
   U1471 : NOR2X1 port map( A => n238, B => n1458, Y => n1445);
   U1472 : NOR2X1 port map( A => n16, B => n164, Y => n1441);
   U1473 : MUX2X1 port map( B => n1635, A => n188, S => n1441, Y => n1442);
   U1474 : NAND2X1 port map( A => n1442, B => n1458, Y => n1443);
   U1475 : NAND2X1 port map( A => n121, B => n1495, Y => n1459);
   U1476 : INVX2 port map( A => n1459, Y => n1523);
   U1477 : MUX2X1 port map( B => n1443, A => n220, S => n1523, Y => n1444);
   U1478 : NOR2X1 port map( A => n1445, B => n1444, Y => n1448);
   U1479 : OAI22X1 port map( A => n1448, B => n1447, C => n1520, D => n1446, Y 
                           => n1449);
   U1480 : OAI21X1 port map( A => n1450, B => n1449, C => n79, Y => n1453);
   U1481 : AOI22X1 port map( A => n1451, B => n231, C => 
                           currentPlainKey_59_port, D => n215, Y => n1452);
   U1482 : NAND3X1 port map( A => n1454, B => n1453, C => n1452, Y => n1273);
   U1483 : AOI22X1 port map( A => n1486, B => n226, C => 
                           currentPlainKey_60_port, D => n215, Y => n1471);
   U1484 : NAND2X1 port map( A => n1531, B => n103, Y => n1467);
   U1485 : AOI22X1 port map( A => n1523, B => n236, C => n1528, D => 
                           RCV_DATA(3), Y => n1463);
   U1486 : NAND2X1 port map( A => n61, B => n1491, Y => n1457);
   U1487 : INVX2 port map( A => n1455, Y => n1456);
   U1488 : AOI22X1 port map( A => currentPlainKey_60_port, B => n1457, C => 
                           n1456, D => n1491, Y => n1460);
   U1489 : NAND2X1 port map( A => n1459, B => n1458, Y => n1472);
   U1490 : NOR2X1 port map( A => n1460, B => n1472, Y => n1461);
   U1491 : NAND2X1 port map( A => n127, B => n1495, Y => n1474);
   U1492 : INVX2 port map( A => n1474, Y => n1521);
   U1493 : MUX2X1 port map( B => n1461, A => n190, S => n1521, Y => n1462);
   U1494 : NAND2X1 port map( A => n1463, B => n1462, Y => n1464);
   U1495 : NAND2X1 port map( A => n55, B => n1464, Y => n1466);
   U1496 : NAND2X1 port map( A => n214, B => n1504, Y => n1465);
   U1497 : NAND3X1 port map( A => n1467, B => n1466, C => n1465, Y => n1469);
   U1498 : MUX2X1 port map( B => n1469, A => n233, S => n1468, Y => n1470);
   U1499 : NAND2X1 port map( A => n1471, B => n1470, Y => n1272);
   U1500 : NAND2X1 port map( A => n123, B => n1495, Y => n1518);
   U1501 : INVX2 port map( A => n1472, Y => n1473);
   U1502 : NAND3X1 port map( A => n1518, B => n1474, C => n1473, Y => n1475);
   U1503 : INVX2 port map( A => n1475, Y => n1499);
   U1504 : OAI21X1 port map( A => n16, B => n168, C => currentPlainKey_61_port,
                           Y => n1477);
   U1505 : OAI21X1 port map( A => n16, B => n1478, C => n1477, Y => n1480);
   U1506 : NOR2X1 port map( A => n220, B => n1518, Y => n1479);
   U1507 : AOI21X1 port map( A => n1499, B => n1480, C => n1479, Y => n1483);
   U1508 : NAND2X1 port map( A => n1521, B => n236, Y => n1482);
   U1509 : AOI22X1 port map( A => n1523, B => RCV_DATA(3), C => n1528, D => 
                           RCV_DATA(4), Y => n1481);
   U1510 : NAND3X1 port map( A => n1483, B => n1482, C => n1481, Y => n1484);
   U1511 : AOI22X1 port map( A => n1485, B => RCV_DATA(5), C => n55, D => n1484
                           , Y => n1489);
   U1512 : NAND2X1 port map( A => n227, B => n1504, Y => n1488);
   U1513 : AOI22X1 port map( A => n1486, B => n231, C => 
                           currentPlainKey_61_port, D => n215, Y => n1487);
   U1514 : NAND3X1 port map( A => n1489, B => n1488, C => n1487, Y => n1271);
   U1515 : AOI22X1 port map( A => n233, B => n1504, C => n219, D => 
                           currentPlainKey_62_port, Y => n1509);
   U1516 : INVX2 port map( A => n1490, Y => n1494);
   U1517 : AOI21X1 port map( A => n89, B => n1491, C => n1620, Y => n1493);
   U1518 : NAND2X1 port map( A => n16, B => n1620, Y => n1492);
   U1519 : OAI21X1 port map( A => n1494, B => n1493, C => n1492, Y => n1496);
   U1520 : MUX2X1 port map( B => n1496, A => n220, S => n115, Y => n1498);
   U1521 : NOR2X1 port map( A => n238, B => n1518, Y => n1497);
   U1522 : AOI21X1 port map( A => n1499, B => n1498, C => n1497, Y => n1501);
   U1523 : NAND2X1 port map( A => n1521, B => RCV_DATA(3), Y => n1500);
   U1524 : NAND2X1 port map( A => n1501, B => n1500, Y => n1502);
   U1525 : AOI22X1 port map( A => n225, B => n1502, C => n1523, D => n103, Y =>
                           n1506);
   U1526 : NAND2X1 port map( A => n1528, B => n19, Y => n1505);
   U1527 : AOI21X1 port map( A => n1506, B => n1505, C => n1504, Y => n1507);
   U1528 : MUX2X1 port map( B => n1507, A => n226, S => n1531, Y => n1508);
   U1529 : NAND2X1 port map( A => n1509, B => n1508, Y => n1270);
   U1530 : NAND2X1 port map( A => n219, B => currentPlainKey_63_port, Y => 
                           n1534);
   U1531 : NOR2X1 port map( A => n1511, B => n166, Y => n1512);
   U1532 : MUX2X1 port map( B => currentPlainKey_63_port, A => n189, S => n1512
                           , Y => n1516);
   U1533 : NOR2X1 port map( A => n1514, B => n1513, Y => n1515);
   U1534 : MUX2X1 port map( B => n1516, A => n220, S => n1515, Y => n1517);
   U1535 : MUX2X1 port map( B => n1517, A => n236, S => n115, Y => n1519);
   U1536 : MUX2X1 port map( B => n1520, A => n1519, S => n1518, Y => n1522);
   U1537 : MUX2X1 port map( B => n1522, A => RCV_DATA(4), S => n1521, Y => 
                           n1525);
   U1538 : INVX2 port map( A => RCV_DATA(5), Y => n1524);
   U1539 : MUX2X1 port map( B => n1525, A => n1524, S => n1523, Y => n1526);
   U1540 : NAND2X1 port map( A => n224, B => n1526, Y => n1530);
   U1541 : MUX2X1 port map( B => n1530, A => n230, S => n1528, Y => n1532);
   U1542 : MUX2X1 port map( B => n1532, A => n51, S => n1531, Y => n1533);
   U1543 : NAND2X1 port map( A => n1534, B => n1533, Y => n1269);
   U1544 : NAND2X1 port map( A => n1535, B => n1605, Y => n1547);
   U1545 : INVX2 port map( A => n1547, Y => n1536);
   U1546 : NAND3X1 port map( A => n17, B => n253, C => n1536, Y => n1545);
   U1547 : NAND2X1 port map( A => address_0_port, B => n1545, Y => n1537);
   U1548 : NAND2X1 port map( A => n1546, B => n1537, Y => n1333);
   U1549 : NAND2X1 port map( A => address_1_port, B => n1545, Y => n1538);
   U1550 : NAND2X1 port map( A => n1546, B => n1538, Y => n1334);
   U1551 : NAND2X1 port map( A => address_2_port, B => n1545, Y => n1539);
   U1552 : NAND2X1 port map( A => n1546, B => n1539, Y => n1335);
   U1553 : MUX2X1 port map( B => n192, A => keyCount_0_port, S => n1542, Y => 
                           n1540);
   U1554 : NAND2X1 port map( A => n1546, B => n1540, Y => n1336);
   U1555 : MUX2X1 port map( B => address_4_port, A => keyCount_1_port, S => 
                           n1542, Y => n1541);
   U1556 : NAND2X1 port map( A => n1546, B => n1541, Y => n1337);
   U1557 : MUX2X1 port map( B => address_5_port, A => keyCount_2_port, S => 
                           n1542, Y => n1543);
   U1558 : NAND2X1 port map( A => n1546, B => n1543, Y => n1338);
   U1559 : OAI21X1 port map( A => n1631, B => n1544, C => n1546, Y => n1339);
   U1560 : OAI21X1 port map( A => n1630, B => n1544, C => n1546, Y => n1340);
   U1561 : OAI21X1 port map( A => n1548, B => n1547, C => parityError, Y => 
                           n1551);
   U1562 : OAI21X1 port map( A => n12, B => n13, C => n1549, Y => n1550);
   U1563 : NAND2X1 port map( A => n1551, B => n1550, Y => nextParityError);
   U1564 : OAI21X1 port map( A => keyCount_0_port, B => n157, C => n135, Y => 
                           n1552);
   U1565 : INVX2 port map( A => n1552, Y => n1607);
   U1566 : NAND2X1 port map( A => n1596, B => n135, Y => n1619);
   U1567 : INVX2 port map( A => n1619, Y => n1610);
   U1568 : NAND2X1 port map( A => keyCount_0_port, B => n1610, Y => n1615);
   U1569 : MUX2X1 port map( B => n1607, A => n1615, S => n1629, Y => n1350);
   U1570 : NAND3X1 port map( A => n1597, B => n14, C => n17, Y => n1555);
   U1571 : NAND3X1 port map( A => n101, B => n253, C => n11, Y => n1554);
   U1572 : OR2X2 port map( A => n1555, B => n1554, Y => n1569);
   U1573 : NAND2X1 port map( A => n1565, B => CLR_RBUFF_port, Y => n1571);
   U1574 : INVX2 port map( A => n1571, Y => n1566);
   U1575 : NAND2X1 port map( A => N1799, B => n1566, Y => n1557);
   U1576 : NAND2X1 port map( A => parityAccumulator_7_port, B => n1569, Y => 
                           n1556);
   U1577 : NAND2X1 port map( A => n1557, B => n1556, Y => n1341);
   U1578 : NAND2X1 port map( A => N1798, B => n1566, Y => n1559);
   U1579 : NAND2X1 port map( A => parityAccumulator_6_port, B => n1569, Y => 
                           n1558);
   U1580 : NAND2X1 port map( A => n1559, B => n1558, Y => n1342);
   U1581 : NAND2X1 port map( A => N1797, B => n1566, Y => n1561);
   U1582 : NAND2X1 port map( A => n1569, B => parityAccumulator_5_port, Y => 
                           n1560);
   U1583 : NAND2X1 port map( A => n1561, B => n1560, Y => n1343);
   U1584 : NAND2X1 port map( A => N1796, B => n1566, Y => n1563);
   U1585 : NAND2X1 port map( A => n1569, B => parityAccumulator_4_port, Y => 
                           n1562);
   U1586 : NAND2X1 port map( A => n1563, B => n1562, Y => n1344);
   U1587 : INVX2 port map( A => n1569, Y => n1565);
   U1588 : NAND2X1 port map( A => N1795, B => n1566, Y => n1564);
   U1589 : OAI21X1 port map( A => n1626, B => n1565, C => n1564, Y => n1345);
   U1590 : NAND2X1 port map( A => N1794, B => n1566, Y => n1567);
   U1591 : OAI21X1 port map( A => n1625, B => n1565, C => n1567, Y => n1346);
   U1592 : INVX2 port map( A => N1793, Y => n1568);
   U1593 : OAI22X1 port map( A => n1624, B => n1565, C => n1571, D => n1568, Y 
                           => n1347);
   U1594 : INVX2 port map( A => N1792, Y => n1570);
   U1595 : OAI22X1 port map( A => n1623, B => n1565, C => n1571, D => n1570, Y 
                           => n1348);
   U1596 : AOI21X1 port map( A => n1580, B => RBUF_FULL, C => n1178, Y => n1572
                           );
   U1597 : NAND2X1 port map( A => n1572, B => n1587, Y => n1576);
   U1598 : NAND2X1 port map( A => n1574, B => n1573, Y => n1575);
   U1599 : NAND2X1 port map( A => n1575, B => n1598, Y => n1581);
   U1600 : NAND2X1 port map( A => n1576, B => n1581, Y => n1591);
   U1601 : NAND2X1 port map( A => n7, B => n1591, Y => n1577);
   U1602 : NAND2X1 port map( A => n1578, B => n1577, Y => n1354);
   U1603 : INVX2 port map( A => keyCount_3_port, Y => n1580);
   U1604 : AND2X2 port map( A => keyCount_2_port, B => keyCount_0_port, Y => 
                           n1579);
   U1605 : NAND3X1 port map( A => keyCount_1_port, B => n1580, C => n1579, Y =>
                           n1595);
   U1606 : INVX2 port map( A => n1595, Y => n1611);
   U1607 : INVX2 port map( A => n1581, Y => n1594);
   U1608 : AOI22X1 port map( A => n1611, B => n1596, C => n1594, D => n9, Y => 
                           n1590);
   U1609 : INVX2 port map( A => RBUF_FULL, Y => n1582);
   U1610 : NAND2X1 port map( A => n1583, B => n1582, Y => n1589);
   U1611 : INVX2 port map( A => OE, Y => n1584);
   U1612 : NAND2X1 port map( A => n1695, B => n1584, Y => n1586);
   U1613 : NAND2X1 port map( A => n1597, B => n17, Y => n1585);
   U1614 : AOI21X1 port map( A => n1587, B => n1586, C => n1585, Y => n1588);
   U1615 : NAND3X1 port map( A => n1590, B => n1589, C => n1588, Y => n1352);
   U1616 : AOI21X1 port map( A => n85, B => n1591, C => n1596, Y => n1592);
   U1617 : NAND3X1 port map( A => n1597, B => n47, C => n1592, Y => n1351);
   U1618 : AOI22X1 port map( A => n1596, B => n1595, C => n1594, D => n194, Y 
                           => n1606);
   U1619 : NAND2X1 port map( A => n1598, B => n1597, Y => n1603);
   U1620 : NAND2X1 port map( A => n1695, B => n1584, Y => n1601);
   U1621 : OAI21X1 port map( A => n1601, B => n14, C => n17, Y => n1602);
   U1622 : AOI21X1 port map( A => RBUF_FULL, B => n1603, C => n1602, Y => n1604
                           );
   U1623 : NAND3X1 port map( A => n1606, B => n1605, C => n1604, Y => n1353);
   U1624 : NOR2X1 port map( A => keyCount_2_port, B => n157, Y => n1609);
   U1625 : OAI21X1 port map( A => keyCount_1_port, B => n157, C => n1607, Y => 
                           n1614);
   U1626 : OAI21X1 port map( A => n1609, B => n1614, C => keyCount_3_port, Y =>
                           n1613);
   U1627 : NAND2X1 port map( A => n1611, B => n1610, Y => n1612);
   U1628 : NAND2X1 port map( A => n1613, B => n1612, Y => n1355);
   U1629 : INVX2 port map( A => n1614, Y => n1618);
   U1630 : INVX2 port map( A => n1615, Y => n1616);
   U1631 : NAND2X1 port map( A => n1616, B => keyCount_1_port, Y => n1617);
   U1632 : MUX2X1 port map( B => n1618, A => n1617, S => n1621, Y => n1349);
   U1633 : MUX2X1 port map( B => n1619, A => n135, S => keyCount_0_port, Y => 
                           n1356);
   U1634 : INVX2 port map( A => keyCount_2_port, Y => n1621);
   U1635 : INVX2 port map( A => parityAccumulator_0_port, Y => n1623);
   U1636 : INVX2 port map( A => parityAccumulator_1_port, Y => n1624);
   U1637 : INVX2 port map( A => parityAccumulator_2_port, Y => n1625);
   U1638 : INVX2 port map( A => parityAccumulator_3_port, Y => n1626);
   U1639 : INVX2 port map( A => keyCount_1_port, Y => n1629);
   U1640 : INVX2 port map( A => address_7_port, Y => n1630);
   U1641 : INVX2 port map( A => address_6_port, Y => n1631);
   U1642 : INVX2 port map( A => currentPlainKey_61_port, Y => n1633);
   U1643 : INVX2 port map( A => currentPlainKey_60_port, Y => n1634);
   U1644 : INVX2 port map( A => currentPlainKey_59_port, Y => n1635);
   U1645 : INVX2 port map( A => currentPlainKey_58_port, Y => n1636);
   U1646 : INVX2 port map( A => currentPlainKey_57_port, Y => n1637);
   U1647 : INVX2 port map( A => currentPlainKey_56_port, Y => n1638);
   U1648 : INVX2 port map( A => currentPlainKey_55_port, Y => n1639);
   U1649 : INVX2 port map( A => currentPlainKey_54_port, Y => n1640);
   U1650 : INVX2 port map( A => currentPlainKey_53_port, Y => n1641);
   U1651 : INVX2 port map( A => currentPlainKey_52_port, Y => n1642);
   U1652 : INVX2 port map( A => currentPlainKey_51_port, Y => n1643);
   U1653 : INVX2 port map( A => currentPlainKey_50_port, Y => n1644);
   U1654 : INVX2 port map( A => currentPlainKey_49_port, Y => n1645);
   U1655 : INVX2 port map( A => currentPlainKey_48_port, Y => n1646);
   U1656 : INVX2 port map( A => currentPlainKey_47_port, Y => n1647);
   U1657 : INVX2 port map( A => currentPlainKey_46_port, Y => n1648);
   U1658 : INVX2 port map( A => currentPlainKey_45_port, Y => n1649);
   U1659 : INVX2 port map( A => currentPlainKey_44_port, Y => n1650);
   U1660 : INVX2 port map( A => currentPlainKey_43_port, Y => n1651);
   U1661 : INVX2 port map( A => currentPlainKey_42_port, Y => n1652);
   U1662 : INVX2 port map( A => currentPlainKey_41_port, Y => n1653);
   U1663 : INVX2 port map( A => currentPlainKey_40_port, Y => n1654);
   U1664 : INVX2 port map( A => currentPlainKey_39_port, Y => n1655);
   U1665 : INVX2 port map( A => currentPlainKey_38_port, Y => n1656);
   U1666 : INVX2 port map( A => currentPlainKey_37_port, Y => n1657);
   U1667 : INVX2 port map( A => currentPlainKey_36_port, Y => n1658);
   U1668 : INVX2 port map( A => currentPlainKey_35_port, Y => n1659);
   U1669 : INVX2 port map( A => currentPlainKey_34_port, Y => n1660);
   U1670 : INVX2 port map( A => currentPlainKey_33_port, Y => n1661);
   U1671 : INVX2 port map( A => currentPlainKey_32_port, Y => n1662);
   U1672 : INVX2 port map( A => currentPlainKey_31_port, Y => n1663);
   U1673 : INVX2 port map( A => currentPlainKey_30_port, Y => n1664);
   U1674 : INVX2 port map( A => currentPlainKey_29_port, Y => n1665);
   U1675 : INVX2 port map( A => currentPlainKey_28_port, Y => n1666);
   U1676 : INVX2 port map( A => currentPlainKey_27_port, Y => n1667);
   U1677 : INVX2 port map( A => currentPlainKey_26_port, Y => n1668);
   U1678 : INVX2 port map( A => currentPlainKey_25_port, Y => n1669);
   U1679 : INVX2 port map( A => currentPlainKey_24_port, Y => n1670);
   U1680 : INVX2 port map( A => currentPlainKey_23_port, Y => n1671);
   U1681 : INVX2 port map( A => currentPlainKey_22_port, Y => n1672);
   U1682 : INVX2 port map( A => currentPlainKey_21_port, Y => n1673);
   U1683 : INVX2 port map( A => currentPlainKey_20_port, Y => n1674);
   U1684 : INVX2 port map( A => currentPlainKey_19_port, Y => n1675);
   U1685 : INVX2 port map( A => currentPlainKey_18_port, Y => n1676);
   U1686 : INVX2 port map( A => currentPlainKey_17_port, Y => n1677);
   U1687 : INVX2 port map( A => currentPlainKey_16_port, Y => n1678);
   U1688 : INVX2 port map( A => currentPlainKey_15_port, Y => n1679);
   U1689 : INVX2 port map( A => currentPlainKey_14_port, Y => n1680);
   U1690 : INVX2 port map( A => currentPlainKey_13_port, Y => n1681);
   U1691 : INVX2 port map( A => currentPlainKey_12_port, Y => n1682);
   U1692 : INVX2 port map( A => currentPlainKey_11_port, Y => n1683);
   U1693 : INVX2 port map( A => currentPlainKey_10_port, Y => n1684);
   U1694 : INVX2 port map( A => currentPlainKey_9_port, Y => n1685);
   U1695 : INVX2 port map( A => currentPlainKey_8_port, Y => n1686);
   U1696 : INVX2 port map( A => currentPlainKey_7_port, Y => n1687);
   U1697 : INVX2 port map( A => currentPlainKey_6_port, Y => n1688);
   U1698 : INVX2 port map( A => currentPlainKey_5_port, Y => n1689);
   U1699 : INVX2 port map( A => currentPlainKey_4_port, Y => n1690);
   U1700 : INVX2 port map( A => SBE, Y => n1695);

end SYN_keyb;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_sr_10bit_1 is

   port( CLK, RST, SHIFT_STROBE, SERIAL_IN : in std_logic;  LOAD_DATA : out 
         std_logic_vector (7 downto 0);  STOP_DATA : out std_logic_vector (1 
         downto 0));

end uart_sr_10bit_1;

architecture SYN_dataflow of uart_sr_10bit_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal LOAD_DATA_7_port, LOAD_DATA_6_port, LOAD_DATA_5_port, 
      LOAD_DATA_4_port, LOAD_DATA_3_port, LOAD_DATA_2_port, LOAD_DATA_1_port, 
      LOAD_DATA_0_port, STOP_DATA_1_port, STOP_DATA_0_port, n3, n12, n14, n16, 
      n18, n20, n22, n24, n26, n28, n30, n32, n33, n1, n2, n4, n5, n6, n7, n8, 
      n9, n10, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, n34, n35 
      : std_logic;

begin
   LOAD_DATA <= ( LOAD_DATA_7_port, LOAD_DATA_6_port, LOAD_DATA_5_port, 
      LOAD_DATA_4_port, LOAD_DATA_3_port, LOAD_DATA_2_port, LOAD_DATA_1_port, 
      LOAD_DATA_0_port );
   STOP_DATA <= ( STOP_DATA_1_port, STOP_DATA_0_port );
   
   present_val_reg_9_inst : DFFSR port map( D => n33, CLK => CLK, R => n15, S 
                           => n32, Q => STOP_DATA_1_port);
   U2 : OAI21X1 port map( A => n35, B => n17, C => n3, Y => n14);
   U3 : NAND2X1 port map( A => LOAD_DATA_0_port, B => n17, Y => n3);
   U4 : OAI22X1 port map( A => n17, B => n34, C => n13, D => n35, Y => n16);
   U6 : OAI22X1 port map( A => n17, B => n31, C => n13, D => n34, Y => n18);
   U8 : OAI22X1 port map( A => n17, B => n29, C => n13, D => n31, Y => n20);
   U10 : OAI22X1 port map( A => n17, B => n27, C => n13, D => n29, Y => n22);
   U12 : OAI22X1 port map( A => n17, B => n25, C => n13, D => n27, Y => n24);
   U14 : OAI22X1 port map( A => n17, B => n23, C => n13, D => n25, Y => n26);
   U16 : OAI22X1 port map( A => n17, B => n21, C => n13, D => n23, Y => n28);
   U18 : OAI22X1 port map( A => n17, B => n19, C => n13, D => n21, Y => n30);
   U22 : OAI21X1 port map( A => n13, B => n19, C => n12, Y => n33);
   U23 : NAND2X1 port map( A => SERIAL_IN, B => n13, Y => n12);
   n32 <= '1';
   present_val_reg_8_inst : DFFSR port map( D => n30, CLK => CLK, R => n15, S 
                           => n10, Q => STOP_DATA_0_port);
   present_val_reg_7_inst : DFFSR port map( D => n28, CLK => CLK, R => n15, S 
                           => n9, Q => LOAD_DATA_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n26, CLK => CLK, R => n15, S 
                           => n8, Q => LOAD_DATA_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n24, CLK => CLK, R => n15, S 
                           => n7, Q => LOAD_DATA_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n22, CLK => CLK, R => n15, S 
                           => n6, Q => LOAD_DATA_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n20, CLK => CLK, R => n15, S 
                           => n5, Q => LOAD_DATA_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n18, CLK => CLK, R => n15, S 
                           => n4, Q => LOAD_DATA_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n16, CLK => CLK, R => n15, S 
                           => n2, Q => LOAD_DATA_1_port);
   present_val_reg_0_inst : DFFSR port map( D => n14, CLK => CLK, R => n15, S 
                           => n1, Q => LOAD_DATA_0_port);
   n1 <= '1';
   n2 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   U21 : INVX2 port map( A => RST, Y => n15);
   U24 : INVX2 port map( A => n13, Y => n17);
   U25 : INVX4 port map( A => n11, Y => n13);
   U26 : INVX2 port map( A => SHIFT_STROBE, Y => n11);
   U27 : INVX2 port map( A => STOP_DATA_1_port, Y => n19);
   U28 : INVX2 port map( A => STOP_DATA_0_port, Y => n21);
   U29 : INVX2 port map( A => LOAD_DATA_7_port, Y => n23);
   U30 : INVX2 port map( A => LOAD_DATA_6_port, Y => n25);
   U31 : INVX2 port map( A => LOAD_DATA_5_port, Y => n27);
   U32 : INVX2 port map( A => LOAD_DATA_4_port, Y => n29);
   U33 : INVX2 port map( A => LOAD_DATA_3_port, Y => n31);
   U35 : INVX2 port map( A => LOAD_DATA_2_port, Y => n34);
   U36 : INVX2 port map( A => LOAD_DATA_1_port, Y => n35);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_sb_check_1 is

   port( RST, CLK, SBC_CLR, SBC_EN : in std_logic;  STOP_DATA : in 
         std_logic_vector (1 downto 0);  SB_DETECT, SBE : out std_logic);

end uart_sb_check_1;

architecture SYN_behavioral of uart_sb_check_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal SBE_prime, sb_detect_flag, n1, n3, n7, n8, n9, n2, n4, n5, n6 : 
      std_logic;

begin
   
   SB_DETECT_reg : DFFSR port map( D => sb_detect_flag, CLK => CLK, R => n2, S 
                           => n3, Q => SB_DETECT);
   SBE_reg : DFFSR port map( D => SBE_prime, CLK => CLK, R => n2, S => n1, Q =>
                           SBE);
   n1 <= '1';
   n3 <= '1';
   U6 : OR2X2 port map( A => SBC_CLR, B => STOP_DATA(0), Y => n7);
   U10 : NOR2X1 port map( A => n7, B => n8, Y => sb_detect_flag);
   U11 : NAND2X1 port map( A => STOP_DATA(1), B => SBC_EN, Y => n8);
   U12 : NOR2X1 port map( A => n6, B => n9, Y => SBE_prime);
   U13 : OAI21X1 port map( A => STOP_DATA(0), B => n4, C => n5, Y => n9);
   U4 : INVX2 port map( A => RST, Y => n2);
   U7 : INVX2 port map( A => STOP_DATA(1), Y => n4);
   U8 : INVX2 port map( A => SBC_CLR, Y => n5);
   U9 : INVX2 port map( A => SBC_EN, Y => n6);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_buf_full_1 is

   port( CLK, RST, CLR_RBUF, SET_RBUF_FULL : in std_logic;  RBUF_FULL : out 
         std_logic);

end uart_rcv_buf_full_1;

architecture SYN_Behavioral of uart_rcv_buf_full_1 is

   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal RBUF_FULL_port, n1, n2, n3 : std_logic;

begin
   RBUF_FULL <= RBUF_FULL_port;
   
   Q_int_reg : DFFSR port map( D => n3, CLK => CLK, R => n1, S => n2, Q => 
                           RBUF_FULL_port);
   U3 : NOR2X1 port map( A => RST, B => CLR_RBUF, Y => n1);
   n2 <= '1';
   U4 : OR2X2 port map( A => RBUF_FULL_port, B => SET_RBUF_FULL, Y => n3);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_buf_1 is

   port( CLK, RST, LOAD_RBUF : in std_logic;  LOAD_DATA : in std_logic_vector 
         (7 downto 0);  RCV_DATA : out std_logic_vector (7 downto 0));

end uart_rcv_buf_1;

architecture SYN_Behavioral of uart_rcv_buf_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, n1, 
      n3, n4, n5, n6, n7, n8, n9, n10, n12, n14, n16, n18, n20, n22, n25, n2, 
      n11, n13, n15, n17, n19, n21, n23, n24, n26 : std_logic;

begin
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   Q_int_reg_7_inst : DFFSR port map( D => n11, CLK => CLK, R => n2, S => n25, 
                           Q => RCV_DATA_7_port);
   Q_int_reg_6_inst : DFFSR port map( D => n13, CLK => CLK, R => n2, S => n22, 
                           Q => RCV_DATA_6_port);
   Q_int_reg_5_inst : DFFSR port map( D => n15, CLK => CLK, R => n2, S => n20, 
                           Q => RCV_DATA_5_port);
   Q_int_reg_4_inst : DFFSR port map( D => n17, CLK => CLK, R => n2, S => n18, 
                           Q => RCV_DATA_4_port);
   Q_int_reg_3_inst : DFFSR port map( D => n19, CLK => CLK, R => n2, S => n16, 
                           Q => RCV_DATA_3_port);
   Q_int_reg_2_inst : DFFSR port map( D => n21, CLK => CLK, R => n2, S => n14, 
                           Q => RCV_DATA_2_port);
   Q_int_reg_1_inst : DFFSR port map( D => n23, CLK => CLK, R => n2, S => n12, 
                           Q => RCV_DATA_1_port);
   Q_int_reg_0_inst : DFFSR port map( D => n24, CLK => CLK, R => n2, S => n10, 
                           Q => RCV_DATA_0_port);
   U3 : AOI22X1 port map( A => LOAD_RBUF, B => LOAD_DATA(0), C => 
                           RCV_DATA_0_port, D => n26, Y => n1);
   U5 : AOI22X1 port map( A => LOAD_DATA(1), B => LOAD_RBUF, C => 
                           RCV_DATA_1_port, D => n26, Y => n3);
   U7 : AOI22X1 port map( A => LOAD_DATA(2), B => LOAD_RBUF, C => 
                           RCV_DATA_2_port, D => n26, Y => n4);
   U9 : AOI22X1 port map( A => LOAD_DATA(3), B => LOAD_RBUF, C => 
                           RCV_DATA_3_port, D => n26, Y => n5);
   U11 : AOI22X1 port map( A => LOAD_DATA(4), B => LOAD_RBUF, C => 
                           RCV_DATA_4_port, D => n26, Y => n6);
   U13 : AOI22X1 port map( A => LOAD_DATA(5), B => LOAD_RBUF, C => 
                           RCV_DATA_5_port, D => n26, Y => n7);
   U15 : AOI22X1 port map( A => LOAD_DATA(6), B => LOAD_RBUF, C => 
                           RCV_DATA_6_port, D => n26, Y => n8);
   U18 : AOI22X1 port map( A => LOAD_DATA(7), B => LOAD_RBUF, C => 
                           RCV_DATA_7_port, D => n26, Y => n9);
   n10 <= '1';
   n12 <= '1';
   n14 <= '1';
   n16 <= '1';
   n18 <= '1';
   n20 <= '1';
   n22 <= '1';
   n25 <= '1';
   U2 : INVX2 port map( A => RST, Y => n2);
   U4 : INVX2 port map( A => n9, Y => n11);
   U6 : INVX2 port map( A => n8, Y => n13);
   U8 : INVX2 port map( A => n7, Y => n15);
   U10 : INVX2 port map( A => n6, Y => n17);
   U12 : INVX2 port map( A => n5, Y => n19);
   U14 : INVX2 port map( A => n4, Y => n21);
   U16 : INVX2 port map( A => n3, Y => n23);
   U17 : INVX2 port map( A => n1, Y => n24);
   U19 : INVX2 port map( A => LOAD_RBUF, Y => n26);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcu_1 is

   port( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT : in std_logic;  RBUF_LOAD
         , TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR : out 
         std_logic);

end uart_rcu_1;

architecture SYN_rcub of uart_rcu_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal RBUF_LOAD_port, TIMER_TRIG_port, CHK_ERROR_port, SET_RBUF_FULL_port, 
      SBC_EN_port, SBC_CLR_port, state_2_port, state_1_port, state_0_port, 
      timerRunning, count_7_port, count_6_port, count_5_port, count_4_port, 
      count_3_port, count_2_port, count_1_port, count_0_port, nextCount_7_port,
      nextCount_6_port, nextCount_5_port, nextCount_4_port, nextCount_3_port, 
      nextCount_2_port, nextCount_1_port, nextCount_0_port, nextState_1_port, 
      nextState_0_port, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, 
      N35, N36, N37, N38, N99, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24_port, n26_port, n27_port, n28_port, 
      n29_port, n30_port, n31_port, n33_port, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      add_46_carry_3_port, add_46_carry_4_port, add_46_carry_5_port, 
      add_46_carry_6_port, n1, n2, n3, n4, n5, n6, n7, n25_port, n32_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n81, n82 : std_logic;

begin
   RBUF_LOAD <= RBUF_LOAD_port;
   TIMER_TRIG <= TIMER_TRIG_port;
   CHK_ERROR <= CHK_ERROR_port;
   SET_RBUF_FULL <= SET_RBUF_FULL_port;
   SBC_EN <= SBC_EN_port;
   SBC_CLR <= SBC_CLR_port;
   
   count_reg_0_inst : DFFSR port map( D => nextCount_0_port, CLK => CLK, R => 
                           n5, S => n33_port, Q => count_0_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n4, S => n31_port, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => n43, CLK => CLK, R => n4, S => 
                           n30_port, Q => state_2_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n4, S => n29_port, Q => state_0_port);
   SBC_CLR_reg : DFFSR port map( D => n78, CLK => CLK, R => n4, S => n28_port, 
                           Q => SBC_CLR_port);
   TIMER_TRIG_reg : DFFSR port map( D => n79, CLK => CLK, R => n4, S => 
                           n27_port, Q => TIMER_TRIG_port);
   RBUF_LOAD_reg : DFFSR port map( D => n80, CLK => CLK, R => n4, S => n26_port
                           , Q => RBUF_LOAD_port);
   timerRunning_reg : DFFSR port map( D => n74, CLK => CLK, R => n4, S => 
                           n24_port, Q => timerRunning);
   nextCount_reg_1_inst : DFFSR port map( D => N32, CLK => CLK, R => n4, S => 
                           n23, Q => nextCount_1_port);
   count_reg_1_inst : DFFSR port map( D => nextCount_1_port, CLK => CLK, R => 
                           n4, S => n22, Q => count_1_port);
   nextCount_reg_0_inst : DFFSR port map( D => N31, CLK => CLK, R => n21, S => 
                           n5, Q => nextCount_0_port);
   nextCount_reg_2_inst : DFFSR port map( D => N33, CLK => CLK, R => n4, S => 
                           n20, Q => nextCount_2_port);
   count_reg_2_inst : DFFSR port map( D => nextCount_2_port, CLK => CLK, R => 
                           n5, S => n19, Q => count_2_port);
   nextCount_reg_3_inst : DFFSR port map( D => N34, CLK => CLK, R => n5, S => 
                           n18, Q => nextCount_3_port);
   count_reg_3_inst : DFFSR port map( D => nextCount_3_port, CLK => CLK, R => 
                           n5, S => n17, Q => count_3_port);
   nextCount_reg_4_inst : DFFSR port map( D => N35, CLK => CLK, R => n5, S => 
                           n16, Q => nextCount_4_port);
   count_reg_4_inst : DFFSR port map( D => nextCount_4_port, CLK => CLK, R => 
                           n5, S => n15, Q => count_4_port);
   nextCount_reg_5_inst : DFFSR port map( D => N36, CLK => CLK, R => n5, S => 
                           n14, Q => nextCount_5_port);
   count_reg_5_inst : DFFSR port map( D => nextCount_5_port, CLK => CLK, R => 
                           n5, S => n13, Q => count_5_port);
   nextCount_reg_6_inst : DFFSR port map( D => N37, CLK => CLK, R => n5, S => 
                           n12, Q => nextCount_6_port);
   count_reg_6_inst : DFFSR port map( D => nextCount_6_port, CLK => CLK, R => 
                           n5, S => n11, Q => count_6_port);
   nextCount_reg_7_inst : DFFSR port map( D => N38, CLK => CLK, R => n5, S => 
                           n10, Q => nextCount_7_port);
   count_reg_7_inst : DFFSR port map( D => nextCount_7_port, CLK => CLK, R => 
                           n5, S => n9, Q => count_7_port);
   SBC_EN_reg : DFFSR port map( D => n76, CLK => CLK, R => n4, S => n8, Q => 
                           SBC_EN_port);
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   n18 <= '1';
   n19 <= '1';
   n20 <= '1';
   n21 <= '1';
   n22 <= '1';
   n23 <= '1';
   n24_port <= '1';
   n26_port <= '1';
   n27_port <= '1';
   n28_port <= '1';
   n29_port <= '1';
   n30_port <= '1';
   n31_port <= '1';
   n33_port <= '1';
   U33 : AND2X2 port map( A => N30, B => timerRunning, Y => N38);
   U34 : AND2X2 port map( A => N29, B => timerRunning, Y => N37);
   U35 : AND2X2 port map( A => N28, B => timerRunning, Y => N36);
   U36 : AND2X2 port map( A => N27, B => timerRunning, Y => N35);
   U37 : AND2X2 port map( A => N26, B => timerRunning, Y => N34);
   U38 : AND2X2 port map( A => N25, B => timerRunning, Y => N33);
   U39 : AND2X2 port map( A => N24, B => timerRunning, Y => N32);
   U54 : OAI21X1 port map( A => n49, B => n45, C => n50, Y => n48);
   U55 : OAI21X1 port map( A => n46, B => n44, C => n45, Y => n50);
   U56 : NAND2X1 port map( A => n51, B => n52, Y => n74);
   U57 : OAI21X1 port map( A => n53, B => n54, C => timerRunning, Y => n52);
   U58 : NAND2X1 port map( A => n55, B => n56, Y => n54);
   U59 : NAND2X1 port map( A => n57, B => n56, Y => n75);
   U60 : NAND3X1 port map( A => n37_port, B => n51, C => CHK_ERROR_port, Y => 
                           n57);
   U61 : OAI21X1 port map( A => n58, B => n82, C => n59, Y => n76);
   U62 : NAND2X1 port map( A => n56, B => n60, Y => n58);
   U63 : NAND2X1 port map( A => n61, B => n40, Y => n56);
   U64 : NAND3X1 port map( A => n62, B => n63, C => n64, Y => n77);
   U65 : NAND3X1 port map( A => n36_port, B => n51, C => SET_RBUF_FULL_port, Y 
                           => n64);
   U66 : NAND2X1 port map( A => n60, B => n63, Y => n53);
   U67 : NAND3X1 port map( A => nextState_0_port, B => nextState_1_port, C => 
                           n61, Y => n63);
   U68 : NAND3X1 port map( A => n38_port, B => n40, C => n61, Y => n62);
   U69 : OAI21X1 port map( A => n65, B => n47, C => n51, Y => n78);
   U70 : OAI21X1 port map( A => n65, B => n81, C => n51, Y => n79);
   U71 : NAND2X1 port map( A => n60, B => n59, Y => n65);
   U72 : NAND3X1 port map( A => nextState_1_port, B => n38_port, C => n41, Y =>
                           n59);
   U73 : NAND2X1 port map( A => n66, B => n55, Y => n80);
   U74 : NAND3X1 port map( A => nextState_1_port, B => n38_port, C => n61, Y =>
                           n55);
   U75 : NAND3X1 port map( A => n60, B => n51, C => RBUF_LOAD_port, Y => n66);
   U76 : NAND3X1 port map( A => nextState_0_port, B => n40, C => n41, Y => n51)
                           ;
   U77 : NAND3X1 port map( A => n38_port, B => n40, C => n41, Y => n60);
   U78 : OAI21X1 port map( A => n42, B => n45, C => n67, Y => n61);
   U79 : NAND3X1 port map( A => state_0_port, B => n45, C => state_1_port, Y =>
                           n67);
   U80 : NAND2X1 port map( A => n68, B => n69, Y => n49);
   U81 : OAI21X1 port map( A => n70, B => n69, C => n68, Y => nextState_1_port)
                           ;
   U82 : NOR2X1 port map( A => N99, B => state_2_port, Y => n70);
   U83 : OAI21X1 port map( A => state_2_port, B => n71, C => n68, Y => 
                           nextState_0_port);
   U84 : NAND2X1 port map( A => state_1_port, B => n46, Y => n68);
   U85 : AOI21X1 port map( A => START_BIT, B => n46, C => n72, Y => n71);
   U86 : OAI21X1 port map( A => N99, B => n69, C => n73, Y => n72);
   U87 : NAND2X1 port map( A => SB_DETECT, B => state_1_port, Y => n73);
   U88 : NAND2X1 port map( A => state_0_port, B => n44, Y => n69);
   U89 : NAND2X1 port map( A => n39, B => timerRunning, Y => N31);
   SET_RBUF_FULL_reg : DFFSR port map( D => n77, CLK => CLK, R => n4, S => n2, 
                           Q => SET_RBUF_FULL_port);
   CHK_ERROR_reg : DFFSR port map( D => n75, CLK => CLK, R => n4, S => n1, Q =>
                           CHK_ERROR_port);
   n1 <= '1';
   n2 <= '1';
   U7 : INVX2 port map( A => RST, Y => n4);
   U8 : INVX2 port map( A => RST, Y => n5);
   U24 : XNOR2X1 port map( A => count_7_port, B => n3, Y => N30);
   U31 : NAND2X1 port map( A => count_6_port, B => add_46_carry_6_port, Y => n3
                           );
   U40 : XOR2X1 port map( A => add_46_carry_6_port, B => count_6_port, Y => N29
                           );
   U41 : AND2X1 port map( A => count_5_port, B => add_46_carry_5_port, Y => 
                           add_46_carry_6_port);
   U42 : XOR2X1 port map( A => add_46_carry_5_port, B => count_5_port, Y => N28
                           );
   U43 : AND2X1 port map( A => count_4_port, B => add_46_carry_4_port, Y => 
                           add_46_carry_5_port);
   U44 : XOR2X1 port map( A => add_46_carry_4_port, B => count_4_port, Y => N27
                           );
   U45 : AND2X1 port map( A => count_3_port, B => add_46_carry_3_port, Y => 
                           add_46_carry_4_port);
   U46 : XOR2X1 port map( A => add_46_carry_3_port, B => count_3_port, Y => N26
                           );
   U47 : AND2X1 port map( A => count_2_port, B => count_1_port, Y => 
                           add_46_carry_3_port);
   U48 : XOR2X1 port map( A => count_1_port, B => count_2_port, Y => N25);
   U49 : INVX2 port map( A => count_1_port, Y => N24);
   U50 : OAI21X1 port map( A => count_0_port, B => count_1_port, C => 
                           count_2_port, Y => n6);
   U51 : NOR2X1 port map( A => n35_port, B => n6, Y => n7);
   U52 : OAI21X1 port map( A => n7, B => count_4_port, C => count_6_port, Y => 
                           n25_port);
   U53 : OAI21X1 port map( A => n34_port, B => n25_port, C => n32_port, Y => 
                           N99);
   U90 : INVX2 port map( A => count_7_port, Y => n32_port);
   U91 : INVX2 port map( A => count_5_port, Y => n34_port);
   U92 : INVX2 port map( A => count_3_port, Y => n35_port);
   U93 : INVX2 port map( A => n53, Y => n36_port);
   U94 : INVX2 port map( A => n58, Y => n37_port);
   U95 : INVX2 port map( A => nextState_0_port, Y => n38_port);
   U96 : INVX2 port map( A => count_0_port, Y => n39);
   U97 : INVX2 port map( A => nextState_1_port, Y => n40);
   U98 : INVX2 port map( A => n61, Y => n41);
   U99 : INVX2 port map( A => n49, Y => n42);
   U100 : INVX2 port map( A => n48, Y => n43);
   U101 : INVX2 port map( A => state_1_port, Y => n44);
   U102 : INVX2 port map( A => state_2_port, Y => n45);
   U103 : INVX2 port map( A => state_0_port, Y => n46);
   U104 : INVX2 port map( A => SBC_CLR_port, Y => n47);
   U105 : INVX2 port map( A => TIMER_TRIG_port, Y => n81);
   U106 : INVX2 port map( A => SBC_EN_port, Y => n82);

end SYN_rcub;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_error_1 is

   port( RST, CLK, RBUF_FULL, CHK_ERROR : in std_logic;  OE : out std_logic);

end uart_error_1;

architecture SYN_behavioral of uart_error_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal OE_prime, n2, n1 : std_logic;

begin
   
   OE_reg : DFFSR port map( D => OE_prime, CLK => CLK, R => n1, S => n2, Q => 
                           OE);
   n2 <= '1';
   U5 : AND2X2 port map( A => RBUF_FULL, B => CHK_ERROR, Y => OE_prime);
   U3 : INVX2 port map( A => RST, Y => n1);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_edge_detector_1 is

   port( CLK, RST, SERIAL_IN : in std_logic;  START_BIT : out std_logic);

end uart_edge_detector_1;

architecture SYN_Behavioral of uart_edge_detector_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal Q_int, Q_int2, n1, n3, n2, n4 : std_logic;

begin
   
   Q_int_reg : DFFSR port map( D => SERIAL_IN, CLK => CLK, R => n2, S => n3, Q 
                           => Q_int);
   Q_int2_reg : DFFSR port map( D => Q_int, CLK => CLK, R => n2, S => n1, Q => 
                           Q_int2);
   n1 <= '1';
   n3 <= '1';
   U7 : NOR2X1 port map( A => Q_int, B => n4, Y => START_BIT);
   U4 : INVX2 port map( A => RST, Y => n2);
   U6 : INVX2 port map( A => Q_int2, Y => n4);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_timer_1 is

   port( CLK, RST, SENDING : in std_logic;  SHIFT_ENABLE_R, SHIFT_ENABLE_E : 
         out std_logic);

end tx_timer_1;

architecture SYN_moore of tx_timer_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal count_3_port, count_2_port, count_1_port, count_0_port, state, 
      nextcount_3_port, nextcount_2_port, nextcount_1_port, nextcount_0_port, 
      nxt_SHIFT_ENABLE_E, n1, n2, n3, n4, n5, n7, n12, n13, n14, n15, n16, n17,
      n18, n6, n8, n9, n10, n11, n19, n20, n21, n22 : std_logic;

begin
   SHIFT_ENABLE_R <= nxt_SHIFT_ENABLE_E;
   
   state_reg : DFFSR port map( D => n8, CLK => CLK, R => n9, S => n7, Q => 
                           state);
   count_reg_0_inst : DFFSR port map( D => nextcount_0_port, CLK => CLK, R => 
                           n9, S => n5, Q => count_0_port);
   count_reg_2_inst : DFFSR port map( D => nextcount_2_port, CLK => CLK, R => 
                           n9, S => n4, Q => count_2_port);
   count_reg_1_inst : DFFSR port map( D => nextcount_1_port, CLK => CLK, R => 
                           n9, S => n3, Q => count_1_port);
   count_reg_3_inst : DFFSR port map( D => nextcount_3_port, CLK => CLK, R => 
                           n9, S => n2, Q => count_3_port);
   SHIFT_ENABLE_E_reg : DFFSR port map( D => nxt_SHIFT_ENABLE_E, CLK => CLK, R 
                           => n9, S => n1, Q => SHIFT_ENABLE_E);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n7 <= '1';
   U14 : NOR2X1 port map( A => n12, B => n13, Y => nextcount_3_port);
   U15 : XNOR2X1 port map( A => count_3_port, B => n14, Y => n12);
   U16 : NOR2X1 port map( A => n15, B => n21, Y => n14);
   U17 : AOI21X1 port map( A => n16, B => state, C => n22, Y => 
                           nextcount_2_port);
   U18 : XNOR2X1 port map( A => n15, B => n21, Y => n16);
   U19 : NAND2X1 port map( A => count_1_port, B => count_0_port, Y => n15);
   U20 : NOR2X1 port map( A => n17, B => n13, Y => nextcount_1_port);
   U21 : NAND3X1 port map( A => n8, B => n18, C => state, Y => n13);
   U22 : XNOR2X1 port map( A => count_0_port, B => count_1_port, Y => n17);
   U23 : OAI21X1 port map( A => count_0_port, B => n22, C => state, Y => 
                           nextcount_0_port);
   U8 : AND2X1 port map( A => n20, B => n19, Y => n6);
   U10 : AND2X2 port map( A => SENDING, B => n6, Y => nxt_SHIFT_ENABLE_E);
   U11 : INVX2 port map( A => n22, Y => n8);
   U12 : INVX1 port map( A => SENDING, Y => n22);
   U13 : INVX2 port map( A => RST, Y => n9);
   U24 : NOR2X1 port map( A => count_0_port, B => count_2_port, Y => n11);
   U25 : INVX2 port map( A => count_1_port, Y => n10);
   U26 : NAND2X1 port map( A => n11, B => n10, Y => n18);
   U27 : INVX2 port map( A => n18, Y => n20);
   U28 : AND2X2 port map( A => count_3_port, B => state, Y => n19);
   U29 : INVX2 port map( A => count_2_port, Y => n21);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_tcu_1 is

   port( clk, rst, p_ready, t_bitstuff : in std_logic;  PRGA_OUT : in 
         std_logic_vector (7 downto 0);  prga_opcode : in std_logic_vector (1 
         downto 0);  t_crc : in std_logic_vector (15 downto 0);  sending, EOP, 
         next_byte : out std_logic;  send_data : out std_logic_vector (7 downto
         0);  t_strobe : out std_logic);

end tx_tcu_1;

architecture SYN_behavioral of tx_tcu_1 is

   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component tx_tcu_1_DW01_inc_0
      port( A : in std_logic_vector (6 downto 0);  SUM : out std_logic_vector 
            (6 downto 0));
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal send_data_7_port, send_data_6_port, send_data_5_port, 
      send_data_4_port, send_data_3_port, send_data_2_port, send_data_1_port, 
      send_data_0_port, state_2_port, state_1_port, state_0_port, count_5_port,
      count_4_port, count_3_port, count_2_port, count_1_port, count_0_port, 
      nextstate_2_port, nextstate_1_port, nextstate_0_port, flop_data_7_port, 
      flop_data_6_port, flop_data_5_port, flop_data_4_port, flop_data_3_port, 
      flop_data_2_port, flop_data_1_port, flop_data_0_port, 
      current_send_data_7_port, current_send_data_6_port, 
      current_send_data_5_port, current_send_data_4_port, 
      current_send_data_3_port, current_send_data_2_port, 
      current_send_data_1_port, current_send_data_0_port, N59, N60, N61, N62, 
      N63, N64, N65, N188, n158, n159, n160, n161, n162, n163, n164, n165, n166
      , n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
      n179, n180, n181, n182, n183, n194, n195, n196, n197, n198, n199, n200, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59_port
      , n60_port, n61_port, n62_port, n63_port, n64_port, n65_port, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n184, n185, n186, n187, n188_port, n189, n190, n191, n192, n193, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256 : std_logic;

begin
   send_data <= ( send_data_7_port, send_data_6_port, send_data_5_port, 
      send_data_4_port, send_data_3_port, send_data_2_port, send_data_1_port, 
      send_data_0_port );
   
   count_reg_0_inst : DFFSR port map( D => n200, CLK => clk, R => n25, S => 
                           n183, Q => count_0_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n25, S => n182, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n25, S => n181, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n25, S => n180, Q => state_2_port);
   count_reg_6_inst : DFFSR port map( D => n199, CLK => clk, R => n25, S => 
                           n179, Q => N188);
   count_reg_1_inst : DFFSR port map( D => n194, CLK => clk, R => n25, S => 
                           n178, Q => count_1_port);
   count_reg_5_inst : DFFSR port map( D => n198, CLK => clk, R => n25, S => 
                           n177, Q => count_5_port);
   count_reg_2_inst : DFFSR port map( D => n195, CLK => clk, R => n25, S => 
                           n176, Q => count_2_port);
   count_reg_3_inst : DFFSR port map( D => n196, CLK => clk, R => n25, S => 
                           n175, Q => count_3_port);
   count_reg_4_inst : DFFSR port map( D => n197, CLK => clk, R => n25, S => 
                           n174, Q => count_4_port);
   flop_data_reg_7_inst : DFFPOSX1 port map( D => n249, CLK => clk, Q => 
                           flop_data_7_port);
   current_send_data_reg_7_inst : DFFPOSX1 port map( D => n173, CLK => clk, Q 
                           => current_send_data_7_port);
   flop_data_reg_6_inst : DFFPOSX1 port map( D => n250, CLK => clk, Q => 
                           flop_data_6_port);
   current_send_data_reg_6_inst : DFFPOSX1 port map( D => n172, CLK => clk, Q 
                           => current_send_data_6_port);
   flop_data_reg_5_inst : DFFPOSX1 port map( D => n251, CLK => clk, Q => 
                           flop_data_5_port);
   current_send_data_reg_5_inst : DFFPOSX1 port map( D => n171, CLK => clk, Q 
                           => current_send_data_5_port);
   flop_data_reg_4_inst : DFFPOSX1 port map( D => n252, CLK => clk, Q => 
                           flop_data_4_port);
   current_send_data_reg_4_inst : DFFPOSX1 port map( D => n170, CLK => clk, Q 
                           => current_send_data_4_port);
   flop_data_reg_3_inst : DFFPOSX1 port map( D => n253, CLK => clk, Q => 
                           flop_data_3_port);
   current_send_data_reg_3_inst : DFFPOSX1 port map( D => n169, CLK => clk, Q 
                           => current_send_data_3_port);
   flop_data_reg_2_inst : DFFPOSX1 port map( D => n254, CLK => clk, Q => 
                           flop_data_2_port);
   current_send_data_reg_2_inst : DFFPOSX1 port map( D => n168, CLK => clk, Q 
                           => current_send_data_2_port);
   flop_data_reg_1_inst : DFFPOSX1 port map( D => n255, CLK => clk, Q => 
                           flop_data_1_port);
   current_send_data_reg_1_inst : DFFPOSX1 port map( D => n167, CLK => clk, Q 
                           => current_send_data_1_port);
   flop_data_reg_0_inst : DFFPOSX1 port map( D => n256, CLK => clk, Q => 
                           flop_data_0_port);
   current_send_data_reg_0_inst : DFFPOSX1 port map( D => n166, CLK => clk, Q 
                           => current_send_data_0_port);
   send_data_reg_7_inst : DFFPOSX1 port map( D => n165, CLK => clk, Q => 
                           send_data_7_port);
   send_data_reg_6_inst : DFFPOSX1 port map( D => n164, CLK => clk, Q => 
                           send_data_6_port);
   send_data_reg_5_inst : DFFPOSX1 port map( D => n163, CLK => clk, Q => 
                           send_data_5_port);
   send_data_reg_4_inst : DFFPOSX1 port map( D => n162, CLK => clk, Q => 
                           send_data_4_port);
   send_data_reg_3_inst : DFFPOSX1 port map( D => n161, CLK => clk, Q => 
                           send_data_3_port);
   send_data_reg_2_inst : DFFPOSX1 port map( D => n160, CLK => clk, Q => 
                           send_data_2_port);
   send_data_reg_1_inst : DFFPOSX1 port map( D => n159, CLK => clk, Q => 
                           send_data_1_port);
   send_data_reg_0_inst : DFFPOSX1 port map( D => n158, CLK => clk, Q => 
                           send_data_0_port);
   n174 <= '1';
   n175 <= '1';
   n176 <= '1';
   n177 <= '1';
   n178 <= '1';
   n179 <= '1';
   n180 <= '1';
   n181 <= '1';
   n182 <= '1';
   n183 <= '1';
   r80 : tx_tcu_1_DW01_inc_0 port map( A(6) => n23, A(5) => count_5_port, A(4) 
                           => n1, A(3) => n2, A(2) => n5, A(1) => count_1_port,
                           A(0) => count_0_port, SUM(6) => N65, SUM(5) => N64, 
                           SUM(4) => N63, SUM(3) => N62, SUM(2) => N61, SUM(1) 
                           => N60, SUM(0) => N59);
   U3 : INVX2 port map( A => count_2_port, Y => n186);
   U4 : INVX2 port map( A => n156, Y => n10);
   U5 : INVX2 port map( A => count_0_port, Y => n150);
   U6 : INVX2 port map( A => n186, Y => n5);
   U7 : BUFX4 port map( A => count_4_port, Y => n1);
   U8 : BUFX4 port map( A => count_3_port, Y => n2);
   U9 : INVX2 port map( A => n187, Y => n3);
   U10 : INVX2 port map( A => n118, Y => n4);
   U11 : OR2X2 port map( A => n104, B => n13, Y => n6);
   U12 : INVX1 port map( A => n134, Y => n84);
   U13 : INVX1 port map( A => n11, Y => n130);
   U14 : NAND2X1 port map( A => n147, B => n146, Y => n7);
   U15 : NAND2X1 port map( A => n8, B => n247, Y => n245);
   U16 : INVX2 port map( A => n7, Y => n8);
   U17 : INVX1 port map( A => n120, Y => n131);
   U18 : OR2X1 port map( A => n9, B => n104, Y => n114);
   U19 : NAND2X1 port map( A => n113, B => n105, Y => n9);
   U20 : AND2X2 port map( A => n5, B => n20, Y => n21);
   U21 : INVX4 port map( A => n24, Y => n30);
   U22 : INVX2 port map( A => n11, Y => n155);
   U23 : OR2X2 port map( A => n11, B => n10, Y => n133);
   U24 : OR2X2 port map( A => n188_port, B => n189, Y => n11);
   U25 : AND2X2 port map( A => n125, B => n88, Y => n12);
   U26 : INVX4 port map( A => n12, Y => n140);
   U27 : INVX1 port map( A => n105, Y => n13);
   U28 : INVX1 port map( A => n133, Y => n119);
   U29 : INVX2 port map( A => state_1_port, Y => n14);
   U30 : INVX1 port map( A => n14, Y => n15);
   U31 : INVX4 port map( A => n14, Y => n16);
   U32 : AND2X2 port map( A => count_1_port, B => n18, Y => n20);
   U33 : AND2X1 port map( A => n154, B => n118, Y => n17);
   U34 : OR2X1 port map( A => n30, B => n29, Y => n22);
   U35 : INVX2 port map( A => rst, Y => n25);
   U36 : NOR2X1 port map( A => t_bitstuff, B => n150, Y => n18);
   U37 : AND2X2 port map( A => state_2_port, B => n16, Y => n19);
   U38 : BUFX4 port map( A => N188, Y => n23);
   U39 : BUFX4 port map( A => state_0_port, Y => n24);
   U40 : XOR2X1 port map( A => n18, B => n3, Y => n109);
   U41 : XOR2X1 port map( A => n21, B => n2, Y => n93);
   U42 : XOR2X1 port map( A => n20, B => n5, Y => n98);
   U43 : OR2X2 port map( A => n22, B => n218, Y => n27);
   U44 : INVX1 port map( A => n87, Y => n118);
   U45 : INVX1 port map( A => n15, Y => n26);
   U46 : INVX2 port map( A => n23, Y => n145);
   U47 : INVX2 port map( A => state_2_port, Y => n58);
   U48 : NAND3X1 port map( A => n24, B => n58, C => n26, Y => n82);
   U49 : NAND3X1 port map( A => n16, B => n58, C => n30, Y => n87);
   U50 : NAND2X1 port map( A => n82, B => n87, Y => n63_port);
   U51 : NAND2X1 port map( A => n63_port, B => n25, Y => n50);
   U52 : NAND2X1 port map( A => state_2_port, B => n26, Y => n29);
   U53 : OAI21X1 port map( A => n184, B => n50, C => n27, Y => n216);
   U54 : NAND2X1 port map( A => n19, B => n30, Y => n59_port);
   U55 : INVX2 port map( A => n59_port, Y => n28);
   U56 : NAND2X1 port map( A => n28, B => n25, Y => n33);
   U57 : INVX2 port map( A => n29, Y => n62_port);
   U58 : NAND2X1 port map( A => n62_port, B => n30, Y => n120);
   U59 : NAND2X1 port map( A => n131, B => n25, Y => n32);
   U60 : INVX2 port map( A => t_crc(15), Y => n31);
   U61 : OAI22X1 port map( A => n157, B => n33, C => n32, D => n31, Y => n217);
   U62 : INVX2 port map( A => n32, Y => n47);
   U63 : INVX2 port map( A => n33, Y => n46);
   U64 : AOI22X1 port map( A => t_crc(14), B => n47, C => PRGA_OUT(6), D => n46
                           , Y => n221);
   U65 : INVX2 port map( A => flop_data_6_port, Y => n80);
   U66 : NAND3X1 port map( A => n241, B => n24, C => n62_port, Y => n49);
   U67 : INVX2 port map( A => t_crc(6), Y => n34);
   U68 : OAI22X1 port map( A => n50, B => n80, C => n49, D => n34, Y => n35);
   U69 : INVX2 port map( A => n35, Y => n222);
   U70 : AOI22X1 port map( A => t_crc(13), B => n47, C => PRGA_OUT(5), D => n46
                           , Y => n224);
   U71 : INVX2 port map( A => flop_data_5_port, Y => n78);
   U72 : INVX2 port map( A => t_crc(5), Y => n36);
   U73 : OAI22X1 port map( A => n50, B => n78, C => n49, D => n36, Y => n37);
   U74 : INVX2 port map( A => n37, Y => n225);
   U75 : AOI22X1 port map( A => t_crc(12), B => n47, C => PRGA_OUT(4), D => n46
                           , Y => n227);
   U76 : INVX2 port map( A => flop_data_4_port, Y => n76);
   U77 : INVX2 port map( A => t_crc(4), Y => n38);
   U78 : OAI22X1 port map( A => n50, B => n76, C => n49, D => n38, Y => n39);
   U79 : INVX2 port map( A => n39, Y => n228);
   U80 : AOI22X1 port map( A => t_crc(11), B => n47, C => PRGA_OUT(3), D => n46
                           , Y => n230);
   U81 : INVX2 port map( A => flop_data_3_port, Y => n74);
   U82 : INVX2 port map( A => t_crc(3), Y => n40);
   U83 : OAI22X1 port map( A => n50, B => n74, C => n49, D => n40, Y => n41);
   U84 : INVX2 port map( A => n41, Y => n231);
   U85 : AOI22X1 port map( A => t_crc(10), B => n47, C => PRGA_OUT(2), D => n46
                           , Y => n233);
   U86 : INVX2 port map( A => flop_data_2_port, Y => n72);
   U87 : INVX2 port map( A => t_crc(2), Y => n42);
   U88 : OAI22X1 port map( A => n50, B => n72, C => n49, D => n42, Y => n43);
   U89 : INVX2 port map( A => n43, Y => n234);
   U90 : AOI22X1 port map( A => t_crc(9), B => n47, C => PRGA_OUT(1), D => n46,
                           Y => n236);
   U91 : INVX2 port map( A => flop_data_1_port, Y => n70);
   U92 : INVX2 port map( A => t_crc(1), Y => n44);
   U93 : OAI22X1 port map( A => n50, B => n70, C => n49, D => n44, Y => n45);
   U94 : INVX2 port map( A => n45, Y => n237);
   U95 : AOI22X1 port map( A => t_crc(8), B => n47, C => PRGA_OUT(0), D => n46,
                           Y => n239);
   U96 : INVX2 port map( A => flop_data_0_port, Y => n68);
   U97 : INVX2 port map( A => t_crc(0), Y => n48);
   U98 : OAI22X1 port map( A => n50, B => n68, C => n49, D => n48, Y => n51);
   U99 : INVX2 port map( A => n51, Y => n240);
   U100 : INVX2 port map( A => count_4_port, Y => n147);
   U101 : INVX2 port map( A => count_5_port, Y => n146);
   U102 : INVX2 port map( A => n82, Y => n132);
   U103 : NAND2X1 port map( A => n149, B => n132, Y => n52);
   U104 : NOR2X1 port map( A => n148, B => n52, Y => t_strobe);
   U105 : NOR3X1 port map( A => n16, B => n24, C => state_2_port, Y => n124);
   U106 : INVX2 port map( A => p_ready, Y => n53);
   U107 : NAND2X1 port map( A => n124, B => n53, Y => n64_port);
   U108 : OAI21X1 port map( A => n156, B => n4, C => n64_port, Y => n54);
   U109 : AOI21X1 port map( A => n19, B => n24, C => n54, Y => n55);
   U110 : INVX2 port map( A => n55, Y => next_byte);
   U111 : NAND2X1 port map( A => n243, B => n23, Y => n57);
   U112 : INVX2 port map( A => n244, Y => n56);
   U113 : NAND2X1 port map( A => n62_port, B => n56, Y => n134);
   U114 : OAI22X1 port map( A => n57, B => n134, C => n154, D => n4, Y => EOP);
   U115 : NAND2X1 port map( A => n62_port, B => n145, Y => n61_port);
   U116 : NAND3X1 port map( A => n24, B => n16, C => n58, Y => n86);
   U117 : NAND2X1 port map( A => n59_port, B => n86, Y => n135);
   U118 : NOR2X1 port map( A => n135, B => n63_port, Y => n60_port);
   U119 : NAND3X1 port map( A => n120, B => n61_port, C => n60_port, Y => 
                           sending);
   U120 : INVX2 port map( A => PRGA_OUT(0), Y => n67);
   U121 : NOR3X1 port map( A => n63_port, B => n19, C => n62_port, Y => n66);
   U122 : AND2X2 port map( A => n64_port, B => n25, Y => n65_port);
   U123 : AND2X2 port map( A => n66, B => n65_port, Y => n81);
   U124 : MUX2X1 port map( B => n68, A => n67, S => n81, Y => n256);
   U125 : INVX2 port map( A => PRGA_OUT(1), Y => n69);
   U126 : MUX2X1 port map( B => n70, A => n69, S => n81, Y => n255);
   U127 : INVX2 port map( A => PRGA_OUT(2), Y => n71);
   U128 : MUX2X1 port map( B => n72, A => n71, S => n81, Y => n254);
   U129 : INVX2 port map( A => PRGA_OUT(3), Y => n73);
   U130 : MUX2X1 port map( B => n74, A => n73, S => n81, Y => n253);
   U131 : INVX2 port map( A => PRGA_OUT(4), Y => n75);
   U132 : MUX2X1 port map( B => n76, A => n75, S => n81, Y => n252);
   U133 : INVX2 port map( A => PRGA_OUT(5), Y => n77);
   U134 : MUX2X1 port map( B => n78, A => n77, S => n81, Y => n251);
   U135 : INVX2 port map( A => PRGA_OUT(6), Y => n79);
   U136 : MUX2X1 port map( B => n80, A => n79, S => n81, Y => n250);
   U137 : MUX2X1 port map( B => n184, A => n157, S => n81, Y => n249);
   U138 : OAI21X1 port map( A => n155, B => n120, C => n82, Y => n83);
   U139 : NAND2X1 port map( A => t_bitstuff, B => n132, Y => n94);
   U140 : OAI21X1 port map( A => n84, B => n83, C => n94, Y => n85);
   U141 : INVX2 port map( A => n85, Y => n139);
   U142 : NAND2X1 port map( A => N63, B => n139, Y => n92);
   U143 : NAND2X1 port map( A => n2, B => n21, Y => n102);
   U144 : OR2X2 port map( A => n155, B => n86, Y => n125);
   U145 : NAND2X1 port map( A => n118, B => n133, Y => n88);
   U146 : NOR2X1 port map( A => n102, B => n12, Y => n90);
   U147 : NAND2X1 port map( A => n102, B => n140, Y => n89);
   U148 : NAND2X1 port map( A => n89, B => n94, Y => n104);
   U149 : MUX2X1 port map( B => n90, A => n104, S => n1, Y => n91);
   U150 : NAND2X1 port map( A => n92, B => n91, Y => n197);
   U151 : NAND2X1 port map( A => N62, B => n139, Y => n97);
   U152 : NAND2X1 port map( A => n93, B => n140, Y => n96);
   U153 : INVX2 port map( A => n94, Y => n142);
   U154 : NAND2X1 port map( A => n142, B => n2, Y => n95);
   U155 : NAND3X1 port map( A => n97, B => n96, C => n95, Y => n196);
   U156 : NAND2X1 port map( A => N61, B => n139, Y => n101);
   U157 : NAND2X1 port map( A => n98, B => n140, Y => n100);
   U158 : NAND2X1 port map( A => n142, B => n5, Y => n99);
   U159 : NAND3X1 port map( A => n101, B => n100, C => n99, Y => n195);
   U160 : NAND2X1 port map( A => N64, B => n139, Y => n108);
   U161 : INVX2 port map( A => n102, Y => n103);
   U162 : NAND3X1 port map( A => n103, B => n1, C => n140, Y => n112);
   U163 : INVX2 port map( A => n112, Y => n106);
   U164 : NAND2X1 port map( A => n140, B => n147, Y => n105);
   U165 : MUX2X1 port map( B => n106, A => n6, S => count_5_port, Y => n107);
   U166 : NAND2X1 port map( A => n108, B => n107, Y => n198);
   U167 : AOI22X1 port map( A => n109, B => n140, C => N60, D => n139, Y => 
                           n111);
   U168 : NAND2X1 port map( A => n142, B => n3, Y => n110);
   U169 : NAND2X1 port map( A => n111, B => n110, Y => n194);
   U170 : NAND2X1 port map( A => N65, B => n139, Y => n117);
   U171 : NOR2X1 port map( A => n146, B => n112, Y => n115);
   U172 : NAND2X1 port map( A => n140, B => n146, Y => n113);
   U173 : MUX2X1 port map( B => n115, A => n114, S => n23, Y => n116);
   U174 : NAND2X1 port map( A => n117, B => n116, Y => n199);
   U175 : NAND2X1 port map( A => n151, B => p_ready, Y => n123);
   U176 : NAND2X1 port map( A => n119, B => n17, Y => n122);
   U177 : AND2X2 port map( A => n120, B => n134, Y => n121);
   U178 : NAND3X1 port map( A => n123, B => n122, C => n121, Y => 
                           nextstate_2_port);
   U179 : NAND2X1 port map( A => n124, B => p_ready, Y => n129);
   U180 : NAND2X1 port map( A => n17, B => n133, Y => n128);
   U181 : INVX2 port map( A => n125, Y => n126);
   U182 : AOI21X1 port map( A => n152, B => n132, C => n126, Y => n127);
   U183 : NAND3X1 port map( A => n129, B => n128, C => n127, Y => 
                           nextstate_1_port);
   U184 : AOI22X1 port map( A => n153, B => n132, C => n131, D => n130, Y => 
                           n138);
   U185 : NAND3X1 port map( A => n17, B => n133, C => p_ready, Y => n137);
   U186 : NOR2X1 port map( A => n135, B => n84, Y => n136);
   U187 : NAND3X1 port map( A => n138, B => n137, C => n136, Y => 
                           nextstate_0_port);
   U188 : XOR2X1 port map( A => n150, B => t_bitstuff, Y => n141);
   U189 : AOI22X1 port map( A => n141, B => n140, C => N59, D => n139, Y => 
                           n144);
   U190 : NAND2X1 port map( A => n142, B => count_0_port, Y => n143);
   U191 : NAND2X1 port map( A => n144, B => n143, Y => n200);
   U192 : NAND2X1 port map( A => n145, B => n150, Y => n148);
   U203 : NOR2X1 port map( A => n16, B => n24, Y => n151);
   U204 : INVX1 port map( A => n153, Y => n152);
   U205 : NAND3X1 port map( A => n149, B => n145, C => count_0_port, Y => n153)
                           ;
   U206 : AND2X1 port map( A => prga_opcode(1), B => prga_opcode(0), Y => n156)
                           ;
   U207 : NAND3X1 port map( A => n1, B => count_1_port, C => count_5_port, Y =>
                           n189);
   U208 : NAND3X1 port map( A => count_0_port, B => n2, C => n190, Y => 
                           n188_port);
   U209 : NOR2X1 port map( A => n23, B => n186, Y => n190);
   U210 : INVX1 port map( A => count_1_port, Y => n187);
   U211 : OAI21X1 port map( A => n191, B => n192, C => n193, Y => n173);
   U212 : INVX1 port map( A => current_send_data_7_port, Y => n192);
   U213 : OAI21X1 port map( A => n191, B => n201, C => n202, Y => n172);
   U214 : INVX1 port map( A => current_send_data_6_port, Y => n201);
   U215 : OAI21X1 port map( A => n191, B => n203, C => n204, Y => n171);
   U216 : INVX1 port map( A => current_send_data_5_port, Y => n203);
   U217 : OAI21X1 port map( A => n191, B => n205, C => n206, Y => n170);
   U218 : INVX1 port map( A => current_send_data_4_port, Y => n205);
   U219 : OAI21X1 port map( A => n191, B => n207, C => n208, Y => n169);
   U220 : INVX1 port map( A => current_send_data_3_port, Y => n207);
   U221 : OAI21X1 port map( A => n191, B => n209, C => n210, Y => n168);
   U222 : INVX1 port map( A => current_send_data_2_port, Y => n209);
   U223 : OAI21X1 port map( A => n191, B => n211, C => n212, Y => n167);
   U224 : INVX1 port map( A => current_send_data_1_port, Y => n211);
   U225 : OAI21X1 port map( A => n191, B => n213, C => n214, Y => n166);
   U226 : INVX1 port map( A => current_send_data_0_port, Y => n213);
   U227 : AOI21X1 port map( A => n24, B => n16, C => rst, Y => n191);
   U228 : NAND2X1 port map( A => n215, B => n193, Y => n165);
   U229 : NOR2X1 port map( A => n216, B => n217, Y => n193);
   U230 : INVX1 port map( A => PRGA_OUT(7), Y => n157);
   U231 : OAI21X1 port map( A => n23, B => t_crc(7), C => n25, Y => n218);
   U232 : INVX1 port map( A => flop_data_7_port, Y => n184);
   U233 : AOI22X1 port map( A => n219, B => current_send_data_7_port, C => 
                           send_data_7_port, D => rst, Y => n215);
   U234 : NAND2X1 port map( A => n220, B => n202, Y => n164);
   U235 : AND2X1 port map( A => n221, B => n222, Y => n202);
   U236 : AOI22X1 port map( A => n219, B => current_send_data_6_port, C => 
                           send_data_6_port, D => rst, Y => n220);
   U237 : NAND2X1 port map( A => n223, B => n204, Y => n163);
   U238 : AND2X1 port map( A => n224, B => n225, Y => n204);
   U239 : AOI22X1 port map( A => n219, B => current_send_data_5_port, C => 
                           send_data_5_port, D => rst, Y => n223);
   U240 : NAND2X1 port map( A => n226, B => n206, Y => n162);
   U241 : AND2X1 port map( A => n227, B => n228, Y => n206);
   U242 : AOI22X1 port map( A => n219, B => current_send_data_4_port, C => 
                           send_data_4_port, D => rst, Y => n226);
   U243 : NAND2X1 port map( A => n229, B => n208, Y => n161);
   U244 : AND2X1 port map( A => n230, B => n231, Y => n208);
   U245 : AOI22X1 port map( A => n219, B => current_send_data_3_port, C => 
                           send_data_3_port, D => rst, Y => n229);
   U246 : NAND2X1 port map( A => n232, B => n210, Y => n160);
   U247 : AND2X1 port map( A => n233, B => n234, Y => n210);
   U248 : AOI22X1 port map( A => n219, B => current_send_data_2_port, C => 
                           send_data_2_port, D => rst, Y => n232);
   U249 : NAND2X1 port map( A => n235, B => n212, Y => n159);
   U250 : AND2X1 port map( A => n236, B => n237, Y => n212);
   U251 : AOI22X1 port map( A => n219, B => current_send_data_1_port, C => 
                           send_data_1_port, D => rst, Y => n235);
   U252 : NAND2X1 port map( A => n238, B => n214, Y => n158);
   U253 : AND2X1 port map( A => n239, B => n240, Y => n214);
   U254 : NOR2X1 port map( A => rst, B => n23, Y => n241);
   U255 : AOI22X1 port map( A => n219, B => current_send_data_0_port, C => 
                           send_data_0_port, D => rst, Y => n238);
   U256 : INVX1 port map( A => n242, Y => n219);
   U257 : NAND3X1 port map( A => n24, B => n25, C => n16, Y => n242);
   U258 : OAI21X1 port map( A => n245, B => n246, C => n24, Y => n244);
   U259 : NAND3X1 port map( A => n5, B => n23, C => n2, Y => n246);
   U260 : NOR2X1 port map( A => count_1_port, B => count_0_port, Y => n247);
   U261 : NAND3X1 port map( A => n149, B => n150, C => n23, Y => n154);
   U262 : NOR2X1 port map( A => n243, B => count_1_port, Y => n149);
   U263 : NAND3X1 port map( A => n186, B => n185, C => n248, Y => n243);
   U264 : NOR2X1 port map( A => count_5_port, B => n1, Y => n248);
   U265 : INVX1 port map( A => count_3_port, Y => n185);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_shiftreg_1 is

   port( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe : in std_logic;  
         send_data : in std_logic_vector (7 downto 0);  d_encode : out 
         std_logic);

end tx_shiftreg_1;

architecture SYN_dataflow of tx_shiftreg_1 is

   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal d_encode_port, present_val_7_port, present_val_6_port, 
      present_val_5_port, present_val_4_port, present_val_3_port, 
      present_val_2_port, present_val_1_port, count_2_port, count_1_port, 
      count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n11, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69 : std_logic;

begin
   d_encode <= d_encode_port;
   
   count_reg_0_inst : DFFSR port map( D => n53, CLK => clk, R => n12, S => n17,
                           Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => n51, CLK => clk, R => n10, S => n17,
                           Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n52, CLK => clk, R => n9, S => n17, 
                           Q => count_2_port);
   present_val_reg_7_inst : DFFSR port map( D => n44, CLK => clk, R => n17, S 
                           => n8, Q => present_val_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n45, CLK => clk, R => n17, S 
                           => n7, Q => present_val_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n46, CLK => clk, R => n17, S 
                           => n6, Q => present_val_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n47, CLK => clk, R => n17, S 
                           => n5, Q => present_val_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n48, CLK => clk, R => n17, S 
                           => n4, Q => present_val_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n49, CLK => clk, R => n17, S 
                           => n3, Q => present_val_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n50, CLK => clk, R => n17, S 
                           => n2, Q => present_val_1_port);
   present_val_reg_0_inst : DFFSR port map( D => n43, CLK => clk, R => n17, S 
                           => n1, Q => d_encode_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n12 <= '1';
   U13 : AND2X2 port map( A => n20, B => n16, Y => n11);
   U15 : INVX4 port map( A => n11, Y => n68);
   U16 : INVX4 port map( A => n69, Y => n65);
   U17 : BUFX4 port map( A => n11, Y => n13);
   U18 : BUFX2 port map( A => n69, Y => n14);
   U19 : INVX2 port map( A => rst, Y => n17);
   U20 : INVX4 port map( A => n15, Y => n16);
   U21 : INVX2 port map( A => n62, Y => n15);
   U22 : INVX2 port map( A => t_bitstuff, Y => n18);
   U23 : NAND2X1 port map( A => SHIFT_ENABLE_R, B => n18, Y => n20);
   U24 : NAND2X1 port map( A => count_1_port, B => count_0_port, Y => n64);
   U25 : INVX2 port map( A => n64, Y => n19);
   U26 : NAND3X1 port map( A => SHIFT_ENABLE_R, B => count_2_port, C => n19, Y 
                           => n62);
   U27 : NAND2X1 port map( A => d_encode_port, B => n13, Y => n24);
   U28 : NAND2X1 port map( A => n68, B => n16, Y => n69);
   U29 : NAND2X1 port map( A => present_val_1_port, B => n65, Y => n23);
   U30 : INVX2 port map( A => send_data(0), Y => n21);
   U31 : OR2X2 port map( A => n16, B => n21, Y => n22);
   U32 : NAND3X1 port map( A => n22, B => n23, C => n24, Y => n43);
   U33 : NAND2X1 port map( A => present_val_1_port, B => n13, Y => n28);
   U34 : NAND2X1 port map( A => present_val_2_port, B => n65, Y => n27);
   U35 : INVX2 port map( A => send_data(1), Y => n25);
   U36 : OR2X2 port map( A => n16, B => n25, Y => n26);
   U37 : NAND3X1 port map( A => n28, B => n27, C => n26, Y => n50);
   U38 : NAND2X1 port map( A => present_val_2_port, B => n13, Y => n32);
   U39 : NAND2X1 port map( A => present_val_3_port, B => n65, Y => n31);
   U40 : INVX2 port map( A => send_data(2), Y => n29);
   U41 : OR2X2 port map( A => n16, B => n29, Y => n30);
   U42 : NAND3X1 port map( A => n32, B => n31, C => n30, Y => n49);
   U43 : NAND2X1 port map( A => present_val_3_port, B => n13, Y => n36);
   U44 : NAND2X1 port map( A => present_val_4_port, B => n65, Y => n35);
   U45 : INVX2 port map( A => send_data(3), Y => n33);
   U46 : OR2X2 port map( A => n16, B => n33, Y => n34);
   U47 : NAND3X1 port map( A => n36, B => n35, C => n34, Y => n48);
   U48 : NAND2X1 port map( A => present_val_4_port, B => n13, Y => n40);
   U49 : NAND2X1 port map( A => present_val_5_port, B => n65, Y => n39);
   U50 : INVX2 port map( A => send_data(4), Y => n37);
   U51 : OR2X2 port map( A => n16, B => n37, Y => n38);
   U52 : NAND3X1 port map( A => n40, B => n39, C => n38, Y => n47);
   U53 : NAND2X1 port map( A => present_val_5_port, B => n13, Y => n55);
   U54 : NAND2X1 port map( A => present_val_6_port, B => n65, Y => n54);
   U55 : INVX2 port map( A => send_data(5), Y => n41);
   U56 : OR2X2 port map( A => n16, B => n41, Y => n42);
   U57 : NAND3X1 port map( A => n55, B => n54, C => n42, Y => n46);
   U58 : NAND2X1 port map( A => present_val_6_port, B => n13, Y => n59);
   U59 : NAND2X1 port map( A => present_val_7_port, B => n65, Y => n58);
   U60 : INVX2 port map( A => send_data(6), Y => n56);
   U61 : OR2X2 port map( A => n16, B => n56, Y => n57);
   U62 : NAND3X1 port map( A => n59, B => n58, C => n57, Y => n45);
   U63 : INVX2 port map( A => present_val_7_port, Y => n61);
   U64 : INVX2 port map( A => send_data(7), Y => n60);
   U65 : OAI22X1 port map( A => n68, B => n61, C => n16, D => n60, Y => n44);
   U66 : NAND2X1 port map( A => count_2_port, B => n16, Y => n63);
   U67 : OAI21X1 port map( A => n64, B => n14, C => n63, Y => n52);
   U68 : NAND2X1 port map( A => n65, B => count_0_port, Y => n67);
   U69 : AND2X2 port map( A => count_0_port, B => n68, Y => n66);
   U70 : MUX2X1 port map( B => n67, A => n66, S => count_1_port, Y => n51);
   U71 : MUX2X1 port map( B => n14, A => n68, S => count_0_port, Y => n53);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_encode_1 is

   port( clk, rst, SHIFT_ENABLE_E, d_encode, EOP : in std_logic;  t_bitstuff, 
         dp_tx_out, dm_tx_out : out std_logic);

end tx_encode_1;

architecture SYN_moore of tx_encode_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal DE_holdout, DE_holdout_BS, state_3_port, state_2_port, state_1_port, 
      state_0_port, nextstate_3_port, nextstate_2_port, nextstate_1_port, 
      nextstate_0_port, DE_holdout_last, DE_holdout_nxt, dm_tx_nxt, n9, n12, 
      n13, n14, n15, n18, n19, n20, n26, n27, n32, n37, n39, n40, n41, n43, n44
      , n49, n50, n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n1, n2, n3,
      n4, n5, n6, n7, n8, n10, n11, n16, n17, n21, n22, n23, n24, n25, n28, n29
      , n30, n31, n33, n34, n35, n36, n38, n42, n45, n46, n47, n48, n51, n52, 
      n53, n63, n65, n66, n67 : std_logic;

begin
   
   DE_holdout_reg : DFFSR port map( D => DE_holdout_nxt, CLK => clk, R => n62, 
                           S => n6, Q => DE_holdout);
   DE_holdout_last_reg : DFFPOSX1 port map( D => n61, CLK => clk, Q => 
                           DE_holdout_last);
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => clk, R => 
                           n6, S => n60, Q => state_3_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n6, S => n59, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n6, S => n58, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n6, S => n57, Q => state_2_port);
   DE_holdout_BS_reg : DFFSR port map( D => n64, CLK => clk, R => n6, S => n56,
                           Q => DE_holdout_BS);
   dp_tx_out_reg : DFFSR port map( D => DE_holdout_nxt, CLK => clk, R => n55, S
                           => n6, Q => dp_tx_out);
   dm_tx_out_reg : DFFSR port map( D => dm_tx_nxt, CLK => clk, R => n6, S => 
                           n54, Q => dm_tx_out);
   U9 : OAI21X1 port map( A => state_1_port, B => n9, C => n13, Y => 
                           nextstate_1_port);
   U11 : OAI21X1 port map( A => n3, B => n15, C => n47, Y => n14);
   U12 : NAND3X1 port map( A => SHIFT_ENABLE_E, B => n53, C => n3, Y => n9);
   U14 : OAI21X1 port map( A => n2, B => n47, C => n18, Y => nextstate_0_port);
   U15 : OAI21X1 port map( A => n19, B => n20, C => SHIFT_ENABLE_E, Y => n18);
   U18 : NOR2X1 port map( A => n3, B => n15, Y => n19);
   U19 : NAND3X1 port map( A => d_encode, B => n26, C => n27, Y => n15);
   U20 : XNOR2X1 port map( A => n66, B => n65, Y => n27);
   U22 : NOR2X1 port map( A => n52, B => SHIFT_ENABLE_E, Y => n12);
   U23 : OAI22X1 port map( A => n6, B => n66, C => rst, D => n65, Y => n61);
   U26 : OAI22X1 port map( A => n5, B => n67, C => n65, D => n32, Y => n64);
   U36 : NOR2X1 port map( A => EOP, B => state_3_port, Y => n26);
   U37 : NOR2X1 port map( A => n4, B => n40, Y => n37);
   U38 : AOI22X1 port map( A => n3, B => n41, C => n48, D => n2, Y => n40);
   U40 : XNOR2X1 port map( A => DE_holdout_BS, B => n44, Y => n41);
   U46 : XOR2X1 port map( A => DE_holdout, B => SHIFT_ENABLE_E, Y => n43);
   U47 : XNOR2X1 port map( A => n49, B => n65, Y => n39);
   U49 : NAND2X1 port map( A => SHIFT_ENABLE_E, B => n63, Y => n49);
   U55 : NAND2X1 port map( A => n44, B => n67, Y => n50);
   U57 : NAND2X1 port map( A => SHIFT_ENABLE_E, B => d_encode, Y => n44);
   n54 <= '1';
   n55 <= '1';
   n56 <= '1';
   n57 <= '1';
   n58 <= '1';
   n59 <= '1';
   n60 <= '1';
   n62 <= '1';
   U3 : INVX1 port map( A => n2, Y => n3);
   U4 : INVX2 port map( A => state_0_port, Y => n2);
   U5 : AND2X2 port map( A => n27, B => d_encode, Y => n1);
   U6 : AND2X2 port map( A => n1, B => n26, Y => n53);
   U7 : INVX2 port map( A => n51, Y => n4);
   U8 : INVX1 port map( A => EOP, Y => n51);
   U10 : INVX2 port map( A => rst, Y => n6);
   U13 : NOR2X1 port map( A => n42, B => n8, Y => n5);
   U16 : INVX1 port map( A => n5, Y => n32);
   U17 : NAND2X1 port map( A => state_2_port, B => state_1_port, Y => n7);
   U21 : NOR3X1 port map( A => state_3_port, B => n7, C => n2, Y => t_bitstuff)
                           ;
   U24 : INVX2 port map( A => n7, Y => n25);
   U25 : NAND3X1 port map( A => n26, B => n2, C => n25, Y => n42);
   U27 : INVX2 port map( A => SHIFT_ENABLE_E, Y => n8);
   U28 : NAND2X1 port map( A => n63, B => n25, Y => n10);
   U29 : OAI21X1 port map( A => n52, B => n10, C => n42, Y => n20);
   U30 : INVX2 port map( A => n42, Y => n11);
   U31 : AOI21X1 port map( A => n14, B => state_1_port, C => n11, Y => n13);
   U32 : INVX2 port map( A => state_2_port, Y => n16);
   U33 : INVX2 port map( A => state_1_port, Y => n33);
   U34 : NAND3X1 port map( A => n2, B => n16, C => n33, Y => n45);
   U35 : NAND2X1 port map( A => n45, B => state_3_port, Y => n31);
   U39 : INVX2 port map( A => n39, Y => n17);
   U41 : NOR2X1 port map( A => n52, B => n17, Y => n21);
   U42 : MUX2X1 port map( B => n21, A => n37, S => n25, Y => n22);
   U43 : NAND2X1 port map( A => n31, B => n22, Y => dm_tx_nxt);
   U44 : OAI21X1 port map( A => n67, B => n44, C => n50, Y => n24);
   U45 : AND2X2 port map( A => n43, B => n2, Y => n23);
   U48 : AOI21X1 port map( A => n3, B => n24, C => n23, Y => n28);
   U50 : MUX2X1 port map( B => n39, A => n28, S => n25, Y => n29);
   U51 : OAI21X1 port map( A => state_3_port, B => n29, C => n51, Y => n30);
   U52 : NAND2X1 port map( A => n31, B => n30, Y => DE_holdout_nxt);
   U53 : NAND2X1 port map( A => n46, B => state_1_port, Y => n35);
   U54 : AOI21X1 port map( A => n53, B => n33, C => n12, Y => n34);
   U56 : MUX2X1 port map( B => n35, A => n34, S => state_2_port, Y => n36);
   U58 : INVX2 port map( A => n36, Y => n38);
   U59 : NAND2X1 port map( A => n42, B => n38, Y => nextstate_2_port);
   U60 : AOI21X1 port map( A => state_3_port, B => n45, C => n51, Y => 
                           nextstate_3_port);
   U61 : INVX2 port map( A => n9, Y => n46);
   U62 : INVX2 port map( A => n12, Y => n47);
   U63 : INVX2 port map( A => n43, Y => n48);
   U64 : INVX2 port map( A => n26, Y => n52);
   U65 : INVX2 port map( A => d_encode, Y => n63);
   U74 : INVX2 port map( A => DE_holdout, Y => n65);
   U75 : INVX2 port map( A => DE_holdout_last, Y => n66);
   U76 : INVX2 port map( A => DE_holdout_BS, Y => n67);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_CRC_CALC_1 is

   port( CLK, RST, EOP, T_STROBE : in std_logic;  PRGA_OPCODE : in 
         std_logic_vector (1 downto 0);  PRGA_OUT : in std_logic_vector (7 
         downto 0);  TX_CRC : out std_logic_vector (15 downto 0));

end tx_CRC_CALC_1;

architecture SYN_txcrcm of tx_CRC_CALC_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal TX_CRC_15_port, TX_CRC_14_port, TX_CRC_13_port, TX_CRC_12_port, 
      TX_CRC_11_port, TX_CRC_10_port, TX_CRC_9_port, TX_CRC_8_port, 
      TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port, TX_CRC_4_port, TX_CRC_3_port
      , TX_CRC_2_port, TX_CRC_1_port, TX_CRC_0_port, n1, n2, n4, n6, n8, n10, 
      n12, n14, n15, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n3, n5, n7, n9, n11, n13, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n79, n80
      : std_logic;

begin
   TX_CRC <= ( TX_CRC_15_port, TX_CRC_14_port, TX_CRC_13_port, TX_CRC_12_port, 
      TX_CRC_11_port, TX_CRC_10_port, TX_CRC_9_port, TX_CRC_8_port, 
      TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port, TX_CRC_4_port, TX_CRC_3_port
      , TX_CRC_2_port, TX_CRC_1_port, TX_CRC_0_port );
   
   current_crc_reg_8_inst : DFFSR port map( D => n70, CLK => CLK, R => n21, S 
                           => n15, Q => TX_CRC_8_port);
   current_crc_reg_15_inst : DFFSR port map( D => n63, CLK => CLK, R => n21, S 
                           => n14, Q => TX_CRC_15_port);
   current_crc_reg_9_inst : DFFSR port map( D => n69, CLK => CLK, R => n21, S 
                           => n12, Q => TX_CRC_9_port);
   current_crc_reg_10_inst : DFFSR port map( D => n68, CLK => CLK, R => n21, S 
                           => n10, Q => TX_CRC_10_port);
   current_crc_reg_11_inst : DFFSR port map( D => n67, CLK => CLK, R => n21, S 
                           => n8, Q => TX_CRC_11_port);
   current_crc_reg_12_inst : DFFSR port map( D => n66, CLK => CLK, R => n21, S 
                           => n6, Q => TX_CRC_12_port);
   current_crc_reg_13_inst : DFFSR port map( D => n65, CLK => CLK, R => n21, S 
                           => n4, Q => TX_CRC_13_port);
   current_crc_reg_14_inst : DFFSR port map( D => n64, CLK => CLK, R => n21, S 
                           => n2, Q => TX_CRC_14_port);
   current_crc_reg_7_inst : DFFSR port map( D => n71, CLK => CLK, R => n21, S 
                           => n1, Q => TX_CRC_7_port);
   n1 <= '1';
   n2 <= '1';
   n4 <= '1';
   n6 <= '1';
   n8 <= '1';
   n10 <= '1';
   n12 <= '1';
   n14 <= '1';
   n15 <= '1';
   U39 : OAI22X1 port map( A => n25, B => n20, C => n38, D => n19, Y => n63);
   U40 : XNOR2X1 port map( A => n40, B => n79, Y => n38);
   U41 : OAI22X1 port map( A => n37, B => n20, C => n19, D => n36, Y => n64);
   U42 : OAI22X1 port map( A => n35, B => n20, C => n19, D => n34, Y => n65);
   U43 : OAI22X1 port map( A => n33, B => n20, C => n19, D => n32, Y => n66);
   U44 : OAI22X1 port map( A => n31, B => n20, C => n19, D => n30, Y => n67);
   U45 : OAI22X1 port map( A => n29, B => n20, C => n19, D => n28, Y => n68);
   U46 : OAI22X1 port map( A => n27, B => n20, C => n41, D => n19, Y => n69);
   U47 : XNOR2X1 port map( A => TX_CRC_1_port, B => n42, Y => n41);
   U48 : OAI22X1 port map( A => n24, B => n20, C => n43, D => n19, Y => n70);
   U49 : XOR2X1 port map( A => n44, B => n45, Y => n43);
   U50 : XNOR2X1 port map( A => TX_CRC_0_port, B => n42, Y => n44);
   U51 : OAI22X1 port map( A => n79, B => n20, C => n46, D => n19, Y => n71);
   U52 : OAI22X1 port map( A => n20, B => n36, C => n47, D => n19, Y => n72);
   U53 : XNOR2X1 port map( A => n48, B => n49, Y => n47);
   U54 : OAI22X1 port map( A => n20, B => n34, C => n50, D => n19, Y => n73);
   U55 : OAI22X1 port map( A => n20, B => n32, C => n51, D => n19, Y => n74);
   U56 : XNOR2X1 port map( A => n52, B => n53, Y => n51);
   U57 : OAI22X1 port map( A => n20, B => n30, C => n54, D => n19, Y => n75);
   U58 : OAI22X1 port map( A => n20, B => n28, C => n55, D => n19, Y => n76);
   U59 : XOR2X1 port map( A => n56, B => n57, Y => n55);
   U60 : OAI22X1 port map( A => n20, B => n26, C => n58, D => n19, Y => n77);
   U61 : XOR2X1 port map( A => n59, B => n60, Y => n58);
   U62 : XOR2X1 port map( A => n42, B => n46, Y => n59);
   U63 : OAI22X1 port map( A => n20, B => n23, C => n40, D => n19, Y => n78);
   U64 : XOR2X1 port map( A => n61, B => n62, Y => n40);
   U65 : XOR2X1 port map( A => n57, B => n42, Y => n62);
   U66 : XNOR2X1 port map( A => n25, B => PRGA_OUT(7), Y => n42);
   U67 : XNOR2X1 port map( A => n24, B => PRGA_OUT(0), Y => n57);
   U68 : XOR2X1 port map( A => n46, B => n60, Y => n61);
   U69 : XOR2X1 port map( A => n54, B => n50, Y => n60);
   U70 : XNOR2X1 port map( A => n53, B => n48, Y => n50);
   U71 : XOR2X1 port map( A => TX_CRC_12_port, B => PRGA_OUT(4), Y => n48);
   U72 : XOR2X1 port map( A => TX_CRC_11_port, B => PRGA_OUT(3), Y => n53);
   U74 : XOR2X1 port map( A => TX_CRC_10_port, B => PRGA_OUT(2), Y => n52);
   U75 : XNOR2X1 port map( A => TX_CRC_9_port, B => PRGA_OUT(1), Y => n56);
   U76 : XNOR2X1 port map( A => n49, B => n45, Y => n46);
   U77 : XNOR2X1 port map( A => n37, B => PRGA_OUT(6), Y => n45);
   U78 : XOR2X1 port map( A => TX_CRC_13_port, B => PRGA_OUT(5), Y => n49);
   U80 : NAND3X1 port map( A => PRGA_OPCODE(0), B => n80, C => T_STROBE, Y => 
                           n39);
   current_crc_reg_6_inst : DFFSR port map( D => n72, CLK => CLK, R => n21, S 
                           => n16, Q => TX_CRC_6_port);
   current_crc_reg_5_inst : DFFSR port map( D => n73, CLK => CLK, R => n21, S 
                           => n13, Q => TX_CRC_5_port);
   current_crc_reg_4_inst : DFFSR port map( D => n74, CLK => CLK, R => n21, S 
                           => n11, Q => TX_CRC_4_port);
   current_crc_reg_3_inst : DFFSR port map( D => n75, CLK => CLK, R => n21, S 
                           => n9, Q => TX_CRC_3_port);
   current_crc_reg_2_inst : DFFSR port map( D => n76, CLK => CLK, R => n21, S 
                           => n7, Q => TX_CRC_2_port);
   current_crc_reg_1_inst : DFFSR port map( D => n77, CLK => CLK, R => n21, S 
                           => n5, Q => TX_CRC_1_port);
   current_crc_reg_0_inst : DFFSR port map( D => n78, CLK => CLK, R => n21, S 
                           => n3, Q => TX_CRC_0_port);
   U5 : INVX4 port map( A => n17, Y => n20);
   n3 <= '1';
   n5 <= '1';
   n7 <= '1';
   n9 <= '1';
   n11 <= '1';
   n13 <= '1';
   n16 <= '1';
   U20 : INVX1 port map( A => EOP, Y => n22);
   U21 : INVX2 port map( A => n39, Y => n18);
   U22 : AND2X2 port map( A => n39, B => n22, Y => n17);
   U23 : INVX2 port map( A => RST, Y => n21);
   U24 : XOR2X1 port map( A => n56, B => n52, Y => n54);
   U25 : INVX2 port map( A => n18, Y => n19);
   U26 : INVX2 port map( A => TX_CRC_0_port, Y => n23);
   U27 : INVX2 port map( A => TX_CRC_8_port, Y => n24);
   U28 : INVX2 port map( A => TX_CRC_15_port, Y => n25);
   U29 : INVX2 port map( A => TX_CRC_1_port, Y => n26);
   U30 : INVX2 port map( A => TX_CRC_9_port, Y => n27);
   U31 : INVX2 port map( A => TX_CRC_2_port, Y => n28);
   U32 : INVX2 port map( A => TX_CRC_10_port, Y => n29);
   U33 : INVX2 port map( A => TX_CRC_3_port, Y => n30);
   U34 : INVX2 port map( A => TX_CRC_11_port, Y => n31);
   U35 : INVX2 port map( A => TX_CRC_4_port, Y => n32);
   U36 : INVX2 port map( A => TX_CRC_12_port, Y => n33);
   U37 : INVX2 port map( A => TX_CRC_5_port, Y => n34);
   U38 : INVX2 port map( A => TX_CRC_13_port, Y => n35);
   U73 : INVX2 port map( A => TX_CRC_6_port, Y => n36);
   U79 : INVX2 port map( A => TX_CRC_14_port, Y => n37);
   U81 : INVX2 port map( A => TX_CRC_7_port, Y => n79);
   U82 : INVX2 port map( A => PRGA_OPCODE(1), Y => n80);

end SYN_txcrcm;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_timer_1 is

   port( CLK, RST, D_EDGE, RCVING : in std_logic;  SHIFT_ENABLE : out std_logic
         );

end rx_timer_1;

architecture SYN_moore of rx_timer_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal count_3_port, count_2_port, count_1_port, count_0_port, state, 
      nextcount_3_port, nextcount_2_port, nextcount_1_port, nextcount_0_port, 
      n1, n2, n3, n4, n6, n15, n17, n18, n20, n21, n22, n23, n5, n7, n8, n9, 
      n10, n11, n12, n13, n14, n16, n19, n24, n25, n26, n27 : std_logic;

begin
   
   state_reg : DFFSR port map( D => n11, CLK => CLK, R => n12, S => n6, Q => 
                           state);
   count_reg_0_inst : DFFSR port map( D => nextcount_0_port, CLK => CLK, R => 
                           n12, S => n4, Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => nextcount_1_port, CLK => CLK, R => 
                           n12, S => n3, Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => nextcount_2_port, CLK => CLK, R => 
                           n12, S => n2, Q => count_2_port);
   count_reg_3_inst : DFFSR port map( D => nextcount_3_port, CLK => CLK, R => 
                           n12, S => n1, Q => count_3_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n6 <= '1';
   U19 : XOR2X1 port map( A => n18, B => n25, Y => n17);
   U20 : NOR2X1 port map( A => count_3_port, B => n26, Y => n15);
   U22 : XOR2X1 port map( A => n21, B => count_2_port, Y => n20);
   U24 : NAND2X1 port map( A => state, B => n23, Y => nextcount_0_port);
   U25 : OAI21X1 port map( A => D_EDGE, B => n27, C => n11, Y => n23);
   U30 : NAND2X1 port map( A => count_0_port, B => count_1_port, Y => n21);
   U32 : XNOR2X1 port map( A => count_0_port, B => count_1_port, Y => n22);
   U7 : INVX2 port map( A => n10, Y => SHIFT_ENABLE);
   U9 : INVX1 port map( A => n7, Y => nextcount_2_port);
   U10 : INVX2 port map( A => RST, Y => n12);
   U11 : NOR2X1 port map( A => n16, B => n25, Y => n5);
   U12 : OAI21X1 port map( A => n8, B => D_EDGE, C => n11, Y => n7);
   U13 : NAND2X1 port map( A => n20, B => state, Y => n8);
   U14 : NOR2X1 port map( A => D_EDGE, B => n14, Y => n9);
   U15 : NAND2X1 port map( A => n5, B => RCVING, Y => n10);
   U16 : BUFX2 port map( A => RCVING, Y => n11);
   U17 : INVX2 port map( A => count_2_port, Y => n13);
   U18 : OAI21X1 port map( A => n22, B => n13, C => n21, Y => n18);
   U21 : XOR2X1 port map( A => n13, B => n22, Y => n25);
   U23 : INVX2 port map( A => state, Y => n14);
   U26 : INVX2 port map( A => n18, Y => n26);
   U27 : NAND3X1 port map( A => count_3_port, B => n9, C => n26, Y => n16);
   U28 : AOI22X1 port map( A => n15, B => n25, C => n17, D => count_3_port, Y 
                           => n19);
   U29 : NAND2X1 port map( A => n11, B => n9, Y => n24);
   U31 : NOR2X1 port map( A => n19, B => n24, Y => nextcount_3_port);
   U33 : NOR2X1 port map( A => n22, B => n24, Y => nextcount_1_port);
   U34 : INVX2 port map( A => count_0_port, Y => n27);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_shift_reg_1 is

   port( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF : in std_logic;  RCV_DATA : 
         out std_logic_vector (7 downto 0));

end rx_shift_reg_1;

architecture SYN_dataflow of rx_shift_reg_1 is

   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      present_val_7_port, present_val_6_port, present_val_5_port, 
      present_val_4_port, present_val_3_port, present_val_2_port, 
      present_val_1_port, present_val_0_port, n2, n6, n8, n10, n12, n14, n16, 
      n18, n21, n23, n24, n26, n27, n29, n30, n32, n33, n35, n36, n38, n39, n41
      , n42, n44, n1, n3, n4, n5, n7, n9, n11, n13, n15, n17, n19, n20, n22, 
      n25, n28, n31, n34, n37, n40, n43, n45, n46, n47, n48, n49, n50 : 
      std_logic;

begin
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   RCV_DATA_reg_7_inst : DFFPOSX1 port map( D => n42, CLK => CLK, Q => 
                           RCV_DATA_7_port);
   RCV_DATA_reg_6_inst : DFFPOSX1 port map( D => n39, CLK => CLK, Q => 
                           RCV_DATA_6_port);
   RCV_DATA_reg_5_inst : DFFPOSX1 port map( D => n36, CLK => CLK, Q => 
                           RCV_DATA_5_port);
   RCV_DATA_reg_4_inst : DFFPOSX1 port map( D => n33, CLK => CLK, Q => 
                           RCV_DATA_4_port);
   RCV_DATA_reg_3_inst : DFFPOSX1 port map( D => n30, CLK => CLK, Q => 
                           RCV_DATA_3_port);
   RCV_DATA_reg_2_inst : DFFPOSX1 port map( D => n27, CLK => CLK, Q => 
                           RCV_DATA_2_port);
   RCV_DATA_reg_1_inst : DFFPOSX1 port map( D => n24, CLK => CLK, Q => 
                           RCV_DATA_1_port);
   RCV_DATA_reg_0_inst : DFFPOSX1 port map( D => n21, CLK => CLK, Q => 
                           RCV_DATA_0_port);
   U2 : OAI21X1 port map( A => RST, B => n50, C => n2, Y => n21);
   U3 : NAND2X1 port map( A => RCV_DATA_0_port, B => RST, Y => n2);
   U6 : OAI21X1 port map( A => RST, B => n49, C => n6, Y => n24);
   U7 : NAND2X1 port map( A => RCV_DATA_1_port, B => RST, Y => n6);
   U10 : OAI21X1 port map( A => RST, B => n48, C => n8, Y => n27);
   U11 : NAND2X1 port map( A => n25, B => RST, Y => n8);
   U14 : OAI21X1 port map( A => RST, B => n47, C => n10, Y => n30);
   U15 : NAND2X1 port map( A => RCV_DATA_3_port, B => RST, Y => n10);
   U18 : OAI21X1 port map( A => RST, B => n46, C => n12, Y => n33);
   U19 : NAND2X1 port map( A => RCV_DATA_4_port, B => RST, Y => n12);
   U22 : OAI21X1 port map( A => RST, B => n45, C => n14, Y => n36);
   U23 : NAND2X1 port map( A => RCV_DATA_5_port, B => RST, Y => n14);
   U26 : OAI21X1 port map( A => RST, B => n43, C => n16, Y => n39);
   U27 : NAND2X1 port map( A => n17, B => RST, Y => n16);
   U30 : OAI21X1 port map( A => RST, B => n40, C => n18, Y => n42);
   U31 : NAND2X1 port map( A => n20, B => RST, Y => n18);
   present_val_reg_0_inst : DFFSR port map( D => n23, CLK => CLK, R => n31, S 
                           => n13, Q => present_val_0_port);
   present_val_reg_7_inst : DFFSR port map( D => n44, CLK => CLK, R => n31, S 
                           => n11, Q => present_val_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n41, CLK => CLK, R => n31, S 
                           => n9, Q => present_val_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n38, CLK => CLK, R => n31, S 
                           => n7, Q => present_val_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n35, CLK => CLK, R => n31, S 
                           => n5, Q => present_val_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n32, CLK => CLK, R => n31, S 
                           => n4, Q => present_val_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n29, CLK => CLK, R => n31, S 
                           => n3, Q => present_val_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n26, CLK => CLK, R => n31, S 
                           => n1, Q => present_val_1_port);
   n1 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n7 <= '1';
   n9 <= '1';
   n11 <= '1';
   n13 <= '1';
   U20 : INVX1 port map( A => RCV_DATA_6_port, Y => n15);
   U21 : INVX2 port map( A => n15, Y => n17);
   U24 : INVX1 port map( A => RCV_DATA_7_port, Y => n19);
   U25 : INVX2 port map( A => n19, Y => n20);
   U28 : INVX1 port map( A => RCV_DATA_2_port, Y => n22);
   U29 : INVX2 port map( A => n22, Y => n25);
   U32 : INVX2 port map( A => RST, Y => n31);
   U33 : AND2X2 port map( A => SHIFT_ENABLE, B => n34, Y => n28);
   U34 : INVX2 port map( A => present_val_7_port, Y => n40);
   U35 : INVX2 port map( A => present_val_6_port, Y => n43);
   U36 : INVX2 port map( A => present_val_5_port, Y => n45);
   U37 : INVX2 port map( A => present_val_4_port, Y => n46);
   U38 : INVX2 port map( A => present_val_3_port, Y => n47);
   U39 : INVX2 port map( A => present_val_2_port, Y => n48);
   U40 : INVX2 port map( A => present_val_1_port, Y => n49);
   U41 : INVX2 port map( A => present_val_0_port, Y => n50);
   U42 : INVX2 port map( A => BITSTUFF, Y => n34);
   U43 : MUX2X1 port map( B => n50, A => n49, S => n28, Y => n23);
   U44 : MUX2X1 port map( B => n49, A => n48, S => n28, Y => n26);
   U45 : MUX2X1 port map( B => n48, A => n47, S => n28, Y => n29);
   U46 : MUX2X1 port map( B => n47, A => n46, S => n28, Y => n32);
   U47 : MUX2X1 port map( B => n46, A => n45, S => n28, Y => n35);
   U48 : MUX2X1 port map( B => n45, A => n43, S => n28, Y => n38);
   U49 : MUX2X1 port map( B => n43, A => n40, S => n28, Y => n41);
   U50 : INVX2 port map( A => D_ORIG, Y => n37);
   U51 : MUX2X1 port map( B => n40, A => n37, S => n28, Y => n44);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_rcu_1 is

   port( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR : in std_logic
         ;  RX_CRC, RX_CHECK_CRC : in std_logic_vector (15 downto 0);  RCV_DATA
         : in std_logic_vector (7 downto 0);  RCVING, W_ENABLE, R_ERROR, 
         CRC_ERROR : out std_logic;  OPCODE : out std_logic_vector (1 downto 0)
         );

end rx_rcu_1;

architecture SYN_moore of rx_rcu_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal CRC_ERROR_port, state_3_port, state_2_port, state_1_port, 
      state_0_port, count_3_port, count_2_port, count_1_port, count_0_port, 
      nextstate_3_port, nextstate_2_port, nextstate_1_port, nextstate_0_port, 
      nxtR_ERROR, curR_ERROR, curCRC_ERROR, N170, n37, n38, n41, n42, n83, n87,
      n88, n94, n149, n150, n151, n152, n155, n156, n158, n159, n161, n162, 
      n163, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31
      , n32, n33, n34, n35, n36, n39, n40, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n84, n85, n86, n89, n90, n91, n92, n93, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n153, n154, n157, n160, n164, n165, n166, n167, n168, 
      n169, n170_port, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223 : std_logic;

begin
   CRC_ERROR <= CRC_ERROR_port;
   
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => CLK, R => 
                           n51, S => n159, Q => state_3_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => CLK, R => 
                           n51, S => n158, Q => state_0_port);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => CLK, R => 
                           n51, S => n156, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => CLK, R => 
                           n51, S => n155, Q => state_1_port);
   count_reg_3_inst : DFFSR port map( D => n163, CLK => CLK, R => n51, S => 
                           n152, Q => count_3_port);
   curCRC_ERROR_reg : DFFPOSX1 port map( D => n151, CLK => CLK, Q => 
                           curCRC_ERROR);
   curR_ERROR_reg : DFFPOSX1 port map( D => n150, CLK => CLK, Q => curR_ERROR);
   R_ERROR_reg : DFFSR port map( D => nxtR_ERROR, CLK => CLK, R => n51, S => 
                           n149, Q => R_ERROR);
   CRC_ERROR_reg : DFFPOSX1 port map( D => n218, CLK => CLK, Q => 
                           CRC_ERROR_port);
   U16 : NAND2X1 port map( A => n37, B => n38, Y => nextstate_2_port);
   U19 : OAI21X1 port map( A => n222, B => n42, C => n47, Y => n41);
   U20 : NAND2X1 port map( A => n184, B => n185, Y => n42);
   U52 : AOI21X1 port map( A => CRC_ERROR_port, B => RST, C => n88, Y => n87);
   U56 : OAI21X1 port map( A => n51, B => n220, C => n94, Y => n150);
   U79 : NOR2X1 port map( A => D_EDGE, B => n49, Y => n83);
   n149 <= '1';
   n152 <= '1';
   n155 <= '1';
   n156 <= '1';
   n158 <= '1';
   n159 <= '1';
   count_reg_0_inst : DFFSR port map( D => n217, CLK => CLK, R => n51, S => n13
                           , Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => n161, CLK => CLK, R => n51, S => n12
                           , Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n162, CLK => CLK, R => n51, S => n11
                           , Q => count_2_port);
   U3 : AND2X2 port map( A => n5, B => n48, Y => n1);
   U4 : AND2X1 port map( A => n65, B => n129, Y => n2);
   U5 : BUFX2 port map( A => n39, Y => n3);
   U6 : BUFX2 port map( A => n35, Y => n4);
   U7 : BUFX4 port map( A => state_1_port, Y => n5);
   U8 : AND2X2 port map( A => n168, B => n85, Y => n6);
   U9 : AND2X2 port map( A => n19, B => n35, Y => n7);
   U10 : AND2X2 port map( A => n50, B => n166, Y => n8);
   U11 : INVX2 port map( A => n14, Y => n170_port);
   U12 : AND2X1 port map( A => n70, B => n16, Y => n9);
   U13 : AND2X2 port map( A => n21, B => n7, Y => n10);
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   U18 : INVX2 port map( A => n48, Y => n14);
   U21 : INVX4 port map( A => n48, Y => n49);
   U22 : NAND2X1 port map( A => n5, B => n170_port, Y => n15);
   U23 : BUFX2 port map( A => n129, Y => n16);
   U24 : BUFX2 port map( A => n5, Y => n47);
   U25 : BUFX2 port map( A => n46, Y => n17);
   U26 : AND2X2 port map( A => n5, B => n14, Y => n52);
   U27 : BUFX2 port map( A => n33, Y => n18);
   U28 : NAND2X1 port map( A => n32, B => n2, Y => W_ENABLE);
   U29 : AND2X2 port map( A => n64, B => n63, Y => n19);
   U30 : INVX1 port map( A => n19, Y => n135);
   U31 : INVX1 port map( A => n54, Y => n20);
   U32 : BUFX2 port map( A => n1, Y => n21);
   U33 : INVX4 port map( A => n50, Y => n54);
   U34 : NAND2X1 port map( A => n21, B => n8, Y => n22);
   U35 : NAND2X1 port map( A => n1, B => n8, Y => n123);
   U36 : NAND2X1 port map( A => n24, B => n9, Y => RCVING);
   U37 : INVX2 port map( A => n175, Y => n23);
   U38 : AND2X2 port map( A => n25, B => n43, Y => n24);
   U39 : INVX1 port map( A => n24, Y => n90);
   U40 : NOR2X1 port map( A => n36, B => n23, Y => n25);
   U41 : NAND2X1 port map( A => n1, B => n7, Y => n179);
   U42 : AND2X2 port map( A => SHIFT_ENABLE, B => n103, Y => n26);
   U43 : AND2X1 port map( A => n111, B => n115, Y => n112);
   U44 : BUFX4 port map( A => state_3_port, Y => n39);
   U45 : AND2X1 port map( A => n46, B => n54, Y => n27);
   U46 : INVX1 port map( A => n47, Y => n73);
   U47 : INVX2 port map( A => n125, Y => n28);
   U48 : AND2X2 port map( A => n39, B => n50, Y => n29);
   U49 : INVX1 port map( A => n29, Y => n153);
   U50 : NAND2X1 port map( A => n65, B => n129, Y => OPCODE(0));
   U51 : AND2X1 port map( A => n118, B => n115, Y => n31);
   U53 : OR2X1 port map( A => RCV_DATA(1), B => RCV_DATA(2), Y => n60);
   U54 : AND2X2 port map( A => n68, B => n179, Y => n32);
   U55 : INVX2 port map( A => RST, Y => n51);
   U57 : AND2X2 port map( A => n39, B => n54, Y => n33);
   U58 : AND2X2 port map( A => SHIFT_ENABLE, B => n103, Y => n34);
   U59 : NOR2X1 port map( A => n50, B => n39, Y => n35);
   U60 : NAND2X1 port map( A => n69, B => n68, Y => n36);
   U61 : INVX1 port map( A => n111, Y => n107);
   U62 : INVX1 port map( A => n105, Y => n110);
   U63 : INVX1 port map( A => n67, Y => n40);
   U64 : INVX1 port map( A => n40, Y => n43);
   U65 : INVX2 port map( A => n71, Y => n44);
   U66 : INVX1 port map( A => n8, Y => n45);
   U67 : AND2X2 port map( A => state_2_port, B => n166, Y => n46);
   U68 : INVX1 port map( A => n17, Y => n71);
   U69 : BUFX4 port map( A => state_0_port, Y => n50);
   U70 : INVX1 port map( A => n178, Y => n125);
   U71 : INVX2 port map( A => state_2_port, Y => n48);
   U72 : INVX1 port map( A => n167, Y => n168);
   U73 : INVX2 port map( A => state_3_port, Y => n166);
   U74 : NAND2X1 port map( A => n52, B => n8, Y => n129);
   U75 : NAND2X1 port map( A => n17, B => n54, Y => n167);
   U76 : NAND2X1 port map( A => n27, B => n47, Y => n65);
   U77 : INVX2 port map( A => n5, Y => n172);
   U78 : NOR2X1 port map( A => n49, B => n172, Y => n53);
   U80 : NAND2X1 port map( A => n53, B => n29, Y => n178);
   U81 : NAND2X1 port map( A => n178, B => n123, Y => n89);
   U82 : INVX2 port map( A => n89, Y => n67);
   U83 : NAND2X1 port map( A => n33, B => n49, Y => n56);
   U84 : OAI21X1 port map( A => n50, B => n170_port, C => n166, Y => n55);
   U85 : MUX2X1 port map( B => n56, A => n55, S => n47, Y => n57);
   U86 : NAND2X1 port map( A => n57, B => n67, Y => OPCODE(1));
   U87 : NAND3X1 port map( A => n33, B => n49, C => n172, Y => n68);
   U88 : INVX2 port map( A => RCV_DATA(0), Y => n58);
   U89 : NAND2X1 port map( A => RCV_DATA(7), B => n58, Y => n59);
   U90 : NOR2X1 port map( A => n60, B => n59, Y => n64);
   U91 : NOR2X1 port map( A => RCV_DATA(4), B => RCV_DATA(3), Y => n62);
   U92 : NOR2X1 port map( A => RCV_DATA(6), B => RCV_DATA(5), Y => n61);
   U93 : AND2X2 port map( A => n62, B => n61, Y => n63);
   U94 : NAND3X1 port map( A => n29, B => n49, C => n172, Y => n177);
   U95 : OAI21X1 port map( A => n47, B => n167, C => n177, Y => n121);
   U96 : INVX2 port map( A => n121, Y => n70);
   U97 : NOR2X1 port map( A => n39, B => n49, Y => n66);
   U98 : NAND3X1 port map( A => n66, B => n50, C => n172, Y => n175);
   U99 : NAND2X1 port map( A => n43, B => n175, Y => n104);
   U100 : NAND2X1 port map( A => n1, B => n166, Y => n69);
   U101 : NAND2X1 port map( A => n83, B => n18, Y => n81);
   U102 : NAND2X1 port map( A => n81, B => n71, Y => n72);
   U103 : NAND3X1 port map( A => curR_ERROR, B => n73, C => n72, Y => n79);
   U104 : NOR2X1 port map( A => n20, B => n15, Y => n75);
   U105 : NAND2X1 port map( A => n19, B => n166, Y => n74);
   U106 : NAND2X1 port map( A => n75, B => n74, Y => n96);
   U107 : NAND2X1 port map( A => n28, B => n175, Y => n77);
   U108 : NOR2X1 port map( A => count_3_port, B => n172, Y => n76);
   U109 : NOR3X1 port map( A => count_0_port, B => count_1_port, C => 
                           count_2_port, Y => n184);
   U110 : NAND2X1 port map( A => n76, B => n184, Y => n84);
   U111 : AOI22X1 port map( A => EOP, B => n77, C => n168, D => n84, Y => n78);
   U112 : NAND3X1 port map( A => n79, B => n96, C => n78, Y => nxtR_ERROR);
   U113 : INVX2 port map( A => n79, Y => n80);
   U114 : OAI21X1 port map( A => n51, B => n80, C => nxtR_ERROR, Y => n94);
   U115 : NAND2X1 port map( A => curCRC_ERROR, B => n51, Y => n86);
   U116 : NAND2X1 port map( A => n8, B => n49, Y => n91);
   U117 : NAND2X1 port map( A => n91, B => n81, Y => n82);
   U118 : NAND2X1 port map( A => n82, B => n172, Y => n99);
   U119 : INVX2 port map( A => n84, Y => n85);
   U120 : NAND3X1 port map( A => n222, B => n51, C => n6, Y => n102);
   U121 : OAI21X1 port map( A => n86, B => n99, C => n102, Y => n88);
   U122 : INVX2 port map( A => count_3_port, Y => n185);
   U123 : NAND2X1 port map( A => n184, B => count_3_port, Y => n124);
   U124 : INVX2 port map( A => n124, Y => n122);
   U125 : AOI22X1 port map( A => n90, B => BS_ERROR, C => n122, D => n89, Y => 
                           n95);
   U126 : OAI22X1 port map( A => n167, B => EOP, C => D_EDGE, D => n91, Y => 
                           n92);
   U127 : MUX2X1 port map( B => n92, A => n18, S => n47, Y => n93);
   U128 : AND2X2 port map( A => n95, B => n93, Y => n37);
   U129 : OAI21X1 port map( A => n41, B => n167, C => n96, Y => n98);
   U130 : NAND2X1 port map( A => EOP, B => n104, Y => n115);
   U131 : NAND2X1 port map( A => n115, B => n177, Y => n97);
   U132 : NOR2X1 port map( A => n98, B => n97, Y => n38);
   U133 : INVX2 port map( A => n99, Y => n100);
   U134 : OAI21X1 port map( A => RST, B => n100, C => curCRC_ERROR, Y => n101);
   U135 : NAND2X1 port map( A => n102, B => n101, Y => n151);
   U136 : INVX2 port map( A => BITSTUFF, Y => n103);
   U137 : NAND3X1 port map( A => count_1_port, B => count_0_port, C => n34, Y 
                           => n105);
   U138 : NAND2X1 port map( A => n104, B => n124, Y => n116);
   U139 : INVX2 port map( A => n116, Y => n118);
   U140 : NAND3X1 port map( A => n110, B => n31, C => count_2_port, Y => n109);
   U141 : NAND2X1 port map( A => n118, B => n105, Y => n111);
   U142 : OAI21X1 port map( A => count_2_port, B => n116, C => n115, Y => n106)
                           ;
   U143 : NOR2X1 port map( A => n107, B => n106, Y => n108);
   U144 : MUX2X1 port map( B => n109, A => n108, S => count_3_port, Y => n163);
   U145 : NAND2X1 port map( A => n31, B => n110, Y => n113);
   U146 : MUX2X1 port map( B => n113, A => n112, S => count_2_port, Y => n162);
   U147 : NAND3X1 port map( A => n26, B => n118, C => n115, Y => n134);
   U148 : INVX2 port map( A => n134, Y => n114);
   U149 : NAND2X1 port map( A => count_0_port, B => n114, Y => n120);
   U150 : INVX2 port map( A => count_0_port, Y => n117);
   U151 : OAI21X1 port map( A => n26, B => n116, C => n115, Y => n132);
   U152 : AOI21X1 port map( A => n118, B => n117, C => n132, Y => n119);
   U153 : MUX2X1 port map( B => n120, A => n119, S => count_1_port, Y => n161);
   U154 : NAND2X1 port map( A => n121, B => EOP, Y => n131);
   U155 : NAND2X1 port map( A => n122, B => n223, Y => n140);
   U156 : OAI21X1 port map( A => n140, B => n175, C => n22, Y => n128);
   U157 : NAND3X1 port map( A => n223, B => n125, C => n124, Y => n126);
   U158 : NAND2X1 port map( A => n32, B => n126, Y => n127);
   U159 : OAI21X1 port map( A => n128, B => n127, C => n221, Y => n130);
   U162 : NAND3X1 port map( A => n131, B => n130, C => n16, Y => 
                           nextstate_1_port);
   U163 : INVX2 port map( A => n132, Y => n133);
   U166 : MUX2X1 port map( B => n134, A => n133, S => count_0_port, Y => n217);
   U169 : NOR2X1 port map( A => n223, B => n45, Y => n138);
   U170 : NAND2X1 port map( A => n4, B => n135, Y => n136);
   U171 : OAI21X1 port map( A => n153, B => n140, C => n136, Y => n137);
   U172 : OAI21X1 port map( A => n138, B => n137, C => n221, Y => n139);
   U173 : NAND2X1 port map( A => n1, B => n139, Y => n165);
   U174 : NAND2X1 port map( A => n29, B => D_EDGE, Y => n143);
   U175 : INVX2 port map( A => n140, Y => n141);
   U176 : NAND3X1 port map( A => n8, B => n141, C => n221, Y => n142);
   U177 : NAND2X1 port map( A => n143, B => n142, Y => n145);
   U178 : NOR2X1 port map( A => n153, B => n223, Y => n144);
   U179 : MUX2X1 port map( B => n145, A => n144, S => n49, Y => n148);
   U180 : OR2X2 port map( A => n219, B => n20, Y => n147);
   U181 : AOI21X1 port map( A => D_EDGE, B => n44, C => n168, Y => n146);
   U182 : NAND3X1 port map( A => n148, B => n147, C => n146, Y => n157);
   U183 : NAND2X1 port map( A => n49, B => n153, Y => n154);
   U184 : MUX2X1 port map( B => n157, A => n154, S => n47, Y => n160);
   U185 : INVX2 port map( A => n160, Y => n164);
   U186 : NAND2X1 port map( A => n165, B => n164, Y => nextstate_0_port);
   U187 : NOR2X1 port map( A => n219, B => n166, Y => n174);
   U188 : AOI22X1 port map( A => n3, B => BS_ERROR, C => D_EDGE, D => n20, Y =>
                           n171);
   U189 : NAND2X1 port map( A => n168, B => EOP, Y => n169);
   U190 : OAI21X1 port map( A => n171, B => n170_port, C => n169, Y => n173);
   U191 : OAI21X1 port map( A => n174, B => n173, C => n172, Y => n183);
   U192 : OAI21X1 port map( A => n18, B => n15, C => n175, Y => n176);
   U193 : AOI22X1 port map( A => n6, B => N170, C => BS_ERROR, D => n176, Y => 
                           n182);
   U194 : OAI21X1 port map( A => EOP, B => n28, C => n177, Y => n180);
   U195 : NOR2X1 port map( A => n180, B => n10, Y => n181);
   U196 : NAND3X1 port map( A => n183, B => n182, C => n181, Y => 
                           nextstate_3_port);
   U197 : XNOR2X1 port map( A => RX_CHECK_CRC(10), B => RX_CRC(10), Y => n190);
   U198 : XNOR2X1 port map( A => RX_CHECK_CRC(9), B => RX_CRC(9), Y => n189);
   U199 : XOR2X1 port map( A => RX_CHECK_CRC(7), B => RX_CRC(7), Y => n187);
   U200 : XOR2X1 port map( A => RX_CHECK_CRC(8), B => RX_CRC(8), Y => n186);
   U201 : NOR2X1 port map( A => n187, B => n186, Y => n188);
   U202 : NAND3X1 port map( A => n190, B => n189, C => n188, Y => n197);
   U203 : XNOR2X1 port map( A => RX_CHECK_CRC(14), B => RX_CRC(14), Y => n195);
   U204 : XNOR2X1 port map( A => RX_CHECK_CRC(13), B => RX_CRC(13), Y => n194);
   U205 : XOR2X1 port map( A => RX_CHECK_CRC(11), B => RX_CRC(11), Y => n192);
   U206 : XOR2X1 port map( A => RX_CHECK_CRC(12), B => RX_CRC(12), Y => n191);
   U207 : NOR2X1 port map( A => n192, B => n191, Y => n193);
   U208 : NAND3X1 port map( A => n195, B => n194, C => n193, Y => n196);
   U209 : NOR2X1 port map( A => n197, B => n196, Y => n213);
   U210 : NOR2X1 port map( A => n214, B => RX_CHECK_CRC(0), Y => n198);
   U211 : OAI22X1 port map( A => RX_CRC(1), B => n198, C => n198, D => n216, Y 
                           => n204);
   U212 : AND2X1 port map( A => RX_CHECK_CRC(0), B => n214, Y => n199);
   U213 : OAI22X1 port map( A => n199, B => n215, C => RX_CHECK_CRC(1), D => 
                           n199, Y => n203);
   U214 : XOR2X1 port map( A => RX_CHECK_CRC(15), B => RX_CRC(15), Y => n201);
   U215 : XOR2X1 port map( A => RX_CHECK_CRC(2), B => RX_CRC(2), Y => n200);
   U216 : NOR2X1 port map( A => n201, B => n200, Y => n202);
   U217 : NAND3X1 port map( A => n204, B => n203, C => n202, Y => n211);
   U218 : XNOR2X1 port map( A => RX_CHECK_CRC(6), B => RX_CRC(6), Y => n209);
   U219 : XNOR2X1 port map( A => RX_CHECK_CRC(5), B => RX_CRC(5), Y => n208);
   U220 : XOR2X1 port map( A => RX_CHECK_CRC(3), B => RX_CRC(3), Y => n206);
   U221 : XOR2X1 port map( A => RX_CHECK_CRC(4), B => RX_CRC(4), Y => n205);
   U222 : NOR2X1 port map( A => n206, B => n205, Y => n207);
   U223 : NAND3X1 port map( A => n209, B => n208, C => n207, Y => n210);
   U224 : NOR2X1 port map( A => n211, B => n210, Y => n212);
   U225 : AND2X1 port map( A => n213, B => n212, Y => N170);
   U226 : INVX2 port map( A => RX_CRC(0), Y => n214);
   U227 : INVX2 port map( A => RX_CRC(1), Y => n215);
   U228 : INVX2 port map( A => RX_CHECK_CRC(1), Y => n216);
   U229 : INVX2 port map( A => n87, Y => n218);
   U230 : INVX2 port map( A => n83, Y => n219);
   U231 : INVX2 port map( A => curR_ERROR, Y => n220);
   U232 : INVX2 port map( A => BS_ERROR, Y => n221);
   U233 : INVX2 port map( A => N170, Y => n222);
   U234 : INVX2 port map( A => EOP, Y => n223);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_eopdetect_1 is

   port( DP1_RX, DM1_RX : in std_logic;  EOP : out std_logic);

end rx_eopdetect_1;

architecture SYN_Behavioral of rx_eopdetect_1 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;

begin
   
   U1 : NOR2X1 port map( A => DP1_RX, B => DM1_RX, Y => EOP);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_edgedetect_1 is

   port( CLK, RST, DP1_RX : in std_logic;  D_EDGE : out std_logic);

end rx_edgedetect_1;

architecture SYN_Behavioral of rx_edgedetect_1 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal DP_hold1, DP_hold2, n1, n3, n2, n4 : std_logic;

begin
   
   DP_hold1_reg : DFFSR port map( D => DP1_RX, CLK => CLK, R => n3, S => n2, Q 
                           => DP_hold1);
   DP_hold2_reg : DFFSR port map( D => DP_hold1, CLK => CLK, R => n1, S => n2, 
                           Q => DP_hold2);
   n1 <= '1';
   n3 <= '1';
   U4 : INVX2 port map( A => RST, Y => n2);
   U6 : XNOR2X1 port map( A => DP_hold2, B => DP_hold1, Y => n4);
   U7 : NOR2X1 port map( A => RST, B => n4, Y => D_EDGE);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_decode_1 is

   port( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP : in std_logic;  D_ORIG, BITSTUFF,
         BS_ERROR : out std_logic);

end rx_decode_1;

architecture SYN_moore of rx_decode_1 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal DP_hold1, DP_hold2, state_3_port, state_2_port, state_1_port, 
      state_0_port, N29, N30, N31, N32, n1, n4, n7, n17, n19, n43, n44, n2, n3,
      n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29_port, n30_port, n31_port, n32_port, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, BS_ERROR_port : std_logic;

begin
   BS_ERROR <= BS_ERROR_port;
   
   DP_hold2_reg : DFFSR port map( D => n44, CLK => CLK, R => n7, S => n9, Q => 
                           DP_hold2);
   state_reg_3_inst : DFFSR port map( D => N32, CLK => CLK, R => n9, S => n4, Q
                           => state_3_port);
   DP_hold1_reg : DFFSR port map( D => n43, CLK => CLK, R => n1, S => n9, Q => 
                           DP_hold1);
   n1 <= '1';
   n4 <= '1';
   n7 <= '1';
   U20 : NAND2X1 port map( A => n17, B => n41, Y => n43);
   U21 : AOI22X1 port map( A => DP_hold1, B => n42, C => DP1_RX, D => n19, Y =>
                           n17);
   U25 : XNOR2X1 port map( A => DP_hold1, B => DP_hold2, Y => D_ORIG);
   state_reg_0_inst : DFFSR port map( D => N29, CLK => CLK, R => n9, S => n6, Q
                           => state_0_port);
   state_reg_2_inst : DFFSR port map( D => N31, CLK => CLK, R => n9, S => n5, Q
                           => state_2_port);
   state_reg_1_inst : DFFSR port map( D => N30, CLK => CLK, R => n9, S => n3, Q
                           => state_1_port);
   U4 : AND2X2 port map( A => state_1_port, B => state_2_port, Y => n2);
   n3 <= '1';
   n5 <= '1';
   n6 <= '1';
   U10 : INVX1 port map( A => SHIFT_ENABLE, Y => n31_port);
   U11 : AND2X1 port map( A => SHIFT_ENABLE, B => state_0_port, Y => n22);
   U12 : INVX2 port map( A => RST, Y => n9);
   U13 : MUX2X1 port map( B => DP_hold1, A => DP_hold2, S => n8, Y => n40);
   U14 : NAND2X1 port map( A => SHIFT_ENABLE, B => n19, Y => n8);
   U15 : INVX2 port map( A => state_0_port, Y => n15);
   U16 : NOR2X1 port map( A => state_1_port, B => state_2_port, Y => n10);
   U17 : NAND3X1 port map( A => state_3_port, B => n15, C => n10, Y => n11);
   U18 : INVX2 port map( A => n11, Y => BS_ERROR_port);
   U19 : NAND2X1 port map( A => n2, B => n15, Y => n19);
   U22 : NOR2X1 port map( A => state_3_port, B => n19, Y => BITSTUFF);
   U23 : INVX2 port map( A => n19, Y => n42);
   U24 : OR2X2 port map( A => EOP, B => state_3_port, Y => n37);
   U26 : INVX2 port map( A => n37, Y => n41);
   U27 : INVX2 port map( A => DP1_RX, Y => n12);
   U28 : XOR2X1 port map( A => n12, B => DP_hold2, Y => n33);
   U29 : INVX2 port map( A => n33, Y => n24);
   U30 : NOR2X1 port map( A => state_0_port, B => n24, Y => n13);
   U31 : MUX2X1 port map( B => n13, A => n24, S => n2, Y => n14);
   U32 : MUX2X1 port map( B => n15, A => n14, S => SHIFT_ENABLE, Y => n16);
   U33 : AND2X2 port map( A => n41, B => n16, Y => N29);
   U34 : INVX2 port map( A => state_2_port, Y => n18);
   U35 : NAND3X1 port map( A => state_1_port, B => n33, C => n18, Y => n35);
   U36 : INVX2 port map( A => n35, Y => n23);
   U37 : INVX2 port map( A => state_1_port, Y => n32_port);
   U38 : NAND2X1 port map( A => n33, B => n32_port, Y => n20);
   U39 : AOI21X1 port map( A => SHIFT_ENABLE, B => n20, C => n18, Y => n21);
   U40 : AOI21X1 port map( A => n23, B => n22, C => n21, Y => n25);
   U41 : NAND2X1 port map( A => n24, B => n42, Y => n29_port);
   U42 : AOI21X1 port map( A => n25, B => n29_port, C => n37, Y => N31);
   U43 : NAND3X1 port map( A => n33, B => n42, C => SHIFT_ENABLE, Y => n28);
   U44 : INVX2 port map( A => EOP, Y => n26);
   U45 : NAND2X1 port map( A => BS_ERROR_port, B => n26, Y => n27);
   U46 : OAI21X1 port map( A => n37, B => n28, C => n27, Y => N32);
   U47 : INVX2 port map( A => n29_port, Y => n30_port);
   U48 : AOI21X1 port map( A => state_1_port, B => n31_port, C => n30_port, Y 
                           => n39);
   U49 : NAND3X1 port map( A => SHIFT_ENABLE, B => n33, C => n32_port, Y => n34
                           );
   U50 : MUX2X1 port map( B => n35, A => n34, S => state_0_port, Y => n36);
   U51 : INVX2 port map( A => n36, Y => n38);
   U52 : AOI21X1 port map( A => n39, B => n38, C => n37, Y => N30);
   U53 : NAND2X1 port map( A => n41, B => n40, Y => n44);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_accumulator_1 is

   port( CLK, RST : in std_logic;  RCV_DATA : in std_logic_vector (7 downto 0);
         W_ENABLE : in std_logic;  rx_CHECK_CRC : out std_logic_vector (15 
         downto 0));

end rx_accumulator_1;

architecture SYN_Behavioral of rx_accumulator_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, rx_CHECK_CRC_13_port, 
      rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, rx_CHECK_CRC_10_port, 
      rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, rx_CHECK_CRC_7_port, 
      rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, rx_CHECK_CRC_4_port, 
      rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, rx_CHECK_CRC_1_port, 
      rx_CHECK_CRC_0_port, n3, n4, n6, n7, n9, n10, n12, n13, n15, n16, n18, 
      n19, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55, n57, n58, n1, n2, n5, n8, n11, n14, n17, 
      n20, n23, n56, n59, n60 : std_logic;

begin
   rx_CHECK_CRC <= ( rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, 
      rx_CHECK_CRC_13_port, rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, 
      rx_CHECK_CRC_10_port, rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, 
      rx_CHECK_CRC_7_port, rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, 
      rx_CHECK_CRC_4_port, rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, 
      rx_CHECK_CRC_1_port, rx_CHECK_CRC_0_port );
   
   present_CHECK_CRC_reg_7_inst : DFFSR port map( D => n58, CLK => CLK, R => n5
                           , S => n57, Q => rx_CHECK_CRC_7_port);
   present_CHECK_CRC_reg_15_inst : DFFSR port map( D => n55, CLK => CLK, R => 
                           n5, S => n54, Q => rx_CHECK_CRC_15_port);
   present_CHECK_CRC_reg_6_inst : DFFSR port map( D => n53, CLK => CLK, R => n5
                           , S => n52, Q => rx_CHECK_CRC_6_port);
   present_CHECK_CRC_reg_14_inst : DFFSR port map( D => n51, CLK => CLK, R => 
                           n5, S => n50, Q => rx_CHECK_CRC_14_port);
   present_CHECK_CRC_reg_5_inst : DFFSR port map( D => n49, CLK => CLK, R => n5
                           , S => n48, Q => rx_CHECK_CRC_5_port);
   present_CHECK_CRC_reg_13_inst : DFFSR port map( D => n47, CLK => CLK, R => 
                           n5, S => n46, Q => rx_CHECK_CRC_13_port);
   present_CHECK_CRC_reg_4_inst : DFFSR port map( D => n45, CLK => CLK, R => n5
                           , S => n44, Q => rx_CHECK_CRC_4_port);
   present_CHECK_CRC_reg_12_inst : DFFSR port map( D => n43, CLK => CLK, R => 
                           n5, S => n42, Q => rx_CHECK_CRC_12_port);
   present_CHECK_CRC_reg_3_inst : DFFSR port map( D => n41, CLK => CLK, R => n5
                           , S => n40, Q => rx_CHECK_CRC_3_port);
   present_CHECK_CRC_reg_11_inst : DFFSR port map( D => n39, CLK => CLK, R => 
                           n5, S => n38, Q => rx_CHECK_CRC_11_port);
   present_CHECK_CRC_reg_2_inst : DFFSR port map( D => n37, CLK => CLK, R => n5
                           , S => n36, Q => rx_CHECK_CRC_2_port);
   present_CHECK_CRC_reg_10_inst : DFFSR port map( D => n35, CLK => CLK, R => 
                           n5, S => n34, Q => rx_CHECK_CRC_10_port);
   present_CHECK_CRC_reg_1_inst : DFFSR port map( D => n33, CLK => CLK, R => n5
                           , S => n32, Q => rx_CHECK_CRC_1_port);
   present_CHECK_CRC_reg_9_inst : DFFSR port map( D => n31, CLK => CLK, R => n5
                           , S => n30, Q => rx_CHECK_CRC_9_port);
   present_CHECK_CRC_reg_0_inst : DFFSR port map( D => n29, CLK => CLK, R => n5
                           , S => n28, Q => rx_CHECK_CRC_0_port);
   present_CHECK_CRC_reg_8_inst : DFFSR port map( D => n27, CLK => CLK, R => n5
                           , S => n26, Q => rx_CHECK_CRC_8_port);
   U2 : OAI21X1 port map( A => n8, B => n60, C => n3, Y => n27);
   U3 : NAND2X1 port map( A => rx_CHECK_CRC_8_port, B => n8, Y => n3);
   U4 : OAI21X1 port map( A => n2, B => n60, C => n4, Y => n29);
   U5 : NAND2X1 port map( A => RCV_DATA(0), B => n2, Y => n4);
   U7 : OAI21X1 port map( A => n8, B => n59, C => n6, Y => n31);
   U8 : NAND2X1 port map( A => rx_CHECK_CRC_9_port, B => n8, Y => n6);
   U9 : OAI21X1 port map( A => n2, B => n59, C => n7, Y => n33);
   U10 : NAND2X1 port map( A => RCV_DATA(1), B => n2, Y => n7);
   U12 : OAI21X1 port map( A => n8, B => n56, C => n9, Y => n35);
   U13 : NAND2X1 port map( A => rx_CHECK_CRC_10_port, B => n8, Y => n9);
   U14 : OAI21X1 port map( A => n2, B => n56, C => n10, Y => n37);
   U15 : NAND2X1 port map( A => RCV_DATA(2), B => n2, Y => n10);
   U17 : OAI21X1 port map( A => n8, B => n23, C => n12, Y => n39);
   U18 : NAND2X1 port map( A => rx_CHECK_CRC_11_port, B => n8, Y => n12);
   U19 : OAI21X1 port map( A => n2, B => n23, C => n13, Y => n41);
   U20 : NAND2X1 port map( A => RCV_DATA(3), B => n2, Y => n13);
   U22 : OAI21X1 port map( A => n8, B => n20, C => n15, Y => n43);
   U23 : NAND2X1 port map( A => rx_CHECK_CRC_12_port, B => n8, Y => n15);
   U24 : OAI21X1 port map( A => n2, B => n20, C => n16, Y => n45);
   U25 : NAND2X1 port map( A => RCV_DATA(4), B => n2, Y => n16);
   U27 : OAI21X1 port map( A => n8, B => n17, C => n18, Y => n47);
   U28 : NAND2X1 port map( A => rx_CHECK_CRC_13_port, B => n8, Y => n18);
   U29 : OAI21X1 port map( A => n2, B => n17, C => n19, Y => n49);
   U30 : NAND2X1 port map( A => RCV_DATA(5), B => n2, Y => n19);
   U32 : OAI21X1 port map( A => n8, B => n14, C => n21, Y => n51);
   U33 : NAND2X1 port map( A => rx_CHECK_CRC_14_port, B => n8, Y => n21);
   U34 : OAI21X1 port map( A => n2, B => n14, C => n22, Y => n53);
   U35 : NAND2X1 port map( A => RCV_DATA(6), B => n2, Y => n22);
   U37 : OAI21X1 port map( A => n8, B => n11, C => n24, Y => n55);
   U38 : NAND2X1 port map( A => rx_CHECK_CRC_15_port, B => n8, Y => n24);
   U41 : OAI21X1 port map( A => n2, B => n11, C => n25, Y => n58);
   U42 : NAND2X1 port map( A => RCV_DATA(7), B => n2, Y => n25);
   n26 <= '1';
   n28 <= '1';
   n30 <= '1';
   n32 <= '1';
   n34 <= '1';
   n36 <= '1';
   n38 <= '1';
   n40 <= '1';
   n42 <= '1';
   n44 <= '1';
   n46 <= '1';
   n48 <= '1';
   n50 <= '1';
   n52 <= '1';
   n54 <= '1';
   n57 <= '1';
   U6 : INVX4 port map( A => n2, Y => n8);
   U11 : INVX4 port map( A => n1, Y => n2);
   U16 : INVX2 port map( A => W_ENABLE, Y => n1);
   U21 : INVX2 port map( A => RST, Y => n5);
   U26 : INVX2 port map( A => rx_CHECK_CRC_7_port, Y => n11);
   U31 : INVX2 port map( A => rx_CHECK_CRC_6_port, Y => n14);
   U36 : INVX2 port map( A => rx_CHECK_CRC_5_port, Y => n17);
   U39 : INVX2 port map( A => rx_CHECK_CRC_4_port, Y => n20);
   U40 : INVX2 port map( A => rx_CHECK_CRC_3_port, Y => n23);
   U43 : INVX2 port map( A => rx_CHECK_CRC_2_port, Y => n56);
   U60 : INVX2 port map( A => rx_CHECK_CRC_1_port, Y => n59);
   U61 : INVX2 port map( A => rx_CHECK_CRC_0_port, Y => n60);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_CRC_CALC_1 is

   port( CLK, RST, W_ENABLE : in std_logic;  OPCODE : in std_logic_vector (1 
         downto 0);  RCV_DATA : in std_logic_vector (7 downto 0);  RX_CRC : out
         std_logic_vector (15 downto 0));

end rx_CRC_CALC_1;

architecture SYN_moore of rx_CRC_CALC_1 is

   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port, current_crc_15_port, 
      current_crc_14_port, current_crc_13_port, current_crc_12_port, 
      current_crc_11_port, current_crc_10_port, current_crc_9_port, 
      current_crc_8_port, current_crc_7_port, current_crc_6_port, 
      current_crc_5_port, current_crc_4_port, current_crc_3_port, 
      current_crc_2_port, current_crc_1_port, current_crc_0_port, 
      cache_1_15_port, cache_1_14_port, cache_1_13_port, cache_1_12_port, 
      cache_1_11_port, cache_1_10_port, cache_1_9_port, cache_1_8_port, 
      cache_1_7_port, cache_1_6_port, cache_1_5_port, cache_1_4_port, 
      cache_1_3_port, cache_1_2_port, cache_1_1_port, cache_1_0_port, n83, n84,
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n101, n103, n105, n107, n109, n111, n113, n115, n117, n119, n121, n123,
      n125, n127, n129, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n100, n102, n104, n106, n108, n110, n112, n114, n116, n118, n120, 
      n122, n124, n126, n128, n130, n131, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n_1029, n_1030, n_1031 : 
      std_logic;

begin
   RX_CRC <= ( RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port );
   
   cache_1_reg_0_inst : DFFPOSX1 port map( D => n129, CLK => CLK, Q => 
                           cache_1_0_port);
   cache_1_reg_8_inst : DFFPOSX1 port map( D => n127, CLK => CLK, Q => 
                           cache_1_8_port);
   cache_1_reg_15_inst : DFFPOSX1 port map( D => n125, CLK => CLK, Q => 
                           cache_1_15_port);
   cache_1_reg_1_inst : DFFPOSX1 port map( D => n123, CLK => CLK, Q => 
                           cache_1_1_port);
   cache_1_reg_9_inst : DFFPOSX1 port map( D => n121, CLK => CLK, Q => 
                           cache_1_9_port);
   cache_1_reg_2_inst : DFFPOSX1 port map( D => n119, CLK => CLK, Q => 
                           cache_1_2_port);
   cache_1_reg_10_inst : DFFPOSX1 port map( D => n117, CLK => CLK, Q => 
                           cache_1_10_port);
   cache_1_reg_3_inst : DFFPOSX1 port map( D => n115, CLK => CLK, Q => 
                           cache_1_3_port);
   cache_1_reg_11_inst : DFFPOSX1 port map( D => n113, CLK => CLK, Q => 
                           cache_1_11_port);
   cache_1_reg_4_inst : DFFPOSX1 port map( D => n111, CLK => CLK, Q => 
                           cache_1_4_port);
   cache_1_reg_12_inst : DFFPOSX1 port map( D => n109, CLK => CLK, Q => 
                           cache_1_12_port);
   cache_1_reg_5_inst : DFFPOSX1 port map( D => n107, CLK => CLK, Q => 
                           cache_1_5_port);
   cache_1_reg_13_inst : DFFPOSX1 port map( D => n105, CLK => CLK, Q => 
                           cache_1_13_port);
   cache_1_reg_6_inst : DFFPOSX1 port map( D => n103, CLK => CLK, Q => 
                           cache_1_6_port);
   cache_1_reg_14_inst : DFFPOSX1 port map( D => n101, CLK => CLK, Q => 
                           cache_1_14_port);
   cache_1_reg_7_inst : DFFPOSX1 port map( D => n99, CLK => CLK, Q => 
                           cache_1_7_port);
   cache_2_reg_15_inst : DFFPOSX1 port map( D => n98, CLK => CLK, Q => 
                           RX_CRC_15_port);
   cache_2_reg_14_inst : DFFPOSX1 port map( D => n97, CLK => CLK, Q => 
                           RX_CRC_14_port);
   cache_2_reg_13_inst : DFFPOSX1 port map( D => n96, CLK => CLK, Q => 
                           RX_CRC_13_port);
   cache_2_reg_12_inst : DFFPOSX1 port map( D => n95, CLK => CLK, Q => 
                           RX_CRC_12_port);
   cache_2_reg_11_inst : DFFPOSX1 port map( D => n94, CLK => CLK, Q => 
                           RX_CRC_11_port);
   cache_2_reg_10_inst : DFFPOSX1 port map( D => n93, CLK => CLK, Q => 
                           RX_CRC_10_port);
   cache_2_reg_9_inst : DFFPOSX1 port map( D => n92, CLK => CLK, Q => 
                           RX_CRC_9_port);
   cache_2_reg_8_inst : DFFPOSX1 port map( D => n91, CLK => CLK, Q => 
                           RX_CRC_8_port);
   cache_2_reg_7_inst : DFFPOSX1 port map( D => n90, CLK => CLK, Q => 
                           RX_CRC_7_port);
   cache_2_reg_6_inst : DFFPOSX1 port map( D => n89, CLK => CLK, Q => 
                           RX_CRC_6_port);
   cache_2_reg_5_inst : DFFPOSX1 port map( D => n88, CLK => CLK, Q => 
                           RX_CRC_5_port);
   cache_2_reg_4_inst : DFFPOSX1 port map( D => n87, CLK => CLK, Q => 
                           RX_CRC_4_port);
   cache_2_reg_3_inst : DFFPOSX1 port map( D => n86, CLK => CLK, Q => 
                           RX_CRC_3_port);
   cache_2_reg_2_inst : DFFPOSX1 port map( D => n85, CLK => CLK, Q => 
                           RX_CRC_2_port);
   cache_2_reg_1_inst : DFFPOSX1 port map( D => n84, CLK => CLK, Q => 
                           RX_CRC_1_port);
   cache_2_reg_0_inst : DFFPOSX1 port map( D => n83, CLK => CLK, Q => 
                           RX_CRC_0_port);
   current_crc_reg_15_inst : DFFSR port map( D => n132, CLK => CLK, R => n35, S
                           => n17, Q => current_crc_15_port);
   current_crc_reg_14_inst : DFFSR port map( D => n133, CLK => CLK, R => n35, S
                           => n16, Q => current_crc_14_port);
   current_crc_reg_13_inst : DFFSR port map( D => n134, CLK => CLK, R => n35, S
                           => n15, Q => current_crc_13_port);
   current_crc_reg_12_inst : DFFSR port map( D => n135, CLK => CLK, R => n35, S
                           => n14, Q => current_crc_12_port);
   current_crc_reg_11_inst : DFFSR port map( D => n136, CLK => CLK, R => n35, S
                           => n13, Q => current_crc_11_port);
   current_crc_reg_10_inst : DFFSR port map( D => n137, CLK => CLK, R => n35, S
                           => n12, Q => current_crc_10_port);
   current_crc_reg_9_inst : DFFSR port map( D => n138, CLK => CLK, R => n35, S 
                           => n11, Q => current_crc_9_port);
   current_crc_reg_8_inst : DFFSR port map( D => n139, CLK => CLK, R => n35, S 
                           => n10, Q => current_crc_8_port);
   current_crc_reg_7_inst : DFFSR port map( D => n140, CLK => CLK, R => n35, S 
                           => n9, Q => current_crc_7_port);
   current_crc_reg_6_inst : DFFSR port map( D => n141, CLK => CLK, R => n35, S 
                           => n8, Q => current_crc_6_port);
   current_crc_reg_5_inst : DFFSR port map( D => n142, CLK => CLK, R => n35, S 
                           => n7, Q => current_crc_5_port);
   current_crc_reg_4_inst : DFFSR port map( D => n143, CLK => CLK, R => n35, S 
                           => n6, Q => current_crc_4_port);
   current_crc_reg_3_inst : DFFSR port map( D => n144, CLK => CLK, R => n35, S 
                           => n5, Q => current_crc_3_port);
   current_crc_reg_2_inst : DFFSR port map( D => n145, CLK => CLK, R => n35, S 
                           => n4, Q => current_crc_2_port);
   current_crc_reg_1_inst : DFFSR port map( D => n146, CLK => CLK, R => n35, S 
                           => n3, Q => current_crc_1_port);
   current_crc_reg_0_inst : DFFSR port map( D => n147, CLK => CLK, R => n35, S 
                           => n2, Q => current_crc_0_port);
   U3 : INVX2 port map( A => n28, Y => n20);
   U4 : XOR2X1 port map( A => n27, B => n25, Y => n1);
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   U21 : INVX2 port map( A => n53, Y => n19);
   U22 : INVX2 port map( A => OPCODE(1), Y => n34);
   U23 : AND2X2 port map( A => n19, B => n35, Y => n18);
   U24 : INVX4 port map( A => n21, Y => n33);
   U25 : AND2X2 port map( A => n19, B => n35, Y => n21);
   U26 : INVX2 port map( A => n22, Y => n30);
   U27 : INVX2 port map( A => n22, Y => n29);
   U28 : AND2X2 port map( A => n54, B => n28, Y => n22);
   U29 : INVX2 port map( A => RST, Y => n35);
   U30 : XNOR2X1 port map( A => n63, B => n27, Y => n64);
   U31 : XNOR2X1 port map( A => RCV_DATA(6), B => current_crc_14_port, Y => 
                           n161);
   U32 : XNOR2X1 port map( A => RCV_DATA(7), B => current_crc_15_port, Y => 
                           n148);
   U33 : XOR2X1 port map( A => RCV_DATA(0), B => current_crc_8_port, Y => n23);
   U34 : XNOR2X1 port map( A => RCV_DATA(5), B => current_crc_13_port, Y => n63
                           );
   U35 : XOR2X1 port map( A => RCV_DATA(1), B => current_crc_9_port, Y => n24);
   U36 : XOR2X1 port map( A => RCV_DATA(3), B => current_crc_11_port, Y => n25)
                           ;
   U37 : XOR2X1 port map( A => RCV_DATA(2), B => current_crc_10_port, Y => n26)
                           ;
   U38 : XOR2X1 port map( A => RCV_DATA(4), B => current_crc_12_port, Y => n27)
                           ;
   U39 : NAND3X1 port map( A => OPCODE(0), B => W_ENABLE, C => n34, Y => n28);
   U40 : INVX8 port map( A => n33, Y => n31);
   U41 : INVX8 port map( A => n33, Y => n32);
   U42 : INVX2 port map( A => RX_CRC_0_port, Y => n36);
   U43 : INVX2 port map( A => cache_1_0_port, Y => n165);
   U44 : NAND3X1 port map( A => OPCODE(0), B => W_ENABLE, C => n34, Y => n53);
   U45 : MUX2X1 port map( B => n36, A => n165, S => n31, Y => n83);
   U46 : INVX2 port map( A => RX_CRC_1_port, Y => n37);
   U47 : INVX2 port map( A => cache_1_1_port, Y => n130);
   U48 : MUX2X1 port map( B => n37, A => n130, S => n32, Y => n84);
   U49 : INVX2 port map( A => RX_CRC_2_port, Y => n38);
   U50 : INVX2 port map( A => cache_1_2_port, Y => n114);
   U51 : MUX2X1 port map( B => n38, A => n114, S => n31, Y => n85);
   U52 : INVX2 port map( A => RX_CRC_3_port, Y => n39);
   U53 : INVX2 port map( A => cache_1_3_port, Y => n100);
   U54 : MUX2X1 port map( B => n39, A => n100, S => n32, Y => n86);
   U55 : INVX2 port map( A => RX_CRC_4_port, Y => n40);
   U56 : INVX2 port map( A => cache_1_4_port, Y => n76);
   U57 : MUX2X1 port map( B => n40, A => n76, S => n31, Y => n87);
   U58 : INVX2 port map( A => RX_CRC_5_port, Y => n41);
   U59 : INVX2 port map( A => cache_1_5_port, Y => n70);
   U60 : MUX2X1 port map( B => n41, A => n70, S => n31, Y => n88);
   U61 : INVX2 port map( A => RX_CRC_6_port, Y => n42);
   U62 : INVX2 port map( A => cache_1_6_port, Y => n62);
   U63 : MUX2X1 port map( B => n42, A => n62, S => n31, Y => n89);
   U64 : INVX2 port map( A => RX_CRC_7_port, Y => n43);
   U65 : INVX2 port map( A => cache_1_7_port, Y => n52);
   U66 : MUX2X1 port map( B => n43, A => n52, S => n32, Y => n90);
   U67 : INVX2 port map( A => RX_CRC_8_port, Y => n44);
   U68 : INVX2 port map( A => cache_1_8_port, Y => n160);
   U69 : MUX2X1 port map( B => n44, A => n160, S => n31, Y => n91);
   U70 : INVX2 port map( A => RX_CRC_9_port, Y => n45);
   U71 : INVX2 port map( A => cache_1_9_port, Y => n122);
   U72 : MUX2X1 port map( B => n45, A => n122, S => n31, Y => n92);
   U73 : INVX2 port map( A => RX_CRC_10_port, Y => n46);
   U74 : INVX2 port map( A => cache_1_10_port, Y => n108);
   U75 : MUX2X1 port map( B => n46, A => n108, S => n31, Y => n93);
   U76 : INVX2 port map( A => RX_CRC_11_port, Y => n47);
   U77 : INVX2 port map( A => cache_1_11_port, Y => n80);
   U78 : MUX2X1 port map( B => n47, A => n80, S => n31, Y => n94);
   U79 : INVX2 port map( A => RX_CRC_12_port, Y => n48);
   U80 : INVX2 port map( A => cache_1_12_port, Y => n73);
   U81 : MUX2X1 port map( B => n48, A => n73, S => n31, Y => n95);
   U82 : INVX2 port map( A => RX_CRC_13_port, Y => n49);
   U83 : INVX2 port map( A => cache_1_13_port, Y => n67);
   U84 : MUX2X1 port map( B => n49, A => n67, S => n31, Y => n96);
   U85 : INVX2 port map( A => RX_CRC_14_port, Y => n50);
   U86 : INVX2 port map( A => cache_1_14_port, Y => n59);
   U87 : MUX2X1 port map( B => n50, A => n59, S => n31, Y => n97);
   U88 : INVX2 port map( A => RX_CRC_15_port, Y => n51);
   U89 : INVX2 port map( A => cache_1_15_port, Y => n153);
   U90 : MUX2X1 port map( B => n51, A => n153, S => n31, Y => n98);
   U91 : INVX2 port map( A => current_crc_7_port, Y => n58);
   U92 : MUX2X1 port map( B => n52, A => n58, S => n18, Y => n99);
   U93 : NAND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n54);
   U94 : INVX2 port map( A => n161, Y => n55);
   U95 : XOR2X1 port map( A => n63, B => n55, Y => n168);
   U96 : INVX2 port map( A => n168, Y => n56);
   U97 : NAND2X1 port map( A => n20, B => n56, Y => n57);
   U98 : OAI21X1 port map( A => n29, B => n58, C => n57, Y => n140);
   U99 : INVX2 port map( A => current_crc_14_port, Y => n61);
   U100 : MUX2X1 port map( B => n59, A => n61, S => n18, Y => n101);
   U101 : NAND2X1 port map( A => current_crc_6_port, B => n20, Y => n60);
   U102 : OAI21X1 port map( A => n30, B => n61, C => n60, Y => n133);
   U103 : INVX2 port map( A => current_crc_6_port, Y => n66);
   U104 : MUX2X1 port map( B => n62, A => n66, S => n32, Y => n103);
   U105 : NAND2X1 port map( A => n20, B => n64, Y => n65);
   U106 : OAI21X1 port map( A => n29, B => n66, C => n65, Y => n141);
   U107 : INVX2 port map( A => current_crc_13_port, Y => n69);
   U108 : MUX2X1 port map( B => n67, A => n69, S => n18, Y => n105);
   U109 : NAND2X1 port map( A => current_crc_5_port, B => n20, Y => n68);
   U110 : OAI21X1 port map( A => n30, B => n69, C => n68, Y => n134);
   U111 : INVX2 port map( A => current_crc_5_port, Y => n72);
   U112 : MUX2X1 port map( B => n70, A => n72, S => n32, Y => n107);
   U113 : NAND2X1 port map( A => n20, B => n1, Y => n71);
   U114 : OAI21X1 port map( A => n29, B => n72, C => n71, Y => n142);
   U115 : INVX2 port map( A => current_crc_12_port, Y => n75);
   U116 : MUX2X1 port map( B => n73, A => n75, S => n32, Y => n109);
   U117 : NAND2X1 port map( A => current_crc_4_port, B => n20, Y => n74);
   U118 : OAI21X1 port map( A => n30, B => n75, C => n74, Y => n135);
   U119 : INVX2 port map( A => current_crc_4_port, Y => n79);
   U120 : MUX2X1 port map( B => n76, A => n79, S => n32, Y => n111);
   U121 : XOR2X1 port map( A => n25, B => n26, Y => n77);
   U122 : NAND2X1 port map( A => n20, B => n77, Y => n78);
   U123 : OAI21X1 port map( A => n29, B => n79, C => n78, Y => n143);
   U124 : INVX2 port map( A => current_crc_11_port, Y => n82);
   U125 : MUX2X1 port map( B => n80, A => n82, S => n32, Y => n113);
   U126 : NAND2X1 port map( A => current_crc_3_port, B => n20, Y => n81);
   U127 : OAI21X1 port map( A => n30, B => n82, C => n81, Y => n136);
   U128 : INVX2 port map( A => current_crc_3_port, Y => n106);
   U129 : MUX2X1 port map( B => n100, A => n106, S => n32, Y => n115);
   U130 : XNOR2X1 port map( A => n26, B => n24, Y => n131);
   U131 : INVX2 port map( A => n131, Y => n102);
   U132 : NAND2X1 port map( A => n20, B => n102, Y => n104);
   U133 : OAI21X1 port map( A => n29, B => n106, C => n104, Y => n144);
   U134 : INVX2 port map( A => current_crc_10_port, Y => n112);
   U135 : MUX2X1 port map( B => n108, A => n112, S => n18, Y => n117);
   U136 : NAND2X1 port map( A => current_crc_2_port, B => n20, Y => n110);
   U137 : OAI21X1 port map( A => n30, B => n112, C => n110, Y => n137);
   U138 : INVX2 port map( A => current_crc_2_port, Y => n120);
   U139 : MUX2X1 port map( B => n114, A => n120, S => n32, Y => n119);
   U140 : XOR2X1 port map( A => n23, B => n24, Y => n116);
   U141 : NAND2X1 port map( A => n20, B => n116, Y => n118);
   U142 : OAI21X1 port map( A => n29, B => n120, C => n118, Y => n145);
   U143 : INVX2 port map( A => current_crc_9_port, Y => n128);
   U144 : MUX2X1 port map( B => n122, A => n128, S => n32, Y => n121);
   U145 : INVX2 port map( A => n148, Y => n166);
   U146 : INVX2 port map( A => current_crc_1_port, Y => n152);
   U147 : XNOR2X1 port map( A => n166, B => n152, Y => n124);
   U148 : NAND2X1 port map( A => n20, B => n124, Y => n126);
   U149 : OAI21X1 port map( A => n30, B => n128, C => n126, Y => n138);
   U150 : MUX2X1 port map( B => n130, A => n152, S => n18, Y => n123);
   U151 : XOR2X1 port map( A => n131, B => n1, Y => n167);
   U152 : INVX2 port map( A => n167, Y => n156);
   U153 : XNOR2X1 port map( A => n168, B => n148, Y => n149);
   U154 : XNOR2X1 port map( A => n156, B => n149, Y => n150);
   U155 : NAND2X1 port map( A => n20, B => n150, Y => n151);
   U156 : OAI21X1 port map( A => n29, B => n152, C => n151, Y => n146);
   U157 : INVX2 port map( A => current_crc_15_port, Y => n159);
   U158 : MUX2X1 port map( B => n153, A => n159, S => n18, Y => n125);
   U159 : FAX1 port map( A => current_crc_7_port, B => n23, C => n166, YC => 
                           n_1029, YS => n154);
   U160 : XNOR2X1 port map( A => n154, B => n168, Y => n155);
   U161 : XOR2X1 port map( A => n156, B => n155, Y => n157);
   U162 : NAND2X1 port map( A => n20, B => n157, Y => n158);
   U163 : OAI21X1 port map( A => n30, B => n159, C => n158, Y => n132);
   U164 : INVX2 port map( A => current_crc_8_port, Y => n164);
   U165 : MUX2X1 port map( B => n160, A => n164, S => n32, Y => n127);
   U166 : INVX2 port map( A => current_crc_0_port, Y => n172);
   U167 : FAX1 port map( A => n166, B => n172, C => n161, YC => n_1030, YS => 
                           n162);
   U168 : NAND2X1 port map( A => n20, B => n162, Y => n163);
   U169 : OAI21X1 port map( A => n29, B => n164, C => n163, Y => n139);
   U170 : MUX2X1 port map( B => n165, A => n172, S => n18, Y => n129);
   U171 : XOR2X1 port map( A => n23, B => n166, Y => n169);
   U172 : FAX1 port map( A => n169, B => n168, C => n167, YC => n_1031, YS => 
                           n170);
   U173 : NAND2X1 port map( A => n20, B => n170, Y => n171);
   U174 : OAI21X1 port map( A => n30, B => n172, C => n171, Y => n147);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RFIFO_1 is

   port( CLK, RST, W_ENABLE, R_ENABLE : in std_logic;  RCV_DATA : in 
         std_logic_vector (7 downto 0);  RCV_OPCODE : in std_logic_vector (1 
         downto 0);  DATA : out std_logic_vector (7 downto 0);  OUT_OPCODE : 
         out std_logic_vector (1 downto 0);  BYTE_COUNT : out std_logic_vector 
         (4 downto 0);  EMPTY, FULL : out std_logic);

end RFIFO_1;

architecture SYN_BRFIFO of RFIFO_1 is

   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, 
      DATA_3_port, DATA_2_port, DATA_1_port, DATA_0_port, OUT_OPCODE_1_port, 
      OUT_OPCODE_0_port, EMPTY_port, FULL_port, readptr_4_port, readptr_3_port,
      readptr_2_port, readptr_1_port, readptr_0_port, writeptr_4_port, 
      writeptr_3_port, writeptr_2_port, writeptr_1_port, writeptr_0_port, state
      , opcode_0_1_port, opcode_0_0_port, opcode_1_1_port, opcode_1_0_port, 
      opcode_2_1_port, opcode_2_0_port, opcode_3_1_port, opcode_3_0_port, 
      opcode_4_1_port, opcode_4_0_port, opcode_5_1_port, opcode_5_0_port, 
      opcode_6_1_port, opcode_6_0_port, opcode_7_1_port, opcode_7_0_port, 
      opcode_8_1_port, opcode_8_0_port, opcode_9_1_port, opcode_9_0_port, 
      opcode_10_1_port, opcode_10_0_port, opcode_11_1_port, opcode_11_0_port, 
      opcode_12_1_port, opcode_12_0_port, opcode_13_1_port, opcode_13_0_port, 
      opcode_14_1_port, opcode_14_0_port, opcode_15_1_port, opcode_15_0_port, 
      opcode_16_1_port, opcode_16_0_port, opcode_17_1_port, opcode_17_0_port, 
      opcode_18_1_port, opcode_18_0_port, opcode_19_1_port, opcode_19_0_port, 
      opcode_20_1_port, opcode_20_0_port, opcode_21_1_port, opcode_21_0_port, 
      opcode_22_1_port, opcode_22_0_port, opcode_23_1_port, opcode_23_0_port, 
      opcode_24_1_port, opcode_24_0_port, opcode_25_1_port, opcode_25_0_port, 
      opcode_26_1_port, opcode_26_0_port, opcode_27_1_port, opcode_27_0_port, 
      opcode_28_1_port, opcode_28_0_port, opcode_29_1_port, opcode_29_0_port, 
      opcode_30_1_port, opcode_30_0_port, opcode_31_1_port, opcode_31_0_port, 
      memory_0_7_port, memory_0_6_port, memory_0_5_port, memory_0_4_port, 
      memory_0_3_port, memory_0_2_port, memory_0_1_port, memory_0_0_port, 
      memory_1_7_port, memory_1_6_port, memory_1_5_port, memory_1_4_port, 
      memory_1_3_port, memory_1_2_port, memory_1_1_port, memory_1_0_port, 
      memory_2_7_port, memory_2_6_port, memory_2_5_port, memory_2_4_port, 
      memory_2_3_port, memory_2_2_port, memory_2_1_port, memory_2_0_port, 
      memory_3_7_port, memory_3_6_port, memory_3_5_port, memory_3_4_port, 
      memory_3_3_port, memory_3_2_port, memory_3_1_port, memory_3_0_port, 
      memory_4_7_port, memory_4_6_port, memory_4_5_port, memory_4_4_port, 
      memory_4_3_port, memory_4_2_port, memory_4_1_port, memory_4_0_port, 
      memory_5_7_port, memory_5_6_port, memory_5_5_port, memory_5_4_port, 
      memory_5_3_port, memory_5_2_port, memory_5_1_port, memory_5_0_port, 
      memory_6_7_port, memory_6_6_port, memory_6_5_port, memory_6_4_port, 
      memory_6_3_port, memory_6_2_port, memory_6_1_port, memory_6_0_port, 
      memory_7_7_port, memory_7_6_port, memory_7_5_port, memory_7_4_port, 
      memory_7_3_port, memory_7_2_port, memory_7_1_port, memory_7_0_port, 
      memory_8_7_port, memory_8_6_port, memory_8_5_port, memory_8_4_port, 
      memory_8_3_port, memory_8_2_port, memory_8_1_port, memory_8_0_port, 
      memory_9_7_port, memory_9_6_port, memory_9_5_port, memory_9_4_port, 
      memory_9_3_port, memory_9_2_port, memory_9_1_port, memory_9_0_port, 
      memory_10_7_port, memory_10_6_port, memory_10_5_port, memory_10_4_port, 
      memory_10_3_port, memory_10_2_port, memory_10_1_port, memory_10_0_port, 
      memory_11_7_port, memory_11_6_port, memory_11_5_port, memory_11_4_port, 
      memory_11_3_port, memory_11_2_port, memory_11_1_port, memory_11_0_port, 
      memory_12_7_port, memory_12_6_port, memory_12_5_port, memory_12_4_port, 
      memory_12_3_port, memory_12_2_port, memory_12_1_port, memory_12_0_port, 
      memory_13_7_port, memory_13_6_port, memory_13_5_port, memory_13_4_port, 
      memory_13_3_port, memory_13_2_port, memory_13_1_port, memory_13_0_port, 
      memory_14_7_port, memory_14_6_port, memory_14_5_port, memory_14_4_port, 
      memory_14_3_port, memory_14_2_port, memory_14_1_port, memory_14_0_port, 
      memory_15_7_port, memory_15_6_port, memory_15_5_port, memory_15_4_port, 
      memory_15_3_port, memory_15_2_port, memory_15_1_port, memory_15_0_port, 
      memory_16_7_port, memory_16_6_port, memory_16_5_port, memory_16_4_port, 
      memory_16_3_port, memory_16_2_port, memory_16_1_port, memory_16_0_port, 
      memory_17_7_port, memory_17_6_port, memory_17_5_port, memory_17_4_port, 
      memory_17_3_port, memory_17_2_port, memory_17_1_port, memory_17_0_port, 
      memory_18_7_port, memory_18_6_port, memory_18_5_port, memory_18_4_port, 
      memory_18_3_port, memory_18_2_port, memory_18_1_port, memory_18_0_port, 
      memory_19_7_port, memory_19_6_port, memory_19_5_port, memory_19_4_port, 
      memory_19_3_port, memory_19_2_port, memory_19_1_port, memory_19_0_port, 
      memory_20_7_port, memory_20_6_port, memory_20_5_port, memory_20_4_port, 
      memory_20_3_port, memory_20_2_port, memory_20_1_port, memory_20_0_port, 
      memory_21_7_port, memory_21_6_port, memory_21_5_port, memory_21_4_port, 
      memory_21_3_port, memory_21_2_port, memory_21_1_port, memory_21_0_port, 
      memory_22_7_port, memory_22_6_port, memory_22_5_port, memory_22_4_port, 
      memory_22_3_port, memory_22_2_port, memory_22_1_port, memory_22_0_port, 
      memory_23_7_port, memory_23_6_port, memory_23_5_port, memory_23_4_port, 
      memory_23_3_port, memory_23_2_port, memory_23_1_port, memory_23_0_port, 
      memory_24_7_port, memory_24_6_port, memory_24_5_port, memory_24_4_port, 
      memory_24_3_port, memory_24_2_port, memory_24_1_port, memory_24_0_port, 
      memory_25_7_port, memory_25_6_port, memory_25_5_port, memory_25_4_port, 
      memory_25_3_port, memory_25_2_port, memory_25_1_port, memory_25_0_port, 
      memory_26_7_port, memory_26_6_port, memory_26_5_port, memory_26_4_port, 
      memory_26_3_port, memory_26_2_port, memory_26_1_port, memory_26_0_port, 
      memory_27_7_port, memory_27_6_port, memory_27_5_port, memory_27_4_port, 
      memory_27_3_port, memory_27_2_port, memory_27_1_port, memory_27_0_port, 
      memory_28_7_port, memory_28_6_port, memory_28_5_port, memory_28_4_port, 
      memory_28_3_port, memory_28_2_port, memory_28_1_port, memory_28_0_port, 
      memory_29_7_port, memory_29_6_port, memory_29_5_port, memory_29_4_port, 
      memory_29_3_port, memory_29_2_port, memory_29_1_port, memory_29_0_port, 
      memory_30_7_port, memory_30_6_port, memory_30_5_port, memory_30_4_port, 
      memory_30_3_port, memory_30_2_port, memory_30_1_port, memory_30_0_port, 
      memory_31_7_port, memory_31_6_port, memory_31_5_port, memory_31_4_port, 
      memory_31_3_port, memory_31_2_port, memory_31_1_port, memory_31_0_port, 
      N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, n847, n848, 
      n849, n850, n851, n853, n854, n855, n856, n857, n858, n859, n860, n861, 
      n862, n863, n864, n866, n867, n868, n869, n870, n871, n872, n873, n874, 
      n875, n876, n879, n880, n881, n882, n883, n884, n885, n886, n889, n890, 
      n891, n892, n893, n894, n895, n896, n899, n900, n901, n902, n903, n904, 
      n905, n906, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038
      , n1039, n1056, n1057, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
      n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, 
      n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, 
      n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
      n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, 
      n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, 
      n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, 
      n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, 
      n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, 
      n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1, n2, n3
      , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338_port, n339_port, n340_port, n341_port,
      n342_port, n343_port, n344_port, n345_port, n346_port, n347_port, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
      n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, 
      n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, 
      n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n852, n865, n877, n878, n887, n888, 
      n897, n898, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1168, 
      n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, 
      n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, 
      n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, 
      n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, 
      n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, 
      n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
      n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, 
      n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, 
      n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, 
      n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, 
      n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, 
      n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, 
      n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
      n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, 
      n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
      n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
      n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415 : std_logic;

begin
   DATA <= ( DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, 
      DATA_2_port, DATA_1_port, DATA_0_port );
   OUT_OPCODE <= ( OUT_OPCODE_1_port, OUT_OPCODE_0_port );
   EMPTY <= EMPTY_port;
   FULL <= FULL_port;
   
   X_Logic1_port <= '1';
   state_reg : DFFSR port map( D => X_Logic1_port, CLK => CLK, R => n177, S => 
                           n868, Q => state);
   readptr_reg_0_inst : DFFSR port map( D => N343, CLK => CLK, R => n177, S => 
                           n867, Q => readptr_0_port);
   readptr_reg_1_inst : DFFSR port map( D => N344, CLK => CLK, R => n177, S => 
                           n866, Q => readptr_1_port);
   readptr_reg_3_inst : DFFSR port map( D => N346, CLK => CLK, R => n177, S => 
                           n864, Q => readptr_3_port);
   readptr_reg_4_inst : DFFSR port map( D => N347, CLK => CLK, R => n177, S => 
                           n863, Q => readptr_4_port);
   writeptr_reg_4_inst : DFFSR port map( D => n862, CLK => CLK, R => n177, S =>
                           n861, Q => writeptr_4_port);
   writeptr_reg_3_inst : DFFSR port map( D => n860, CLK => CLK, R => n177, S =>
                           n859, Q => writeptr_3_port);
   writeptr_reg_0_inst : DFFSR port map( D => n858, CLK => CLK, R => n177, S =>
                           n857, Q => writeptr_0_port);
   writeptr_reg_1_inst : DFFSR port map( D => n856, CLK => CLK, R => n177, S =>
                           n855, Q => writeptr_1_port);
   writeptr_reg_2_inst : DFFSR port map( D => n854, CLK => CLK, R => n177, S =>
                           n853, Q => writeptr_2_port);
   FULL_reg : DFFPOSX1 port map( D => n1414, CLK => CLK, Q => FULL_port);
   BYTE_COUNT_reg_4_inst : DFFSR port map( D => N342, CLK => CLK, R => n177, S 
                           => n851, Q => BYTE_COUNT(4));
   BYTE_COUNT_reg_3_inst : DFFSR port map( D => N341, CLK => CLK, R => n177, S 
                           => n850, Q => BYTE_COUNT(3));
   BYTE_COUNT_reg_2_inst : DFFSR port map( D => N340, CLK => CLK, R => n177, S 
                           => n849, Q => BYTE_COUNT(2));
   BYTE_COUNT_reg_1_inst : DFFSR port map( D => N339, CLK => CLK, R => n177, S 
                           => n848, Q => BYTE_COUNT(1));
   BYTE_COUNT_reg_0_inst : DFFSR port map( D => N338, CLK => CLK, R => n177, S 
                           => n847, Q => BYTE_COUNT(0));
   memory_reg_0_7_inst : DFFPOSX1 port map( D => n1389, CLK => CLK, Q => 
                           memory_0_7_port);
   memory_reg_0_6_inst : DFFPOSX1 port map( D => n1388, CLK => CLK, Q => 
                           memory_0_6_port);
   memory_reg_0_5_inst : DFFPOSX1 port map( D => n1387, CLK => CLK, Q => 
                           memory_0_5_port);
   memory_reg_0_4_inst : DFFPOSX1 port map( D => n1386, CLK => CLK, Q => 
                           memory_0_4_port);
   memory_reg_0_3_inst : DFFPOSX1 port map( D => n1385, CLK => CLK, Q => 
                           memory_0_3_port);
   memory_reg_0_2_inst : DFFPOSX1 port map( D => n1384, CLK => CLK, Q => 
                           memory_0_2_port);
   memory_reg_0_1_inst : DFFPOSX1 port map( D => n1383, CLK => CLK, Q => 
                           memory_0_1_port);
   memory_reg_0_0_inst : DFFPOSX1 port map( D => n1382, CLK => CLK, Q => 
                           memory_0_0_port);
   memory_reg_1_7_inst : DFFPOSX1 port map( D => n1397, CLK => CLK, Q => 
                           memory_1_7_port);
   memory_reg_1_6_inst : DFFPOSX1 port map( D => n1396, CLK => CLK, Q => 
                           memory_1_6_port);
   memory_reg_1_5_inst : DFFPOSX1 port map( D => n1395, CLK => CLK, Q => 
                           memory_1_5_port);
   memory_reg_1_4_inst : DFFPOSX1 port map( D => n1394, CLK => CLK, Q => 
                           memory_1_4_port);
   memory_reg_1_3_inst : DFFPOSX1 port map( D => n1393, CLK => CLK, Q => 
                           memory_1_3_port);
   memory_reg_1_2_inst : DFFPOSX1 port map( D => n1392, CLK => CLK, Q => 
                           memory_1_2_port);
   memory_reg_1_1_inst : DFFPOSX1 port map( D => n1391, CLK => CLK, Q => 
                           memory_1_1_port);
   memory_reg_1_0_inst : DFFPOSX1 port map( D => n1390, CLK => CLK, Q => 
                           memory_1_0_port);
   memory_reg_2_7_inst : DFFPOSX1 port map( D => n1405, CLK => CLK, Q => 
                           memory_2_7_port);
   memory_reg_2_6_inst : DFFPOSX1 port map( D => n1404, CLK => CLK, Q => 
                           memory_2_6_port);
   memory_reg_2_5_inst : DFFPOSX1 port map( D => n1403, CLK => CLK, Q => 
                           memory_2_5_port);
   memory_reg_2_4_inst : DFFPOSX1 port map( D => n1402, CLK => CLK, Q => 
                           memory_2_4_port);
   memory_reg_2_3_inst : DFFPOSX1 port map( D => n1401, CLK => CLK, Q => 
                           memory_2_3_port);
   memory_reg_2_2_inst : DFFPOSX1 port map( D => n1400, CLK => CLK, Q => 
                           memory_2_2_port);
   memory_reg_2_1_inst : DFFPOSX1 port map( D => n1399, CLK => CLK, Q => 
                           memory_2_1_port);
   memory_reg_2_0_inst : DFFPOSX1 port map( D => n1398, CLK => CLK, Q => 
                           memory_2_0_port);
   memory_reg_3_7_inst : DFFPOSX1 port map( D => n1413, CLK => CLK, Q => 
                           memory_3_7_port);
   memory_reg_3_6_inst : DFFPOSX1 port map( D => n1412, CLK => CLK, Q => 
                           memory_3_6_port);
   memory_reg_3_5_inst : DFFPOSX1 port map( D => n1411, CLK => CLK, Q => 
                           memory_3_5_port);
   memory_reg_3_4_inst : DFFPOSX1 port map( D => n1410, CLK => CLK, Q => 
                           memory_3_4_port);
   memory_reg_3_3_inst : DFFPOSX1 port map( D => n1409, CLK => CLK, Q => 
                           memory_3_3_port);
   memory_reg_3_2_inst : DFFPOSX1 port map( D => n1408, CLK => CLK, Q => 
                           memory_3_2_port);
   memory_reg_3_1_inst : DFFPOSX1 port map( D => n1407, CLK => CLK, Q => 
                           memory_3_1_port);
   memory_reg_3_0_inst : DFFPOSX1 port map( D => n1406, CLK => CLK, Q => 
                           memory_3_0_port);
   memory_reg_4_7_inst : DFFPOSX1 port map( D => n869, CLK => CLK, Q => 
                           memory_4_7_port);
   memory_reg_4_6_inst : DFFPOSX1 port map( D => n870, CLK => CLK, Q => 
                           memory_4_6_port);
   memory_reg_4_5_inst : DFFPOSX1 port map( D => n871, CLK => CLK, Q => 
                           memory_4_5_port);
   memory_reg_4_4_inst : DFFPOSX1 port map( D => n872, CLK => CLK, Q => 
                           memory_4_4_port);
   memory_reg_4_3_inst : DFFPOSX1 port map( D => n873, CLK => CLK, Q => 
                           memory_4_3_port);
   memory_reg_4_2_inst : DFFPOSX1 port map( D => n874, CLK => CLK, Q => 
                           memory_4_2_port);
   memory_reg_4_1_inst : DFFPOSX1 port map( D => n875, CLK => CLK, Q => 
                           memory_4_1_port);
   memory_reg_4_0_inst : DFFPOSX1 port map( D => n876, CLK => CLK, Q => 
                           memory_4_0_port);
   memory_reg_5_7_inst : DFFPOSX1 port map( D => n879, CLK => CLK, Q => 
                           memory_5_7_port);
   memory_reg_5_6_inst : DFFPOSX1 port map( D => n880, CLK => CLK, Q => 
                           memory_5_6_port);
   memory_reg_5_5_inst : DFFPOSX1 port map( D => n881, CLK => CLK, Q => 
                           memory_5_5_port);
   memory_reg_5_4_inst : DFFPOSX1 port map( D => n882, CLK => CLK, Q => 
                           memory_5_4_port);
   memory_reg_5_3_inst : DFFPOSX1 port map( D => n883, CLK => CLK, Q => 
                           memory_5_3_port);
   memory_reg_5_2_inst : DFFPOSX1 port map( D => n884, CLK => CLK, Q => 
                           memory_5_2_port);
   memory_reg_5_1_inst : DFFPOSX1 port map( D => n885, CLK => CLK, Q => 
                           memory_5_1_port);
   memory_reg_5_0_inst : DFFPOSX1 port map( D => n886, CLK => CLK, Q => 
                           memory_5_0_port);
   memory_reg_6_7_inst : DFFPOSX1 port map( D => n889, CLK => CLK, Q => 
                           memory_6_7_port);
   memory_reg_6_6_inst : DFFPOSX1 port map( D => n890, CLK => CLK, Q => 
                           memory_6_6_port);
   memory_reg_6_5_inst : DFFPOSX1 port map( D => n891, CLK => CLK, Q => 
                           memory_6_5_port);
   memory_reg_6_4_inst : DFFPOSX1 port map( D => n892, CLK => CLK, Q => 
                           memory_6_4_port);
   memory_reg_6_3_inst : DFFPOSX1 port map( D => n893, CLK => CLK, Q => 
                           memory_6_3_port);
   memory_reg_6_2_inst : DFFPOSX1 port map( D => n894, CLK => CLK, Q => 
                           memory_6_2_port);
   memory_reg_6_1_inst : DFFPOSX1 port map( D => n895, CLK => CLK, Q => 
                           memory_6_1_port);
   memory_reg_6_0_inst : DFFPOSX1 port map( D => n896, CLK => CLK, Q => 
                           memory_6_0_port);
   memory_reg_7_7_inst : DFFPOSX1 port map( D => n899, CLK => CLK, Q => 
                           memory_7_7_port);
   memory_reg_7_6_inst : DFFPOSX1 port map( D => n900, CLK => CLK, Q => 
                           memory_7_6_port);
   memory_reg_7_5_inst : DFFPOSX1 port map( D => n901, CLK => CLK, Q => 
                           memory_7_5_port);
   memory_reg_7_4_inst : DFFPOSX1 port map( D => n902, CLK => CLK, Q => 
                           memory_7_4_port);
   memory_reg_7_3_inst : DFFPOSX1 port map( D => n903, CLK => CLK, Q => 
                           memory_7_3_port);
   memory_reg_7_2_inst : DFFPOSX1 port map( D => n904, CLK => CLK, Q => 
                           memory_7_2_port);
   memory_reg_7_1_inst : DFFPOSX1 port map( D => n905, CLK => CLK, Q => 
                           memory_7_1_port);
   memory_reg_7_0_inst : DFFPOSX1 port map( D => n906, CLK => CLK, Q => 
                           memory_7_0_port);
   memory_reg_8_7_inst : DFFPOSX1 port map( D => n1167, CLK => CLK, Q => 
                           memory_8_7_port);
   memory_reg_8_6_inst : DFFPOSX1 port map( D => n1166, CLK => CLK, Q => 
                           memory_8_6_port);
   memory_reg_8_5_inst : DFFPOSX1 port map( D => n1165, CLK => CLK, Q => 
                           memory_8_5_port);
   memory_reg_8_4_inst : DFFPOSX1 port map( D => n1164, CLK => CLK, Q => 
                           memory_8_4_port);
   memory_reg_8_3_inst : DFFPOSX1 port map( D => n1163, CLK => CLK, Q => 
                           memory_8_3_port);
   memory_reg_8_2_inst : DFFPOSX1 port map( D => n1162, CLK => CLK, Q => 
                           memory_8_2_port);
   memory_reg_8_1_inst : DFFPOSX1 port map( D => n1161, CLK => CLK, Q => 
                           memory_8_1_port);
   memory_reg_8_0_inst : DFFPOSX1 port map( D => n1160, CLK => CLK, Q => 
                           memory_8_0_port);
   memory_reg_9_7_inst : DFFPOSX1 port map( D => n1159, CLK => CLK, Q => 
                           memory_9_7_port);
   memory_reg_9_6_inst : DFFPOSX1 port map( D => n1158, CLK => CLK, Q => 
                           memory_9_6_port);
   memory_reg_9_5_inst : DFFPOSX1 port map( D => n1157, CLK => CLK, Q => 
                           memory_9_5_port);
   memory_reg_9_4_inst : DFFPOSX1 port map( D => n1156, CLK => CLK, Q => 
                           memory_9_4_port);
   memory_reg_9_3_inst : DFFPOSX1 port map( D => n1155, CLK => CLK, Q => 
                           memory_9_3_port);
   memory_reg_9_2_inst : DFFPOSX1 port map( D => n1154, CLK => CLK, Q => 
                           memory_9_2_port);
   memory_reg_9_1_inst : DFFPOSX1 port map( D => n1153, CLK => CLK, Q => 
                           memory_9_1_port);
   memory_reg_9_0_inst : DFFPOSX1 port map( D => n1152, CLK => CLK, Q => 
                           memory_9_0_port);
   memory_reg_10_7_inst : DFFPOSX1 port map( D => n1151, CLK => CLK, Q => 
                           memory_10_7_port);
   memory_reg_10_6_inst : DFFPOSX1 port map( D => n1150, CLK => CLK, Q => 
                           memory_10_6_port);
   memory_reg_10_5_inst : DFFPOSX1 port map( D => n1149, CLK => CLK, Q => 
                           memory_10_5_port);
   memory_reg_10_4_inst : DFFPOSX1 port map( D => n1148, CLK => CLK, Q => 
                           memory_10_4_port);
   memory_reg_10_3_inst : DFFPOSX1 port map( D => n1147, CLK => CLK, Q => 
                           memory_10_3_port);
   memory_reg_10_2_inst : DFFPOSX1 port map( D => n1146, CLK => CLK, Q => 
                           memory_10_2_port);
   memory_reg_10_1_inst : DFFPOSX1 port map( D => n1145, CLK => CLK, Q => 
                           memory_10_1_port);
   memory_reg_10_0_inst : DFFPOSX1 port map( D => n1144, CLK => CLK, Q => 
                           memory_10_0_port);
   memory_reg_11_7_inst : DFFPOSX1 port map( D => n1143, CLK => CLK, Q => 
                           memory_11_7_port);
   memory_reg_11_6_inst : DFFPOSX1 port map( D => n1142, CLK => CLK, Q => 
                           memory_11_6_port);
   memory_reg_11_5_inst : DFFPOSX1 port map( D => n1141, CLK => CLK, Q => 
                           memory_11_5_port);
   memory_reg_11_4_inst : DFFPOSX1 port map( D => n1140, CLK => CLK, Q => 
                           memory_11_4_port);
   memory_reg_11_3_inst : DFFPOSX1 port map( D => n1139, CLK => CLK, Q => 
                           memory_11_3_port);
   memory_reg_11_2_inst : DFFPOSX1 port map( D => n1138, CLK => CLK, Q => 
                           memory_11_2_port);
   memory_reg_11_1_inst : DFFPOSX1 port map( D => n1137, CLK => CLK, Q => 
                           memory_11_1_port);
   memory_reg_11_0_inst : DFFPOSX1 port map( D => n1136, CLK => CLK, Q => 
                           memory_11_0_port);
   memory_reg_12_7_inst : DFFPOSX1 port map( D => n1374, CLK => CLK, Q => 
                           memory_12_7_port);
   memory_reg_12_6_inst : DFFPOSX1 port map( D => n1375, CLK => CLK, Q => 
                           memory_12_6_port);
   memory_reg_12_5_inst : DFFPOSX1 port map( D => n1376, CLK => CLK, Q => 
                           memory_12_5_port);
   memory_reg_12_4_inst : DFFPOSX1 port map( D => n1377, CLK => CLK, Q => 
                           memory_12_4_port);
   memory_reg_12_3_inst : DFFPOSX1 port map( D => n1378, CLK => CLK, Q => 
                           memory_12_3_port);
   memory_reg_12_2_inst : DFFPOSX1 port map( D => n1379, CLK => CLK, Q => 
                           memory_12_2_port);
   memory_reg_12_1_inst : DFFPOSX1 port map( D => n1380, CLK => CLK, Q => 
                           memory_12_1_port);
   memory_reg_12_0_inst : DFFPOSX1 port map( D => n1381, CLK => CLK, Q => 
                           memory_12_0_port);
   memory_reg_13_7_inst : DFFPOSX1 port map( D => n1366, CLK => CLK, Q => 
                           memory_13_7_port);
   memory_reg_13_6_inst : DFFPOSX1 port map( D => n1367, CLK => CLK, Q => 
                           memory_13_6_port);
   memory_reg_13_5_inst : DFFPOSX1 port map( D => n1368, CLK => CLK, Q => 
                           memory_13_5_port);
   memory_reg_13_4_inst : DFFPOSX1 port map( D => n1369, CLK => CLK, Q => 
                           memory_13_4_port);
   memory_reg_13_3_inst : DFFPOSX1 port map( D => n1370, CLK => CLK, Q => 
                           memory_13_3_port);
   memory_reg_13_2_inst : DFFPOSX1 port map( D => n1371, CLK => CLK, Q => 
                           memory_13_2_port);
   memory_reg_13_1_inst : DFFPOSX1 port map( D => n1372, CLK => CLK, Q => 
                           memory_13_1_port);
   memory_reg_13_0_inst : DFFPOSX1 port map( D => n1373, CLK => CLK, Q => 
                           memory_13_0_port);
   memory_reg_14_7_inst : DFFPOSX1 port map( D => n1358, CLK => CLK, Q => 
                           memory_14_7_port);
   memory_reg_14_6_inst : DFFPOSX1 port map( D => n1359, CLK => CLK, Q => 
                           memory_14_6_port);
   memory_reg_14_5_inst : DFFPOSX1 port map( D => n1360, CLK => CLK, Q => 
                           memory_14_5_port);
   memory_reg_14_4_inst : DFFPOSX1 port map( D => n1361, CLK => CLK, Q => 
                           memory_14_4_port);
   memory_reg_14_3_inst : DFFPOSX1 port map( D => n1362, CLK => CLK, Q => 
                           memory_14_3_port);
   memory_reg_14_2_inst : DFFPOSX1 port map( D => n1363, CLK => CLK, Q => 
                           memory_14_2_port);
   memory_reg_14_1_inst : DFFPOSX1 port map( D => n1364, CLK => CLK, Q => 
                           memory_14_1_port);
   memory_reg_14_0_inst : DFFPOSX1 port map( D => n1365, CLK => CLK, Q => 
                           memory_14_0_port);
   memory_reg_15_7_inst : DFFPOSX1 port map( D => n1350, CLK => CLK, Q => 
                           memory_15_7_port);
   memory_reg_15_6_inst : DFFPOSX1 port map( D => n1351, CLK => CLK, Q => 
                           memory_15_6_port);
   memory_reg_15_5_inst : DFFPOSX1 port map( D => n1352, CLK => CLK, Q => 
                           memory_15_5_port);
   memory_reg_15_4_inst : DFFPOSX1 port map( D => n1353, CLK => CLK, Q => 
                           memory_15_4_port);
   memory_reg_15_3_inst : DFFPOSX1 port map( D => n1354, CLK => CLK, Q => 
                           memory_15_3_port);
   memory_reg_15_2_inst : DFFPOSX1 port map( D => n1355, CLK => CLK, Q => 
                           memory_15_2_port);
   memory_reg_15_1_inst : DFFPOSX1 port map( D => n1356, CLK => CLK, Q => 
                           memory_15_1_port);
   memory_reg_15_0_inst : DFFPOSX1 port map( D => n1357, CLK => CLK, Q => 
                           memory_15_0_port);
   memory_reg_16_7_inst : DFFPOSX1 port map( D => n1135, CLK => CLK, Q => 
                           memory_16_7_port);
   memory_reg_16_6_inst : DFFPOSX1 port map( D => n1134, CLK => CLK, Q => 
                           memory_16_6_port);
   memory_reg_16_5_inst : DFFPOSX1 port map( D => n1133, CLK => CLK, Q => 
                           memory_16_5_port);
   memory_reg_16_4_inst : DFFPOSX1 port map( D => n1132, CLK => CLK, Q => 
                           memory_16_4_port);
   memory_reg_16_3_inst : DFFPOSX1 port map( D => n1131, CLK => CLK, Q => 
                           memory_16_3_port);
   memory_reg_16_2_inst : DFFPOSX1 port map( D => n1130, CLK => CLK, Q => 
                           memory_16_2_port);
   memory_reg_16_1_inst : DFFPOSX1 port map( D => n1129, CLK => CLK, Q => 
                           memory_16_1_port);
   memory_reg_16_0_inst : DFFPOSX1 port map( D => n1128, CLK => CLK, Q => 
                           memory_16_0_port);
   memory_reg_17_7_inst : DFFPOSX1 port map( D => n1127, CLK => CLK, Q => 
                           memory_17_7_port);
   memory_reg_17_6_inst : DFFPOSX1 port map( D => n1126, CLK => CLK, Q => 
                           memory_17_6_port);
   memory_reg_17_5_inst : DFFPOSX1 port map( D => n1125, CLK => CLK, Q => 
                           memory_17_5_port);
   memory_reg_17_4_inst : DFFPOSX1 port map( D => n1124, CLK => CLK, Q => 
                           memory_17_4_port);
   memory_reg_17_3_inst : DFFPOSX1 port map( D => n1123, CLK => CLK, Q => 
                           memory_17_3_port);
   memory_reg_17_2_inst : DFFPOSX1 port map( D => n1122, CLK => CLK, Q => 
                           memory_17_2_port);
   memory_reg_17_1_inst : DFFPOSX1 port map( D => n1121, CLK => CLK, Q => 
                           memory_17_1_port);
   memory_reg_17_0_inst : DFFPOSX1 port map( D => n1120, CLK => CLK, Q => 
                           memory_17_0_port);
   memory_reg_18_7_inst : DFFPOSX1 port map( D => n1119, CLK => CLK, Q => 
                           memory_18_7_port);
   memory_reg_18_6_inst : DFFPOSX1 port map( D => n1118, CLK => CLK, Q => 
                           memory_18_6_port);
   memory_reg_18_5_inst : DFFPOSX1 port map( D => n1117, CLK => CLK, Q => 
                           memory_18_5_port);
   memory_reg_18_4_inst : DFFPOSX1 port map( D => n1116, CLK => CLK, Q => 
                           memory_18_4_port);
   memory_reg_18_3_inst : DFFPOSX1 port map( D => n1115, CLK => CLK, Q => 
                           memory_18_3_port);
   memory_reg_18_2_inst : DFFPOSX1 port map( D => n1114, CLK => CLK, Q => 
                           memory_18_2_port);
   memory_reg_18_1_inst : DFFPOSX1 port map( D => n1113, CLK => CLK, Q => 
                           memory_18_1_port);
   memory_reg_18_0_inst : DFFPOSX1 port map( D => n1112, CLK => CLK, Q => 
                           memory_18_0_port);
   memory_reg_19_7_inst : DFFPOSX1 port map( D => n1111, CLK => CLK, Q => 
                           memory_19_7_port);
   memory_reg_19_6_inst : DFFPOSX1 port map( D => n1110, CLK => CLK, Q => 
                           memory_19_6_port);
   memory_reg_19_5_inst : DFFPOSX1 port map( D => n1109, CLK => CLK, Q => 
                           memory_19_5_port);
   memory_reg_19_4_inst : DFFPOSX1 port map( D => n1108, CLK => CLK, Q => 
                           memory_19_4_port);
   memory_reg_19_3_inst : DFFPOSX1 port map( D => n1107, CLK => CLK, Q => 
                           memory_19_3_port);
   memory_reg_19_2_inst : DFFPOSX1 port map( D => n1106, CLK => CLK, Q => 
                           memory_19_2_port);
   memory_reg_19_1_inst : DFFPOSX1 port map( D => n1105, CLK => CLK, Q => 
                           memory_19_1_port);
   memory_reg_19_0_inst : DFFPOSX1 port map( D => n1104, CLK => CLK, Q => 
                           memory_19_0_port);
   memory_reg_20_7_inst : DFFPOSX1 port map( D => n1342, CLK => CLK, Q => 
                           memory_20_7_port);
   memory_reg_20_6_inst : DFFPOSX1 port map( D => n1343, CLK => CLK, Q => 
                           memory_20_6_port);
   memory_reg_20_5_inst : DFFPOSX1 port map( D => n1344, CLK => CLK, Q => 
                           memory_20_5_port);
   memory_reg_20_4_inst : DFFPOSX1 port map( D => n1345, CLK => CLK, Q => 
                           memory_20_4_port);
   memory_reg_20_3_inst : DFFPOSX1 port map( D => n1346, CLK => CLK, Q => 
                           memory_20_3_port);
   memory_reg_20_2_inst : DFFPOSX1 port map( D => n1347, CLK => CLK, Q => 
                           memory_20_2_port);
   memory_reg_20_1_inst : DFFPOSX1 port map( D => n1348, CLK => CLK, Q => 
                           memory_20_1_port);
   memory_reg_20_0_inst : DFFPOSX1 port map( D => n1349, CLK => CLK, Q => 
                           memory_20_0_port);
   memory_reg_21_7_inst : DFFPOSX1 port map( D => n1334, CLK => CLK, Q => 
                           memory_21_7_port);
   memory_reg_21_6_inst : DFFPOSX1 port map( D => n1335, CLK => CLK, Q => 
                           memory_21_6_port);
   memory_reg_21_5_inst : DFFPOSX1 port map( D => n1336, CLK => CLK, Q => 
                           memory_21_5_port);
   memory_reg_21_4_inst : DFFPOSX1 port map( D => n1337, CLK => CLK, Q => 
                           memory_21_4_port);
   memory_reg_21_3_inst : DFFPOSX1 port map( D => n1338, CLK => CLK, Q => 
                           memory_21_3_port);
   memory_reg_21_2_inst : DFFPOSX1 port map( D => n1339, CLK => CLK, Q => 
                           memory_21_2_port);
   memory_reg_21_1_inst : DFFPOSX1 port map( D => n1340, CLK => CLK, Q => 
                           memory_21_1_port);
   memory_reg_21_0_inst : DFFPOSX1 port map( D => n1341, CLK => CLK, Q => 
                           memory_21_0_port);
   memory_reg_22_7_inst : DFFPOSX1 port map( D => n1326, CLK => CLK, Q => 
                           memory_22_7_port);
   memory_reg_22_6_inst : DFFPOSX1 port map( D => n1327, CLK => CLK, Q => 
                           memory_22_6_port);
   memory_reg_22_5_inst : DFFPOSX1 port map( D => n1328, CLK => CLK, Q => 
                           memory_22_5_port);
   memory_reg_22_4_inst : DFFPOSX1 port map( D => n1329, CLK => CLK, Q => 
                           memory_22_4_port);
   memory_reg_22_3_inst : DFFPOSX1 port map( D => n1330, CLK => CLK, Q => 
                           memory_22_3_port);
   memory_reg_22_2_inst : DFFPOSX1 port map( D => n1331, CLK => CLK, Q => 
                           memory_22_2_port);
   memory_reg_22_1_inst : DFFPOSX1 port map( D => n1332, CLK => CLK, Q => 
                           memory_22_1_port);
   memory_reg_22_0_inst : DFFPOSX1 port map( D => n1333, CLK => CLK, Q => 
                           memory_22_0_port);
   memory_reg_23_7_inst : DFFPOSX1 port map( D => n1318, CLK => CLK, Q => 
                           memory_23_7_port);
   memory_reg_23_6_inst : DFFPOSX1 port map( D => n1319, CLK => CLK, Q => 
                           memory_23_6_port);
   memory_reg_23_5_inst : DFFPOSX1 port map( D => n1320, CLK => CLK, Q => 
                           memory_23_5_port);
   memory_reg_23_4_inst : DFFPOSX1 port map( D => n1321, CLK => CLK, Q => 
                           memory_23_4_port);
   memory_reg_23_3_inst : DFFPOSX1 port map( D => n1322, CLK => CLK, Q => 
                           memory_23_3_port);
   memory_reg_23_2_inst : DFFPOSX1 port map( D => n1323, CLK => CLK, Q => 
                           memory_23_2_port);
   memory_reg_23_1_inst : DFFPOSX1 port map( D => n1324, CLK => CLK, Q => 
                           memory_23_1_port);
   memory_reg_23_0_inst : DFFPOSX1 port map( D => n1325, CLK => CLK, Q => 
                           memory_23_0_port);
   memory_reg_24_7_inst : DFFPOSX1 port map( D => n1310, CLK => CLK, Q => 
                           memory_24_7_port);
   memory_reg_24_6_inst : DFFPOSX1 port map( D => n1311, CLK => CLK, Q => 
                           memory_24_6_port);
   memory_reg_24_5_inst : DFFPOSX1 port map( D => n1312, CLK => CLK, Q => 
                           memory_24_5_port);
   memory_reg_24_4_inst : DFFPOSX1 port map( D => n1313, CLK => CLK, Q => 
                           memory_24_4_port);
   memory_reg_24_3_inst : DFFPOSX1 port map( D => n1314, CLK => CLK, Q => 
                           memory_24_3_port);
   memory_reg_24_2_inst : DFFPOSX1 port map( D => n1315, CLK => CLK, Q => 
                           memory_24_2_port);
   memory_reg_24_1_inst : DFFPOSX1 port map( D => n1316, CLK => CLK, Q => 
                           memory_24_1_port);
   memory_reg_24_0_inst : DFFPOSX1 port map( D => n1317, CLK => CLK, Q => 
                           memory_24_0_port);
   memory_reg_25_7_inst : DFFPOSX1 port map( D => n1302, CLK => CLK, Q => 
                           memory_25_7_port);
   memory_reg_25_6_inst : DFFPOSX1 port map( D => n1303, CLK => CLK, Q => 
                           memory_25_6_port);
   memory_reg_25_5_inst : DFFPOSX1 port map( D => n1304, CLK => CLK, Q => 
                           memory_25_5_port);
   memory_reg_25_4_inst : DFFPOSX1 port map( D => n1305, CLK => CLK, Q => 
                           memory_25_4_port);
   memory_reg_25_3_inst : DFFPOSX1 port map( D => n1306, CLK => CLK, Q => 
                           memory_25_3_port);
   memory_reg_25_2_inst : DFFPOSX1 port map( D => n1307, CLK => CLK, Q => 
                           memory_25_2_port);
   memory_reg_25_1_inst : DFFPOSX1 port map( D => n1308, CLK => CLK, Q => 
                           memory_25_1_port);
   memory_reg_25_0_inst : DFFPOSX1 port map( D => n1309, CLK => CLK, Q => 
                           memory_25_0_port);
   memory_reg_26_7_inst : DFFPOSX1 port map( D => n1294, CLK => CLK, Q => 
                           memory_26_7_port);
   memory_reg_26_6_inst : DFFPOSX1 port map( D => n1295, CLK => CLK, Q => 
                           memory_26_6_port);
   memory_reg_26_5_inst : DFFPOSX1 port map( D => n1296, CLK => CLK, Q => 
                           memory_26_5_port);
   memory_reg_26_4_inst : DFFPOSX1 port map( D => n1297, CLK => CLK, Q => 
                           memory_26_4_port);
   memory_reg_26_3_inst : DFFPOSX1 port map( D => n1298, CLK => CLK, Q => 
                           memory_26_3_port);
   memory_reg_26_2_inst : DFFPOSX1 port map( D => n1299, CLK => CLK, Q => 
                           memory_26_2_port);
   memory_reg_26_1_inst : DFFPOSX1 port map( D => n1300, CLK => CLK, Q => 
                           memory_26_1_port);
   memory_reg_26_0_inst : DFFPOSX1 port map( D => n1301, CLK => CLK, Q => 
                           memory_26_0_port);
   memory_reg_27_7_inst : DFFPOSX1 port map( D => n1286, CLK => CLK, Q => 
                           memory_27_7_port);
   memory_reg_27_6_inst : DFFPOSX1 port map( D => n1287, CLK => CLK, Q => 
                           memory_27_6_port);
   memory_reg_27_5_inst : DFFPOSX1 port map( D => n1288, CLK => CLK, Q => 
                           memory_27_5_port);
   memory_reg_27_4_inst : DFFPOSX1 port map( D => n1289, CLK => CLK, Q => 
                           memory_27_4_port);
   memory_reg_27_3_inst : DFFPOSX1 port map( D => n1290, CLK => CLK, Q => 
                           memory_27_3_port);
   memory_reg_27_2_inst : DFFPOSX1 port map( D => n1291, CLK => CLK, Q => 
                           memory_27_2_port);
   memory_reg_27_1_inst : DFFPOSX1 port map( D => n1292, CLK => CLK, Q => 
                           memory_27_1_port);
   memory_reg_27_0_inst : DFFPOSX1 port map( D => n1293, CLK => CLK, Q => 
                           memory_27_0_port);
   memory_reg_28_7_inst : DFFPOSX1 port map( D => n1103, CLK => CLK, Q => 
                           memory_28_7_port);
   memory_reg_28_6_inst : DFFPOSX1 port map( D => n1102, CLK => CLK, Q => 
                           memory_28_6_port);
   memory_reg_28_5_inst : DFFPOSX1 port map( D => n1101, CLK => CLK, Q => 
                           memory_28_5_port);
   memory_reg_28_4_inst : DFFPOSX1 port map( D => n1100, CLK => CLK, Q => 
                           memory_28_4_port);
   memory_reg_28_3_inst : DFFPOSX1 port map( D => n1099, CLK => CLK, Q => 
                           memory_28_3_port);
   memory_reg_28_2_inst : DFFPOSX1 port map( D => n1098, CLK => CLK, Q => 
                           memory_28_2_port);
   memory_reg_28_1_inst : DFFPOSX1 port map( D => n1097, CLK => CLK, Q => 
                           memory_28_1_port);
   memory_reg_28_0_inst : DFFPOSX1 port map( D => n1096, CLK => CLK, Q => 
                           memory_28_0_port);
   memory_reg_29_7_inst : DFFPOSX1 port map( D => n1095, CLK => CLK, Q => 
                           memory_29_7_port);
   memory_reg_29_6_inst : DFFPOSX1 port map( D => n1094, CLK => CLK, Q => 
                           memory_29_6_port);
   memory_reg_29_5_inst : DFFPOSX1 port map( D => n1093, CLK => CLK, Q => 
                           memory_29_5_port);
   memory_reg_29_4_inst : DFFPOSX1 port map( D => n1092, CLK => CLK, Q => 
                           memory_29_4_port);
   memory_reg_29_3_inst : DFFPOSX1 port map( D => n1091, CLK => CLK, Q => 
                           memory_29_3_port);
   memory_reg_29_2_inst : DFFPOSX1 port map( D => n1090, CLK => CLK, Q => 
                           memory_29_2_port);
   memory_reg_29_1_inst : DFFPOSX1 port map( D => n1089, CLK => CLK, Q => 
                           memory_29_1_port);
   memory_reg_29_0_inst : DFFPOSX1 port map( D => n1088, CLK => CLK, Q => 
                           memory_29_0_port);
   memory_reg_30_7_inst : DFFPOSX1 port map( D => n1087, CLK => CLK, Q => 
                           memory_30_7_port);
   memory_reg_30_6_inst : DFFPOSX1 port map( D => n1086, CLK => CLK, Q => 
                           memory_30_6_port);
   memory_reg_30_5_inst : DFFPOSX1 port map( D => n1085, CLK => CLK, Q => 
                           memory_30_5_port);
   memory_reg_30_4_inst : DFFPOSX1 port map( D => n1084, CLK => CLK, Q => 
                           memory_30_4_port);
   memory_reg_30_3_inst : DFFPOSX1 port map( D => n1083, CLK => CLK, Q => 
                           memory_30_3_port);
   memory_reg_30_2_inst : DFFPOSX1 port map( D => n1082, CLK => CLK, Q => 
                           memory_30_2_port);
   memory_reg_30_1_inst : DFFPOSX1 port map( D => n1081, CLK => CLK, Q => 
                           memory_30_1_port);
   memory_reg_30_0_inst : DFFPOSX1 port map( D => n1080, CLK => CLK, Q => 
                           memory_30_0_port);
   memory_reg_31_7_inst : DFFPOSX1 port map( D => n1079, CLK => CLK, Q => 
                           memory_31_7_port);
   memory_reg_31_6_inst : DFFPOSX1 port map( D => n1078, CLK => CLK, Q => 
                           memory_31_6_port);
   memory_reg_31_5_inst : DFFPOSX1 port map( D => n1077, CLK => CLK, Q => 
                           memory_31_5_port);
   memory_reg_31_4_inst : DFFPOSX1 port map( D => n1076, CLK => CLK, Q => 
                           memory_31_4_port);
   memory_reg_31_3_inst : DFFPOSX1 port map( D => n1075, CLK => CLK, Q => 
                           memory_31_3_port);
   memory_reg_31_2_inst : DFFPOSX1 port map( D => n1074, CLK => CLK, Q => 
                           memory_31_2_port);
   memory_reg_31_1_inst : DFFPOSX1 port map( D => n1073, CLK => CLK, Q => 
                           memory_31_1_port);
   memory_reg_31_0_inst : DFFPOSX1 port map( D => n1072, CLK => CLK, Q => 
                           memory_31_0_port);
   opcode_reg_0_1_inst : DFFPOSX1 port map( D => n610, CLK => CLK, Q => 
                           opcode_0_1_port);
   opcode_reg_0_0_inst : DFFPOSX1 port map( D => n611, CLK => CLK, Q => 
                           opcode_0_0_port);
   opcode_reg_1_1_inst : DFFPOSX1 port map( D => n652, CLK => CLK, Q => 
                           opcode_1_1_port);
   opcode_reg_1_0_inst : DFFPOSX1 port map( D => n653, CLK => CLK, Q => 
                           opcode_1_0_port);
   opcode_reg_2_1_inst : DFFPOSX1 port map( D => n654, CLK => CLK, Q => 
                           opcode_2_1_port);
   opcode_reg_2_0_inst : DFFPOSX1 port map( D => n655, CLK => CLK, Q => 
                           opcode_2_0_port);
   opcode_reg_3_1_inst : DFFPOSX1 port map( D => n624, CLK => CLK, Q => 
                           opcode_3_1_port);
   opcode_reg_3_0_inst : DFFPOSX1 port map( D => n625, CLK => CLK, Q => 
                           opcode_3_0_port);
   opcode_reg_4_1_inst : DFFPOSX1 port map( D => n640, CLK => CLK, Q => 
                           opcode_4_1_port);
   opcode_reg_4_0_inst : DFFPOSX1 port map( D => n641, CLK => CLK, Q => 
                           opcode_4_0_port);
   opcode_reg_5_1_inst : DFFPOSX1 port map( D => n614, CLK => CLK, Q => 
                           opcode_5_1_port);
   opcode_reg_5_0_inst : DFFPOSX1 port map( D => n615, CLK => CLK, Q => 
                           opcode_5_0_port);
   opcode_reg_6_1_inst : DFFPOSX1 port map( D => n600, CLK => CLK, Q => 
                           opcode_6_1_port);
   opcode_reg_6_0_inst : DFFPOSX1 port map( D => n601, CLK => CLK, Q => 
                           opcode_6_0_port);
   opcode_reg_7_1_inst : DFFPOSX1 port map( D => n608, CLK => CLK, Q => 
                           opcode_7_1_port);
   opcode_reg_7_0_inst : DFFPOSX1 port map( D => n609, CLK => CLK, Q => 
                           opcode_7_0_port);
   opcode_reg_8_1_inst : DFFPOSX1 port map( D => n634, CLK => CLK, Q => 
                           opcode_8_1_port);
   opcode_reg_8_0_inst : DFFPOSX1 port map( D => n635, CLK => CLK, Q => 
                           opcode_8_0_port);
   opcode_reg_9_1_inst : DFFPOSX1 port map( D => n622, CLK => CLK, Q => 
                           opcode_9_1_port);
   opcode_reg_9_0_inst : DFFPOSX1 port map( D => n623, CLK => CLK, Q => 
                           opcode_9_0_port);
   opcode_reg_10_1_inst : DFFPOSX1 port map( D => n646, CLK => CLK, Q => 
                           opcode_10_1_port);
   opcode_reg_10_0_inst : DFFPOSX1 port map( D => n647, CLK => CLK, Q => 
                           opcode_10_0_port);
   opcode_reg_11_1_inst : DFFPOSX1 port map( D => n1057, CLK => CLK, Q => 
                           opcode_11_1_port);
   opcode_reg_11_0_inst : DFFPOSX1 port map( D => n1056, CLK => CLK, Q => 
                           opcode_11_0_port);
   opcode_reg_12_1_inst : DFFPOSX1 port map( D => n642, CLK => CLK, Q => 
                           opcode_12_1_port);
   opcode_reg_12_0_inst : DFFPOSX1 port map( D => n643, CLK => CLK, Q => 
                           opcode_12_0_port);
   opcode_reg_13_1_inst : DFFPOSX1 port map( D => n638, CLK => CLK, Q => 
                           opcode_13_1_port);
   opcode_reg_13_0_inst : DFFPOSX1 port map( D => n639, CLK => CLK, Q => 
                           opcode_13_0_port);
   opcode_reg_14_1_inst : DFFPOSX1 port map( D => n636, CLK => CLK, Q => 
                           opcode_14_1_port);
   opcode_reg_14_0_inst : DFFPOSX1 port map( D => n637, CLK => CLK, Q => 
                           opcode_14_0_port);
   opcode_reg_15_1_inst : DFFPOSX1 port map( D => n648, CLK => CLK, Q => 
                           opcode_15_1_port);
   opcode_reg_15_0_inst : DFFPOSX1 port map( D => n649, CLK => CLK, Q => 
                           opcode_15_0_port);
   opcode_reg_16_1_inst : DFFPOSX1 port map( D => n626, CLK => CLK, Q => 
                           opcode_16_1_port);
   opcode_reg_16_0_inst : DFFPOSX1 port map( D => n627, CLK => CLK, Q => 
                           opcode_16_0_port);
   opcode_reg_17_1_inst : DFFPOSX1 port map( D => n612, CLK => CLK, Q => 
                           opcode_17_1_port);
   opcode_reg_17_0_inst : DFFPOSX1 port map( D => n613, CLK => CLK, Q => 
                           opcode_17_0_port);
   opcode_reg_18_1_inst : DFFPOSX1 port map( D => n602, CLK => CLK, Q => 
                           opcode_18_1_port);
   opcode_reg_18_0_inst : DFFPOSX1 port map( D => n603, CLK => CLK, Q => 
                           opcode_18_0_port);
   opcode_reg_19_1_inst : DFFPOSX1 port map( D => n628, CLK => CLK, Q => 
                           opcode_19_1_port);
   opcode_reg_19_0_inst : DFFPOSX1 port map( D => n629, CLK => CLK, Q => 
                           opcode_19_0_port);
   opcode_reg_20_1_inst : DFFPOSX1 port map( D => n658, CLK => CLK, Q => 
                           opcode_20_1_port);
   opcode_reg_20_0_inst : DFFPOSX1 port map( D => n659, CLK => CLK, Q => 
                           opcode_20_0_port);
   opcode_reg_21_1_inst : DFFPOSX1 port map( D => n660, CLK => CLK, Q => 
                           opcode_21_1_port);
   opcode_reg_21_0_inst : DFFPOSX1 port map( D => n661, CLK => CLK, Q => 
                           opcode_21_0_port);
   opcode_reg_22_1_inst : DFFPOSX1 port map( D => n620, CLK => CLK, Q => 
                           opcode_22_1_port);
   opcode_reg_22_0_inst : DFFPOSX1 port map( D => n621, CLK => CLK, Q => 
                           opcode_22_0_port);
   opcode_reg_23_1_inst : DFFPOSX1 port map( D => n618, CLK => CLK, Q => 
                           opcode_23_1_port);
   opcode_reg_23_0_inst : DFFPOSX1 port map( D => n619, CLK => CLK, Q => 
                           opcode_23_0_port);
   opcode_reg_24_1_inst : DFFPOSX1 port map( D => n606, CLK => CLK, Q => 
                           opcode_24_1_port);
   opcode_reg_24_0_inst : DFFPOSX1 port map( D => n607, CLK => CLK, Q => 
                           opcode_24_0_port);
   opcode_reg_25_1_inst : DFFPOSX1 port map( D => n656, CLK => CLK, Q => 
                           opcode_25_1_port);
   opcode_reg_25_0_inst : DFFPOSX1 port map( D => n657, CLK => CLK, Q => 
                           opcode_25_0_port);
   opcode_reg_26_1_inst : DFFPOSX1 port map( D => n630, CLK => CLK, Q => 
                           opcode_26_1_port);
   opcode_reg_26_0_inst : DFFPOSX1 port map( D => n631, CLK => CLK, Q => 
                           opcode_26_0_port);
   opcode_reg_27_1_inst : DFFPOSX1 port map( D => n650, CLK => CLK, Q => 
                           opcode_27_1_port);
   opcode_reg_27_0_inst : DFFPOSX1 port map( D => n651, CLK => CLK, Q => 
                           opcode_27_0_port);
   opcode_reg_28_1_inst : DFFPOSX1 port map( D => n644, CLK => CLK, Q => 
                           opcode_28_1_port);
   opcode_reg_28_0_inst : DFFPOSX1 port map( D => n645, CLK => CLK, Q => 
                           opcode_28_0_port);
   opcode_reg_29_1_inst : DFFPOSX1 port map( D => n632, CLK => CLK, Q => 
                           opcode_29_1_port);
   opcode_reg_29_0_inst : DFFPOSX1 port map( D => n633, CLK => CLK, Q => 
                           opcode_29_0_port);
   opcode_reg_30_1_inst : DFFPOSX1 port map( D => n616, CLK => CLK, Q => 
                           opcode_30_1_port);
   opcode_reg_30_0_inst : DFFPOSX1 port map( D => n617, CLK => CLK, Q => 
                           opcode_30_0_port);
   opcode_reg_31_1_inst : DFFPOSX1 port map( D => n604, CLK => CLK, Q => 
                           opcode_31_1_port);
   opcode_reg_31_0_inst : DFFPOSX1 port map( D => n605, CLK => CLK, Q => 
                           opcode_31_0_port);
   DATA_reg_7_inst : DFFPOSX1 port map( D => n1039, CLK => CLK, Q => 
                           DATA_7_port);
   DATA_reg_6_inst : DFFPOSX1 port map( D => n1038, CLK => CLK, Q => 
                           DATA_6_port);
   DATA_reg_5_inst : DFFPOSX1 port map( D => n1037, CLK => CLK, Q => 
                           DATA_5_port);
   DATA_reg_4_inst : DFFPOSX1 port map( D => n1036, CLK => CLK, Q => 
                           DATA_4_port);
   DATA_reg_3_inst : DFFPOSX1 port map( D => n1035, CLK => CLK, Q => 
                           DATA_3_port);
   DATA_reg_2_inst : DFFPOSX1 port map( D => n1034, CLK => CLK, Q => 
                           DATA_2_port);
   DATA_reg_1_inst : DFFPOSX1 port map( D => n1033, CLK => CLK, Q => 
                           DATA_1_port);
   DATA_reg_0_inst : DFFPOSX1 port map( D => n1032, CLK => CLK, Q => 
                           DATA_0_port);
   OUT_OPCODE_reg_1_inst : DFFPOSX1 port map( D => n1031, CLK => CLK, Q => 
                           OUT_OPCODE_1_port);
   OUT_OPCODE_reg_0_inst : DFFPOSX1 port map( D => n1030, CLK => CLK, Q => 
                           OUT_OPCODE_0_port);
   EMPTY_reg : DFFPOSX1 port map( D => n1415, CLK => CLK, Q => EMPTY_port);
   n847 <= '1';
   n848 <= '1';
   n849 <= '1';
   n850 <= '1';
   n851 <= '1';
   n853 <= '1';
   n855 <= '1';
   n857 <= '1';
   n859 <= '1';
   n861 <= '1';
   n863 <= '1';
   n864 <= '1';
   n866 <= '1';
   n867 <= '1';
   n868 <= '1';
   readptr_reg_2_inst : DFFSR port map( D => N345, CLK => CLK, R => n177, S => 
                           n23, Q => readptr_2_port);
   U3 : INVX1 port map( A => n94, Y => n568);
   U4 : INVX4 port map( A => n50, Y => n51);
   U5 : INVX2 port map( A => n338_port, Y => n512);
   U6 : INVX2 port map( A => n348, Y => n514);
   U7 : INVX2 port map( A => n248, Y => n1);
   U8 : INVX2 port map( A => n248, Y => n33);
   U9 : AND2X1 port map( A => n2, B => writeptr_1_port, Y => n86);
   U10 : BUFX2 port map( A => writeptr_0_port, Y => n2);
   U11 : INVX1 port map( A => writeptr_0_port, Y => n230);
   U12 : INVX4 port map( A => n338_port, Y => n3);
   U13 : INVX4 port map( A => n348, Y => n4);
   U14 : INVX1 port map( A => n542, Y => n5);
   U15 : INVX2 port map( A => n5, Y => n6);
   U16 : INVX1 port map( A => n573, Y => n7);
   U17 : INVX2 port map( A => n7, Y => n8);
   U18 : BUFX4 port map( A => n106, Y => n92);
   U19 : MUX2X1 port map( B => n170, A => opcode_6_0_port, S => n323, Y => n324
                           );
   U20 : INVX2 port map( A => n323, Y => n492);
   U21 : MUX2X1 port map( B => n170, A => opcode_2_0_port, S => n343_port, Y =>
                           n344_port);
   U22 : INVX2 port map( A => n29, Y => n555);
   U23 : INVX2 port map( A => n348, Y => n48);
   U24 : INVX2 port map( A => n338_port, Y => n47);
   U25 : AND2X2 port map( A => n1262, B => n120, Y => n9);
   U26 : AND2X1 port map( A => n1273, B => n120, Y => n10);
   U27 : AND2X2 port map( A => n1283, B => n120, Y => n11);
   U28 : AND2X2 port map( A => n1252, B => n1262, Y => n12);
   U29 : AND2X2 port map( A => n1282, B => n1252, Y => n13);
   U30 : AND2X1 port map( A => n1273, B => n1252, Y => n14);
   U31 : AND2X1 port map( A => n1253, B => n1252, Y => n15);
   U32 : AND2X2 port map( A => n1274, B => n1252, Y => n16);
   U33 : AND2X2 port map( A => n1283, B => n1252, Y => n17);
   U34 : AND2X1 port map( A => n1252, B => n1263, Y => n18);
   U35 : AND2X1 port map( A => n1253, B => n120, Y => n19);
   U36 : AND2X1 port map( A => n1274, B => n120, Y => n20);
   U37 : AND2X1 port map( A => n1263, B => n120, Y => n21);
   U38 : AND2X2 port map( A => n1282, B => n120, Y => n22);
   U39 : INVX1 port map( A => RCV_DATA(0), Y => n515);
   U40 : INVX1 port map( A => RCV_DATA(1), Y => n516);
   U41 : INVX1 port map( A => RCV_DATA(3), Y => n517);
   U42 : INVX1 port map( A => RCV_DATA(5), Y => n519);
   n23 <= '1';
   U44 : INVX1 port map( A => n553, Y => n554);
   U45 : INVX1 port map( A => RCV_DATA(4), Y => n518);
   U46 : INVX2 port map( A => n225, Y => n24);
   U47 : INVX2 port map( A => n225, Y => n394);
   U48 : INVX1 port map( A => n230, Y => n25);
   U49 : INVX1 port map( A => n547, Y => n26);
   U50 : INVX2 port map( A => n26, Y => n27);
   U51 : BUFX2 port map( A => n537, Y => n28);
   U52 : INVX1 port map( A => RCV_DATA(6), Y => n520);
   U53 : AND2X2 port map( A => n2, B => writeptr_1_port, Y => n29);
   U54 : INVX1 port map( A => RCV_DATA(7), Y => n521);
   U55 : INVX1 port map( A => n149, Y => n229);
   U56 : BUFX2 port map( A => n107, Y => n30);
   U57 : INVX2 port map( A => n272, Y => n31);
   U58 : INVX2 port map( A => n272, Y => n434);
   U59 : AND2X2 port map( A => n271, B => n308, Y => n32);
   U60 : INVX2 port map( A => n244, Y => n34);
   U61 : INVX2 port map( A => n244, Y => n404);
   U62 : NOR2X1 port map( A => n87, B => n85, Y => n35);
   U63 : INVX4 port map( A => n663, Y => n36);
   U64 : INVX1 port map( A => n82, Y => n37);
   U65 : XNOR2X1 port map( A => n547, B => n36, Y => n90);
   U66 : INVX1 port map( A => n566, Y => n38);
   U67 : INVX4 port map( A => n41, Y => n73);
   U68 : INVX2 port map( A => n333, Y => n39);
   U69 : INVX2 port map( A => n343_port, Y => n40);
   U70 : NAND2X1 port map( A => n271, B => n308, Y => n41);
   U71 : INVX2 port map( A => n264, Y => n42);
   U72 : INVX2 port map( A => n264, Y => n43);
   U73 : INVX2 port map( A => n264, Y => n433);
   U74 : INVX2 port map( A => n256, Y => n44);
   U75 : INVX2 port map( A => n256, Y => n430);
   U76 : INVX2 port map( A => n252, Y => n45);
   U77 : INVX2 port map( A => n252, Y => n46);
   U78 : INVX2 port map( A => n252, Y => n421);
   U79 : INVX1 port map( A => n574, Y => n49);
   U80 : INVX1 port map( A => writeptr_4_port, Y => n574);
   U81 : INVX2 port map( A => readptr_1_port, Y => n50);
   U82 : BUFX2 port map( A => n37, Y => n52);
   U83 : NAND2X1 port map( A => RCV_OPCODE(1), B => RCV_OPCODE(0), Y => n53);
   U84 : NAND2X1 port map( A => RCV_OPCODE(0), B => RCV_OPCODE(1), Y => n54);
   U85 : INVX2 port map( A => n243, Y => n55);
   U86 : INVX2 port map( A => n243, Y => n271);
   U87 : INVX2 port map( A => n260, Y => n56);
   U88 : INVX2 port map( A => n260, Y => n432);
   U89 : INVX2 port map( A => n323, Y => n57);
   U90 : INVX2 port map( A => n323, Y => n58);
   U91 : INVX1 port map( A => n235, Y => n59);
   U92 : INVX1 port map( A => n231, Y => n60);
   U93 : INVX1 port map( A => n221, Y => n61);
   U94 : INVX1 port map( A => n216, Y => n62);
   U95 : INVX1 port map( A => n211, Y => n63);
   U96 : INVX2 port map( A => n207, Y => n64);
   U97 : INVX2 port map( A => n207, Y => n365);
   U98 : INVX4 port map( A => n284, Y => n65);
   U99 : INVX2 port map( A => n284, Y => n451);
   U100 : INVX4 port map( A => n328, Y => n66);
   U101 : INVX2 port map( A => n328, Y => n501);
   U102 : INVX2 port map( A => n279, Y => n67);
   U103 : INVX2 port map( A => n279, Y => n442);
   U104 : AND2X2 port map( A => n239, B => n353, Y => n106);
   U105 : NAND2X1 port map( A => n578, B => n68, Y => n577);
   U106 : NOR2X1 port map( A => n565, B => n94, Y => n68);
   U107 : AND2X2 port map( A => n353, B => n354, Y => n69);
   U108 : AND2X2 port map( A => n353, B => n354, Y => n70);
   U109 : INVX2 port map( A => n333, Y => n71);
   U110 : INVX4 port map( A => n333, Y => n510);
   U111 : INVX4 port map( A => n343_port, Y => n513);
   U112 : INVX2 port map( A => n577, Y => n583);
   U113 : BUFX2 port map( A => n555, Y => n72);
   U114 : INVX2 port map( A => readptr_0_port, Y => n74);
   U115 : INVX2 port map( A => n74, Y => n75);
   U116 : INVX1 port map( A => n74, Y => n76);
   U117 : INVX4 port map( A => n51, Y => n594);
   U118 : AND2X2 port map( A => n51, B => n663, Y => n120);
   U119 : AND2X2 port map( A => n51, B => n36, Y => n121);
   U120 : INVX1 port map( A => n150, Y => n77);
   U121 : INVX2 port map( A => n569, Y => n78);
   U122 : INVX4 port map( A => n150, Y => n151);
   U123 : AND2X1 port map( A => n563, B => n562, Y => n564);
   U124 : INVX1 port map( A => n558, Y => n89);
   U125 : INVX4 port map( A => n278, Y => n472);
   U126 : INVX4 port map( A => n206, Y => n239);
   U127 : AND2X2 port map( A => n353, B => n354, Y => n79);
   U128 : AND2X2 port map( A => n353, B => n354, Y => n80);
   U129 : AND2X2 port map( A => R_ENABLE, B => n181, Y => n81);
   U130 : INVX2 port map( A => n81, Y => n597);
   U131 : BUFX2 port map( A => n230, Y => n82);
   U132 : INVX2 port map( A => n471, Y => n83);
   U133 : BUFX4 port map( A => readptr_4_port, Y => n84);
   U134 : AND2X2 port map( A => n524, B => n178, Y => n85);
   U135 : INVX1 port map( A => n85, Y => n522);
   U136 : XOR2X1 port map( A => n317, B => n88, Y => n87);
   U137 : INVX1 port map( A => n87, Y => n541);
   U138 : XNOR2X1 port map( A => n94, B => n153, Y => n88);
   U139 : INVX1 port map( A => n558, Y => n581);
   U140 : INVX1 port map( A => n90, Y => n540);
   U141 : INVX1 port map( A => n77, Y => n215);
   U142 : INVX8 port map( A => n148, Y => n149);
   U143 : NAND3X1 port map( A => n90, B => n35, C => n204, Y => n91);
   U144 : BUFX4 port map( A => n106, Y => n93);
   U145 : BUFX4 port map( A => writeptr_3_port, Y => n94);
   U146 : INVX2 port map( A => n21, Y => n131);
   U147 : INVX2 port map( A => n18, Y => n143);
   U148 : INVX2 port map( A => n14, Y => n144);
   U149 : INVX2 port map( A => n19, Y => n128);
   U150 : INVX2 port map( A => n20, Y => n133);
   U151 : AND2X1 port map( A => writeptr_4_port, B => n124, Y => n122);
   U152 : AND2X2 port map( A => n578, B => n353, Y => n95);
   U153 : INVX2 port map( A => n172, Y => n170);
   U154 : INVX2 port map( A => n176, Y => n174);
   U155 : INVX2 port map( A => n176, Y => n173);
   U156 : AND2X2 port map( A => n308, B => n578, Y => n96);
   U157 : AND2X2 port map( A => n472, B => n471, Y => n97);
   U158 : AND2X2 port map( A => n569, B => n578, Y => n98);
   U159 : AND2X2 port map( A => n471, B => n578, Y => n99);
   U160 : AND2X2 port map( A => n293, B => n578, Y => n100);
   U161 : AND2X2 port map( A => n283, B => n578, Y => n101);
   U162 : AND2X2 port map( A => n303, B => n578, Y => n102);
   U163 : INVX2 port map( A => RCV_OPCODE(0), Y => n172);
   U164 : INVX1 port map( A => RCV_OPCODE(1), Y => n176);
   U165 : AND2X2 port map( A => n277, B => W_ENABLE, Y => n103);
   U166 : AND2X2 port map( A => W_ENABLE, B => n91, Y => n104);
   U167 : AND2X2 port map( A => n288, B => n578, Y => n105);
   U168 : AND2X2 port map( A => n148, B => n2, Y => n107);
   U169 : INVX2 port map( A => RST, Y => n177);
   U170 : AND2X2 port map( A => n276, B => n574, Y => n108);
   U171 : AND2X2 port map( A => n1283, B => n121, Y => n109);
   U172 : AND2X2 port map( A => n1253, B => n121, Y => n110);
   U173 : AND2X2 port map( A => n1274, B => n121, Y => n111);
   U174 : AND2X2 port map( A => n1263, B => n121, Y => n112);
   U175 : AND2X2 port map( A => n1282, B => n121, Y => n113);
   U176 : AND2X2 port map( A => n1251, B => n121, Y => n114);
   U177 : AND2X2 port map( A => n1262, B => n121, Y => n115);
   U178 : AND2X2 port map( A => n1273, B => n121, Y => n116);
   U179 : XNOR2X1 port map( A => n573, B => n537, Y => n542);
   U180 : AND2X2 port map( A => n124, B => n574, Y => n117);
   U181 : INVX2 port map( A => n12, Y => n142);
   U182 : INVX4 port map( A => n13, Y => n146);
   U183 : INVX2 port map( A => n139, Y => n140);
   U184 : INVX1 port map( A => n838, Y => n139);
   U185 : INVX4 port map( A => n16, Y => n145);
   U186 : INVX4 port map( A => n17, Y => n147);
   U187 : INVX2 port map( A => n15, Y => n141);
   U188 : INVX4 port map( A => n22, Y => n136);
   U189 : INVX2 port map( A => n129, Y => n130);
   U190 : INVX1 port map( A => n839, Y => n129);
   U191 : INVX2 port map( A => n9, Y => n132);
   U192 : INVX2 port map( A => n10, Y => n134);
   U193 : INVX4 port map( A => n11, Y => n135);
   U194 : INVX2 port map( A => n119, Y => n137);
   U195 : INVX2 port map( A => n119, Y => n138);
   U196 : INVX2 port map( A => n155, Y => n154);
   U197 : INVX2 port map( A => n157, Y => n156);
   U198 : INVX2 port map( A => RCV_DATA(2), Y => n158);
   U199 : INVX2 port map( A => RCV_DATA(2), Y => n159);
   U200 : INVX2 port map( A => n161, Y => n160);
   U201 : INVX2 port map( A => n165, Y => n164);
   U202 : INVX2 port map( A => n163, Y => n162);
   U203 : INVX2 port map( A => n167, Y => n166);
   U204 : INVX2 port map( A => n169, Y => n168);
   U205 : AND2X2 port map( A => writeptr_4_port, B => n276, Y => n118);
   U206 : OR2X2 port map( A => n597, B => n182, Y => n119);
   U207 : XOR2X1 port map( A => n151, B => n51, Y => n123);
   U208 : INVX2 port map( A => writeptr_1_port, Y => n150);
   U209 : INVX2 port map( A => readptr_3_port, Y => n152);
   U210 : NOR2X1 port map( A => RST, B => n94, Y => n124);
   U211 : INVX2 port map( A => n517, Y => n161);
   U212 : INVX2 port map( A => n519, Y => n165);
   U213 : INVX2 port map( A => n515, Y => n155);
   U214 : INVX2 port map( A => n516, Y => n157);
   U215 : INVX2 port map( A => n518, Y => n163);
   U216 : INVX2 port map( A => n520, Y => n167);
   U217 : INVX2 port map( A => n521, Y => n169);
   U218 : BUFX2 port map( A => n352, Y => n125);
   U219 : BUFX4 port map( A => n352, Y => n126);
   U220 : INVX2 port map( A => writeptr_2_port, Y => n148);
   U221 : INVX1 port map( A => n337, Y => n471);
   U222 : INVX1 port map( A => n317, Y => n569);
   U223 : INVX1 port map( A => n172, Y => n171);
   U224 : INVX1 port map( A => n176, Y => n175);
   U225 : INVX4 port map( A => n318, Y => n127);
   U226 : INVX2 port map( A => n318, Y => n483);
   U227 : INVX4 port map( A => n563, Y => n578);
   U228 : INVX4 port map( A => n211, Y => n374);
   U229 : INVX4 port map( A => n216, Y => n383);
   U230 : INVX4 port map( A => n221, Y => n392);
   U231 : INVX4 port map( A => n231, Y => n395);
   U232 : INVX4 port map( A => n235, Y => n396);
   U233 : INVX4 port map( A => n289, Y => n460);
   U234 : INVX4 port map( A => n294, Y => n469);
   U235 : INVX4 port map( A => n304, Y => n473);
   U236 : INVX4 port map( A => n309, Y => n474);
   U237 : INVX4 port map( A => n313, Y => n475);
   U238 : AND2X2 port map( A => n1253, B => n1254, Y => n841);
   U239 : AND2X2 port map( A => n1251, B => n1254, Y => n840);
   U240 : AND2X2 port map( A => n1254, B => n1263, Y => n865);
   U241 : AND2X2 port map( A => n1254, B => n1262, Y => n852);
   U242 : AND2X2 port map( A => n1274, B => n1254, Y => n909);
   U243 : AND2X2 port map( A => n1273, B => n1254, Y => n908);
   U244 : AND2X2 port map( A => n1283, B => n1254, Y => n916);
   U245 : AND2X2 port map( A => n1282, B => n1254, Y => n915);
   U246 : INVX8 port map( A => n152, Y => n153);
   U247 : INVX2 port map( A => memory_16_7_port, Y => n780);
   U248 : INVX2 port map( A => memory_17_7_port, Y => n788);
   U249 : INVX2 port map( A => memory_18_7_port, Y => n796);
   U250 : INVX2 port map( A => readptr_2_port, Y => n663);
   U251 : INVX2 port map( A => memory_19_7_port, Y => n804);
   U252 : NAND2X1 port map( A => n1251, B => n120, Y => n839);
   U253 : INVX2 port map( A => memory_24_7_port, Y => n706);
   U254 : INVX2 port map( A => memory_25_7_port, Y => n698);
   U255 : INVX2 port map( A => memory_26_7_port, Y => n690);
   U256 : INVX2 port map( A => memory_27_7_port, Y => n682);
   U257 : INVX2 port map( A => memory_3_7_port, Y => n745);
   U258 : INVX2 port map( A => memory_2_7_port, Y => n737);
   U259 : INVX2 port map( A => memory_1_7_port, Y => n729);
   U260 : INVX2 port map( A => memory_0_7_port, Y => n721);
   U261 : INVX2 port map( A => memory_8_7_port, Y => n748);
   U262 : INVX2 port map( A => memory_9_7_port, Y => n756);
   U263 : INVX2 port map( A => memory_10_7_port, Y => n764);
   U264 : INVX2 port map( A => memory_11_7_port, Y => n772);
   U265 : INVX2 port map( A => memory_16_6_port, Y => n781);
   U266 : INVX2 port map( A => memory_17_6_port, Y => n789);
   U267 : INVX2 port map( A => memory_18_6_port, Y => n797);
   U268 : INVX2 port map( A => memory_19_6_port, Y => n805);
   U269 : INVX2 port map( A => memory_24_6_port, Y => n707);
   U270 : INVX2 port map( A => memory_25_6_port, Y => n699);
   U271 : INVX2 port map( A => memory_26_6_port, Y => n691);
   U272 : INVX2 port map( A => memory_27_6_port, Y => n683);
   U273 : INVX2 port map( A => memory_3_6_port, Y => n744);
   U274 : INVX2 port map( A => memory_2_6_port, Y => n736);
   U275 : INVX2 port map( A => memory_1_6_port, Y => n728);
   U276 : INVX2 port map( A => memory_0_6_port, Y => n720);
   U277 : INVX2 port map( A => memory_8_6_port, Y => n749);
   U278 : INVX2 port map( A => memory_9_6_port, Y => n757);
   U279 : INVX2 port map( A => memory_10_6_port, Y => n765);
   U280 : INVX2 port map( A => memory_11_6_port, Y => n773);
   U281 : INVX2 port map( A => memory_16_5_port, Y => n782);
   U282 : INVX2 port map( A => memory_17_5_port, Y => n790);
   U283 : INVX2 port map( A => memory_18_5_port, Y => n798);
   U284 : INVX2 port map( A => memory_19_5_port, Y => n806);
   U285 : INVX2 port map( A => memory_24_5_port, Y => n708);
   U286 : INVX2 port map( A => memory_25_5_port, Y => n700);
   U287 : INVX2 port map( A => memory_26_5_port, Y => n692);
   U288 : INVX2 port map( A => memory_27_5_port, Y => n684);
   U289 : INVX2 port map( A => memory_3_5_port, Y => n743);
   U290 : INVX2 port map( A => memory_2_5_port, Y => n735);
   U291 : INVX2 port map( A => memory_1_5_port, Y => n727);
   U292 : INVX2 port map( A => memory_0_5_port, Y => n719);
   U293 : INVX2 port map( A => memory_8_5_port, Y => n750);
   U294 : INVX2 port map( A => memory_9_5_port, Y => n758);
   U295 : INVX2 port map( A => memory_10_5_port, Y => n766);
   U296 : INVX2 port map( A => memory_11_5_port, Y => n774);
   U297 : INVX2 port map( A => memory_16_4_port, Y => n783);
   U298 : INVX2 port map( A => memory_17_4_port, Y => n791);
   U299 : INVX2 port map( A => memory_18_4_port, Y => n799);
   U300 : INVX2 port map( A => memory_19_4_port, Y => n807);
   U301 : INVX2 port map( A => memory_24_4_port, Y => n709);
   U302 : INVX2 port map( A => memory_25_4_port, Y => n701);
   U303 : INVX2 port map( A => memory_26_4_port, Y => n693);
   U304 : INVX2 port map( A => memory_27_4_port, Y => n685);
   U305 : INVX2 port map( A => memory_3_4_port, Y => n742);
   U306 : INVX2 port map( A => memory_2_4_port, Y => n734);
   U307 : INVX2 port map( A => memory_1_4_port, Y => n726);
   U308 : INVX2 port map( A => memory_0_4_port, Y => n718);
   U309 : INVX2 port map( A => memory_8_4_port, Y => n751);
   U310 : INVX2 port map( A => memory_9_4_port, Y => n759);
   U311 : INVX2 port map( A => memory_10_4_port, Y => n767);
   U312 : INVX2 port map( A => memory_11_4_port, Y => n775);
   U313 : INVX2 port map( A => memory_16_3_port, Y => n784);
   U314 : INVX2 port map( A => memory_17_3_port, Y => n792);
   U315 : INVX2 port map( A => memory_18_3_port, Y => n800);
   U316 : INVX2 port map( A => memory_19_3_port, Y => n808);
   U317 : INVX2 port map( A => memory_24_3_port, Y => n710);
   U318 : INVX2 port map( A => memory_25_3_port, Y => n702);
   U319 : INVX2 port map( A => memory_26_3_port, Y => n694);
   U320 : INVX2 port map( A => memory_27_3_port, Y => n686);
   U321 : INVX2 port map( A => memory_3_3_port, Y => n741);
   U322 : INVX2 port map( A => memory_2_3_port, Y => n733);
   U323 : INVX2 port map( A => memory_1_3_port, Y => n725);
   U324 : INVX2 port map( A => memory_0_3_port, Y => n717);
   U325 : INVX2 port map( A => memory_8_3_port, Y => n752);
   U326 : INVX2 port map( A => memory_9_3_port, Y => n760);
   U327 : INVX2 port map( A => memory_10_3_port, Y => n768);
   U328 : INVX2 port map( A => memory_11_3_port, Y => n776);
   U329 : INVX2 port map( A => memory_16_2_port, Y => n785);
   U330 : INVX2 port map( A => memory_17_2_port, Y => n793);
   U331 : INVX2 port map( A => memory_18_2_port, Y => n801);
   U332 : INVX2 port map( A => memory_19_2_port, Y => n809);
   U333 : INVX2 port map( A => memory_24_2_port, Y => n711);
   U334 : INVX2 port map( A => memory_25_2_port, Y => n703);
   U335 : INVX2 port map( A => memory_26_2_port, Y => n695);
   U336 : INVX2 port map( A => memory_27_2_port, Y => n687);
   U337 : INVX2 port map( A => memory_3_2_port, Y => n740);
   U338 : INVX2 port map( A => memory_2_2_port, Y => n732);
   U339 : INVX2 port map( A => memory_1_2_port, Y => n724);
   U340 : INVX2 port map( A => memory_0_2_port, Y => n716);
   U341 : INVX2 port map( A => memory_8_2_port, Y => n753);
   U342 : INVX2 port map( A => memory_9_2_port, Y => n761);
   U343 : INVX2 port map( A => memory_10_2_port, Y => n769);
   U344 : INVX2 port map( A => memory_11_2_port, Y => n777);
   U345 : INVX2 port map( A => memory_16_1_port, Y => n786);
   U346 : INVX2 port map( A => memory_17_1_port, Y => n794);
   U347 : INVX2 port map( A => memory_18_1_port, Y => n802);
   U348 : INVX2 port map( A => memory_19_1_port, Y => n810);
   U349 : INVX2 port map( A => memory_24_1_port, Y => n712);
   U350 : INVX2 port map( A => memory_25_1_port, Y => n704);
   U351 : INVX2 port map( A => memory_26_1_port, Y => n696);
   U352 : INVX2 port map( A => memory_27_1_port, Y => n688);
   U353 : INVX2 port map( A => memory_3_1_port, Y => n739);
   U354 : INVX2 port map( A => memory_2_1_port, Y => n731);
   U355 : INVX2 port map( A => memory_1_1_port, Y => n723);
   U356 : INVX2 port map( A => memory_0_1_port, Y => n715);
   U357 : INVX2 port map( A => memory_8_1_port, Y => n754);
   U358 : INVX2 port map( A => memory_9_1_port, Y => n762);
   U359 : INVX2 port map( A => memory_10_1_port, Y => n770);
   U360 : INVX2 port map( A => memory_11_1_port, Y => n778);
   U361 : INVX2 port map( A => memory_16_0_port, Y => n787);
   U362 : INVX2 port map( A => memory_17_0_port, Y => n795);
   U363 : INVX2 port map( A => memory_18_0_port, Y => n803);
   U364 : INVX2 port map( A => memory_19_0_port, Y => n811);
   U365 : INVX2 port map( A => memory_24_0_port, Y => n713);
   U366 : INVX2 port map( A => memory_25_0_port, Y => n705);
   U367 : INVX2 port map( A => memory_26_0_port, Y => n697);
   U368 : INVX2 port map( A => memory_27_0_port, Y => n689);
   U369 : INVX2 port map( A => memory_3_0_port, Y => n738);
   U370 : INVX2 port map( A => memory_2_0_port, Y => n730);
   U371 : INVX2 port map( A => memory_1_0_port, Y => n722);
   U372 : INVX2 port map( A => memory_0_0_port, Y => n714);
   U373 : INVX2 port map( A => memory_8_0_port, Y => n755);
   U374 : INVX2 port map( A => memory_9_0_port, Y => n763);
   U375 : INVX2 port map( A => memory_10_0_port, Y => n771);
   U376 : INVX2 port map( A => memory_11_0_port, Y => n779);
   U377 : INVX2 port map( A => opcode_16_1_port, Y => n820);
   U378 : INVX2 port map( A => opcode_17_1_port, Y => n822);
   U379 : INVX2 port map( A => opcode_18_1_port, Y => n824);
   U380 : INVX2 port map( A => opcode_19_1_port, Y => n826);
   U381 : INVX2 port map( A => opcode_24_1_port, Y => n672);
   U382 : INVX2 port map( A => opcode_25_1_port, Y => n670);
   U383 : INVX2 port map( A => opcode_26_1_port, Y => n668);
   U384 : INVX2 port map( A => opcode_27_1_port, Y => n666);
   U385 : INVX2 port map( A => opcode_3_1_port, Y => n681);
   U386 : INVX2 port map( A => opcode_2_1_port, Y => n679);
   U387 : INVX2 port map( A => opcode_1_1_port, Y => n677);
   U388 : INVX2 port map( A => opcode_0_1_port, Y => n675);
   U389 : INVX2 port map( A => opcode_8_1_port, Y => n812);
   U390 : INVX2 port map( A => opcode_9_1_port, Y => n814);
   U391 : INVX2 port map( A => opcode_10_1_port, Y => n816);
   U392 : INVX2 port map( A => opcode_11_1_port, Y => n818);
   U393 : INVX2 port map( A => opcode_16_0_port, Y => n821);
   U394 : INVX2 port map( A => opcode_17_0_port, Y => n823);
   U395 : INVX2 port map( A => opcode_18_0_port, Y => n825);
   U396 : INVX2 port map( A => opcode_19_0_port, Y => n827);
   U397 : INVX2 port map( A => n75, Y => n662);
   U398 : INVX2 port map( A => n153, Y => n664);
   U399 : INVX2 port map( A => opcode_24_0_port, Y => n673);
   U400 : INVX2 port map( A => opcode_25_0_port, Y => n671);
   U401 : INVX2 port map( A => opcode_26_0_port, Y => n669);
   U402 : INVX2 port map( A => opcode_27_0_port, Y => n667);
   U403 : INVX2 port map( A => opcode_3_0_port, Y => n680);
   U404 : INVX2 port map( A => opcode_2_0_port, Y => n678);
   U405 : INVX2 port map( A => opcode_1_0_port, Y => n676);
   U406 : INVX2 port map( A => opcode_0_0_port, Y => n674);
   U407 : INVX2 port map( A => n84, Y => n665);
   U408 : INVX2 port map( A => opcode_8_0_port, Y => n813);
   U409 : INVX2 port map( A => opcode_9_0_port, Y => n815);
   U410 : INVX2 port map( A => opcode_10_0_port, Y => n817);
   U411 : INVX2 port map( A => opcode_11_0_port, Y => n819);
   U412 : NAND2X1 port map( A => n75, B => n82, Y => n524);
   U413 : NAND2X1 port map( A => n37, B => n662, Y => n178);
   U414 : NOR2X1 port map( A => n123, B => n522, Y => n180);
   U415 : XNOR2X1 port map( A => n149, B => n36, Y => n527);
   U416 : XNOR2X1 port map( A => n94, B => n153, Y => n532);
   U417 : XNOR2X1 port map( A => writeptr_4_port, B => n84, Y => n537);
   U418 : AND2X2 port map( A => n532, B => n537, Y => n179);
   U419 : NAND3X1 port map( A => n180, B => n527, C => n179, Y => n181);
   U420 : MUX2X1 port map( B => n181, A => n747, S => RST, Y => n1415);
   U421 : INVX2 port map( A => OUT_OPCODE_0_port, Y => n184);
   U422 : INVX2 port map( A => n1241, Y => n183);
   U423 : NAND2X1 port map( A => n177, B => state, Y => n182);
   U424 : MUX2X1 port map( B => n184, A => n183, S => n137, Y => n1030);
   U425 : INVX2 port map( A => OUT_OPCODE_1_port, Y => n186);
   U426 : INVX2 port map( A => n1214, Y => n185);
   U427 : MUX2X1 port map( B => n186, A => n185, S => n138, Y => n1031);
   U428 : INVX2 port map( A => DATA_0_port, Y => n188);
   U429 : INVX2 port map( A => n1187, Y => n187);
   U430 : MUX2X1 port map( B => n188, A => n187, S => n137, Y => n1032);
   U431 : INVX2 port map( A => DATA_1_port, Y => n190);
   U432 : INVX2 port map( A => n1064, Y => n189);
   U433 : MUX2X1 port map( B => n190, A => n189, S => n138, Y => n1033);
   U434 : INVX2 port map( A => DATA_2_port, Y => n192);
   U435 : INVX2 port map( A => n1025, Y => n191);
   U436 : MUX2X1 port map( B => n192, A => n191, S => n137, Y => n1034);
   U437 : INVX2 port map( A => DATA_3_port, Y => n194);
   U438 : INVX2 port map( A => n998, Y => n193);
   U439 : MUX2X1 port map( B => n194, A => n193, S => n138, Y => n1035);
   U440 : INVX2 port map( A => DATA_4_port, Y => n196);
   U441 : INVX2 port map( A => n971, Y => n195);
   U442 : MUX2X1 port map( B => n196, A => n195, S => n137, Y => n1036);
   U443 : INVX2 port map( A => DATA_5_port, Y => n198);
   U444 : INVX2 port map( A => n944, Y => n197);
   U445 : MUX2X1 port map( B => n198, A => n197, S => n138, Y => n1037);
   U446 : INVX2 port map( A => DATA_6_port, Y => n200);
   U447 : INVX2 port map( A => n917, Y => n199);
   U448 : MUX2X1 port map( B => n200, A => n199, S => n137, Y => n1038);
   U449 : INVX2 port map( A => DATA_7_port, Y => n202);
   U450 : INVX2 port map( A => n828, Y => n201);
   U451 : MUX2X1 port map( B => n202, A => n201, S => n138, Y => n1039);
   U452 : NAND2X1 port map( A => n30, B => n215, Y => n347_port);
   U453 : INVX2 port map( A => n347_port, Y => n308);
   U454 : INVX2 port map( A => n54, Y => n566);
   U455 : NAND2X1 port map( A => n107, B => n151, Y => n337);
   U456 : NAND2X1 port map( A => n555, B => n149, Y => n203);
   U457 : NAND2X1 port map( A => n337, B => n203, Y => n547);
   U458 : NAND2X1 port map( A => n149, B => n29, Y => n317);
   U459 : NOR2X1 port map( A => n87, B => n85, Y => n205);
   U460 : XNOR2X1 port map( A => n151, B => n25, Y => n553);
   U461 : XNOR2X1 port map( A => n553, B => n594, Y => n544);
   U462 : NAND3X1 port map( A => n94, B => n86, C => n149, Y => n573);
   U463 : AND2X2 port map( A => n544, B => n542, Y => n204);
   U464 : NAND3X1 port map( A => n90, B => n205, C => n204, Y => n277);
   U465 : NAND2X1 port map( A => W_ENABLE, B => n277, Y => n558);
   U466 : NAND2X1 port map( A => n566, B => n581, Y => n563);
   U467 : NAND2X1 port map( A => n96, B => n117, Y => n210);
   U468 : NAND2X1 port map( A => n94, B => n177, Y => n298);
   U469 : INVX2 port map( A => n298, Y => n276);
   U470 : NAND3X1 port map( A => n118, B => n103, C => n53, Y => n206);
   U471 : NAND2X1 port map( A => n239, B => n569, Y => n207);
   U472 : MUX2X1 port map( B => opcode_31_0_port, A => n171, S => n365, Y => 
                           n208);
   U473 : NAND2X1 port map( A => n210, B => n208, Y => n605);
   U474 : MUX2X1 port map( B => opcode_31_1_port, A => n175, S => n365, Y => 
                           n209);
   U475 : NAND2X1 port map( A => n210, B => n209, Y => n604);
   U476 : OR2X2 port map( A => n77, B => n52, Y => n556);
   U477 : INVX2 port map( A => n556, Y => n220);
   U478 : NAND2X1 port map( A => n220, B => n229, Y => n565);
   U479 : INVX2 port map( A => n565, Y => n353);
   U480 : NAND2X1 port map( A => n117, B => n95, Y => n214);
   U481 : NAND3X1 port map( A => n149, B => n77, C => n82, Y => n322);
   U482 : INVX2 port map( A => n322, Y => n283);
   U483 : NAND2X1 port map( A => n239, B => n283, Y => n211);
   U484 : MUX2X1 port map( B => opcode_30_0_port, A => n171, S => n374, Y => 
                           n212);
   U485 : NAND2X1 port map( A => n214, B => n212, Y => n617);
   U486 : MUX2X1 port map( B => opcode_30_1_port, A => n175, S => n374, Y => 
                           n213);
   U487 : NAND2X1 port map( A => n214, B => n213, Y => n616);
   U488 : NAND2X1 port map( A => n98, B => n118, Y => n219);
   U489 : NAND3X1 port map( A => n149, B => n52, C => n215, Y => n327);
   U490 : INVX2 port map( A => n327, Y => n288);
   U491 : NAND2X1 port map( A => n239, B => n288, Y => n216);
   U492 : MUX2X1 port map( B => opcode_29_0_port, A => n171, S => n383, Y => 
                           n217);
   U493 : NAND2X1 port map( A => n219, B => n217, Y => n633);
   U494 : MUX2X1 port map( B => opcode_29_1_port, A => n175, S => n383, Y => 
                           n218);
   U495 : NAND2X1 port map( A => n219, B => n218, Y => n632);
   U496 : NAND2X1 port map( A => n101, B => n118, Y => n224);
   U497 : NAND2X1 port map( A => n220, B => n149, Y => n332);
   U498 : INVX2 port map( A => n332, Y => n293);
   U499 : NAND2X1 port map( A => n239, B => n293, Y => n221);
   U500 : MUX2X1 port map( B => opcode_28_0_port, A => n171, S => n392, Y => 
                           n222);
   U501 : NAND2X1 port map( A => n224, B => n222, Y => n645);
   U502 : MUX2X1 port map( B => opcode_28_1_port, A => n175, S => n392, Y => 
                           n223);
   U503 : NAND2X1 port map( A => n224, B => n223, Y => n644);
   U504 : NAND2X1 port map( A => n105, B => n118, Y => n228);
   U505 : NAND2X1 port map( A => n239, B => n471, Y => n225);
   U506 : MUX2X1 port map( B => opcode_27_0_port, A => n171, S => n394, Y => 
                           n226);
   U507 : NAND2X1 port map( A => n228, B => n226, Y => n651);
   U508 : MUX2X1 port map( B => opcode_27_1_port, A => n175, S => n394, Y => 
                           n227);
   U509 : NAND2X1 port map( A => n228, B => n227, Y => n650);
   U510 : NAND2X1 port map( A => n100, B => n118, Y => n234);
   U511 : NAND3X1 port map( A => n77, B => n82, C => n229, Y => n342_port);
   U512 : INVX2 port map( A => n342_port, Y => n303);
   U513 : NAND2X1 port map( A => n239, B => n303, Y => n231);
   U514 : MUX2X1 port map( B => opcode_26_0_port, A => n171, S => n395, Y => 
                           n232);
   U515 : NAND2X1 port map( A => n234, B => n232, Y => n631);
   U516 : MUX2X1 port map( B => opcode_26_1_port, A => n175, S => n395, Y => 
                           n233);
   U517 : NAND2X1 port map( A => n234, B => n233, Y => n630);
   U518 : NAND2X1 port map( A => n99, B => n118, Y => n238);
   U519 : NAND2X1 port map( A => n239, B => n308, Y => n235);
   U520 : MUX2X1 port map( B => opcode_25_0_port, A => n171, S => n396, Y => 
                           n236);
   U521 : NAND2X1 port map( A => n238, B => n236, Y => n657);
   U522 : MUX2X1 port map( B => opcode_25_1_port, A => n175, S => n396, Y => 
                           n237);
   U523 : NAND2X1 port map( A => n238, B => n237, Y => n656);
   U524 : NAND2X1 port map( A => n102, B => n118, Y => n242);
   U525 : MUX2X1 port map( B => opcode_24_0_port, A => n170, S => n92, Y => 
                           n240);
   U526 : NAND2X1 port map( A => n242, B => n240, Y => n607);
   U527 : MUX2X1 port map( B => opcode_24_1_port, A => n174, S => n92, Y => 
                           n241);
   U528 : NAND2X1 port map( A => n242, B => n241, Y => n606);
   U529 : NAND2X1 port map( A => n96, B => n118, Y => n247);
   U530 : NAND3X1 port map( A => n122, B => n53, C => n103, Y => n243);
   U531 : NAND2X1 port map( A => n55, B => n569, Y => n244);
   U532 : MUX2X1 port map( B => opcode_23_0_port, A => n170, S => n404, Y => 
                           n245);
   U533 : NAND2X1 port map( A => n247, B => n245, Y => n619);
   U534 : MUX2X1 port map( B => opcode_23_1_port, A => n174, S => n404, Y => 
                           n246);
   U535 : NAND2X1 port map( A => n247, B => n246, Y => n618);
   U536 : NAND2X1 port map( A => n118, B => n95, Y => n251);
   U537 : NAND2X1 port map( A => n55, B => n283, Y => n248);
   U538 : MUX2X1 port map( B => opcode_22_0_port, A => n170, S => n1, Y => n249
                           );
   U539 : NAND2X1 port map( A => n251, B => n249, Y => n621);
   U540 : MUX2X1 port map( B => opcode_22_1_port, A => n174, S => n1, Y => n250
                           );
   U541 : NAND2X1 port map( A => n251, B => n250, Y => n620);
   U542 : NAND2X1 port map( A => n98, B => n122, Y => n255);
   U543 : NAND2X1 port map( A => n271, B => n288, Y => n252);
   U544 : MUX2X1 port map( B => opcode_21_0_port, A => n170, S => n421, Y => 
                           n253);
   U545 : NAND2X1 port map( A => n255, B => n253, Y => n661);
   U546 : MUX2X1 port map( B => opcode_21_1_port, A => n174, S => n421, Y => 
                           n254);
   U547 : NAND2X1 port map( A => n255, B => n254, Y => n660);
   U548 : NAND2X1 port map( A => n101, B => n122, Y => n259);
   U549 : NAND2X1 port map( A => n271, B => n293, Y => n256);
   U550 : MUX2X1 port map( B => opcode_20_0_port, A => n170, S => n430, Y => 
                           n257);
   U551 : NAND2X1 port map( A => n259, B => n257, Y => n659);
   U552 : MUX2X1 port map( B => opcode_20_1_port, A => n174, S => n430, Y => 
                           n258);
   U553 : NAND2X1 port map( A => n259, B => n258, Y => n658);
   U554 : NAND2X1 port map( A => n105, B => n122, Y => n263);
   U555 : NAND2X1 port map( A => n55, B => n471, Y => n260);
   U556 : MUX2X1 port map( B => opcode_19_0_port, A => n170, S => n432, Y => 
                           n261);
   U557 : NAND2X1 port map( A => n263, B => n261, Y => n629);
   U558 : MUX2X1 port map( B => opcode_19_1_port, A => n174, S => n432, Y => 
                           n262);
   U559 : NAND2X1 port map( A => n263, B => n262, Y => n628);
   U560 : NAND2X1 port map( A => n100, B => n122, Y => n267);
   U561 : NAND2X1 port map( A => n271, B => n303, Y => n264);
   U562 : MUX2X1 port map( B => opcode_18_0_port, A => n170, S => n433, Y => 
                           n265);
   U563 : NAND2X1 port map( A => n267, B => n265, Y => n603);
   U564 : MUX2X1 port map( B => opcode_18_1_port, A => n174, S => n433, Y => 
                           n266);
   U565 : NAND2X1 port map( A => n267, B => n266, Y => n602);
   U566 : NAND2X1 port map( A => n99, B => n122, Y => n270);
   U567 : MUX2X1 port map( B => opcode_17_0_port, A => n170, S => n73, Y => 
                           n268);
   U568 : NAND2X1 port map( A => n270, B => n268, Y => n613);
   U569 : MUX2X1 port map( B => opcode_17_1_port, A => n174, S => n73, Y => 
                           n269);
   U570 : NAND2X1 port map( A => n270, B => n269, Y => n612);
   U571 : NAND2X1 port map( A => n102, B => n122, Y => n275);
   U572 : NAND2X1 port map( A => n353, B => n55, Y => n272);
   U573 : MUX2X1 port map( B => opcode_16_0_port, A => n170, S => n434, Y => 
                           n273);
   U574 : NAND2X1 port map( A => n275, B => n273, Y => n627);
   U575 : MUX2X1 port map( B => opcode_16_1_port, A => n174, S => n434, Y => 
                           n274);
   U576 : NAND2X1 port map( A => n275, B => n274, Y => n626);
   U577 : NAND2X1 port map( A => n96, B => n122, Y => n282);
   U578 : NAND3X1 port map( A => n108, B => n104, C => n54, Y => n278);
   U579 : NAND2X1 port map( A => n472, B => n569, Y => n279);
   U580 : MUX2X1 port map( B => opcode_15_0_port, A => n170, S => n442, Y => 
                           n280);
   U581 : NAND2X1 port map( A => n282, B => n280, Y => n649);
   U582 : MUX2X1 port map( B => opcode_15_1_port, A => n174, S => n442, Y => 
                           n281);
   U583 : NAND2X1 port map( A => n282, B => n281, Y => n648);
   U584 : NAND2X1 port map( A => n122, B => n95, Y => n287);
   U585 : NAND2X1 port map( A => n472, B => n283, Y => n284);
   U586 : MUX2X1 port map( B => opcode_14_0_port, A => n170, S => n451, Y => 
                           n285);
   U587 : NAND2X1 port map( A => n287, B => n285, Y => n637);
   U588 : MUX2X1 port map( B => opcode_14_1_port, A => n174, S => n451, Y => 
                           n286);
   U589 : NAND2X1 port map( A => n287, B => n286, Y => n636);
   U590 : NAND2X1 port map( A => n98, B => n108, Y => n292);
   U591 : NAND2X1 port map( A => n472, B => n288, Y => n289);
   U592 : MUX2X1 port map( B => opcode_13_0_port, A => n170, S => n460, Y => 
                           n290);
   U593 : NAND2X1 port map( A => n292, B => n290, Y => n639);
   U594 : MUX2X1 port map( B => opcode_13_1_port, A => n174, S => n460, Y => 
                           n291);
   U595 : NAND2X1 port map( A => n292, B => n291, Y => n638);
   U596 : NAND2X1 port map( A => n101, B => n108, Y => n297);
   U597 : NAND2X1 port map( A => n472, B => n293, Y => n294);
   U598 : MUX2X1 port map( B => opcode_12_0_port, A => n171, S => n469, Y => 
                           n295);
   U599 : NAND2X1 port map( A => n297, B => n295, Y => n643);
   U600 : MUX2X1 port map( B => opcode_12_1_port, A => n173, S => n469, Y => 
                           n296);
   U601 : NAND2X1 port map( A => n297, B => n296, Y => n642);
   U602 : MUX2X1 port map( B => n83, A => n327, S => n566, Y => n300);
   U603 : NOR2X1 port map( A => n558, B => n298, Y => n299);
   U604 : NAND3X1 port map( A => n300, B => n574, C => n299, Y => n301);
   U605 : INVX2 port map( A => n301, Y => n302);
   U606 : MUX2X1 port map( B => n819, A => n172, S => n302, Y => n1056);
   U607 : MUX2X1 port map( B => n818, A => n176, S => n302, Y => n1057);
   U608 : NAND2X1 port map( A => n100, B => n108, Y => n307);
   U609 : NAND2X1 port map( A => n472, B => n303, Y => n304);
   U610 : MUX2X1 port map( B => opcode_10_0_port, A => n170, S => n473, Y => 
                           n305);
   U611 : NAND2X1 port map( A => n307, B => n305, Y => n647);
   U612 : MUX2X1 port map( B => opcode_10_1_port, A => n173, S => n473, Y => 
                           n306);
   U613 : NAND2X1 port map( A => n307, B => n306, Y => n646);
   U614 : NAND2X1 port map( A => n99, B => n108, Y => n312);
   U615 : NAND2X1 port map( A => n472, B => n308, Y => n309);
   U616 : MUX2X1 port map( B => opcode_9_0_port, A => n170, S => n474, Y => 
                           n310);
   U617 : NAND2X1 port map( A => n312, B => n310, Y => n623);
   U618 : MUX2X1 port map( B => opcode_9_1_port, A => n173, S => n474, Y => 
                           n311);
   U619 : NAND2X1 port map( A => n312, B => n311, Y => n622);
   U620 : NAND2X1 port map( A => n102, B => n108, Y => n316);
   U621 : NAND2X1 port map( A => n472, B => n353, Y => n313);
   U622 : MUX2X1 port map( B => opcode_8_0_port, A => n170, S => n475, Y => 
                           n314);
   U623 : NAND2X1 port map( A => n316, B => n314, Y => n635);
   U624 : MUX2X1 port map( B => opcode_8_1_port, A => n173, S => n475, Y => 
                           n315);
   U625 : NAND2X1 port map( A => n316, B => n315, Y => n634);
   U626 : NAND2X1 port map( A => n96, B => n108, Y => n321);
   U627 : NAND3X1 port map( A => n53, B => n117, C => n104, Y => n352);
   U628 : OR2X2 port map( A => n126, B => n78, Y => n318);
   U629 : MUX2X1 port map( B => opcode_7_0_port, A => n170, S => n483, Y => 
                           n319);
   U630 : NAND2X1 port map( A => n321, B => n319, Y => n609);
   U631 : MUX2X1 port map( B => opcode_7_1_port, A => n173, S => n483, Y => 
                           n320);
   U632 : NAND2X1 port map( A => n321, B => n320, Y => n608);
   U633 : NAND2X1 port map( A => n108, B => n95, Y => n326);
   U634 : OR2X2 port map( A => n125, B => n322, Y => n323);
   U635 : NAND2X1 port map( A => n326, B => n324, Y => n601);
   U636 : MUX2X1 port map( B => opcode_6_1_port, A => n173, S => n492, Y => 
                           n325);
   U637 : NAND2X1 port map( A => n326, B => n325, Y => n600);
   U638 : NAND2X1 port map( A => n98, B => n117, Y => n331);
   U639 : OR2X2 port map( A => n125, B => n327, Y => n328);
   U640 : MUX2X1 port map( B => opcode_5_0_port, A => n170, S => n501, Y => 
                           n329);
   U641 : NAND2X1 port map( A => n331, B => n329, Y => n615);
   U642 : MUX2X1 port map( B => opcode_5_1_port, A => n173, S => n501, Y => 
                           n330);
   U643 : NAND2X1 port map( A => n331, B => n330, Y => n614);
   U644 : NAND2X1 port map( A => n101, B => n117, Y => n336);
   U645 : OR2X2 port map( A => n126, B => n332, Y => n333);
   U646 : MUX2X1 port map( B => opcode_4_0_port, A => n171, S => n510, Y => 
                           n334);
   U647 : NAND2X1 port map( A => n336, B => n334, Y => n641);
   U648 : MUX2X1 port map( B => opcode_4_1_port, A => n173, S => n510, Y => 
                           n335);
   U649 : NAND2X1 port map( A => n336, B => n335, Y => n640);
   U650 : NAND2X1 port map( A => n105, B => n117, Y => n341_port);
   U651 : OR2X2 port map( A => n126, B => n83, Y => n338_port);
   U652 : MUX2X1 port map( B => opcode_3_0_port, A => n170, S => n512, Y => 
                           n339_port);
   U653 : NAND2X1 port map( A => n341_port, B => n339_port, Y => n625);
   U654 : MUX2X1 port map( B => opcode_3_1_port, A => n173, S => n512, Y => 
                           n340_port);
   U655 : NAND2X1 port map( A => n341_port, B => n340_port, Y => n624);
   U656 : NAND2X1 port map( A => n100, B => n117, Y => n346_port);
   U657 : OR2X2 port map( A => n126, B => n342_port, Y => n343_port);
   U658 : NAND2X1 port map( A => n346_port, B => n344_port, Y => n655);
   U659 : MUX2X1 port map( B => opcode_2_1_port, A => n173, S => n513, Y => 
                           n345_port);
   U660 : NAND2X1 port map( A => n346_port, B => n345_port, Y => n654);
   U661 : NAND2X1 port map( A => n99, B => n117, Y => n351);
   U662 : OR2X2 port map( A => n126, B => n347_port, Y => n348);
   U663 : MUX2X1 port map( B => opcode_1_0_port, A => n170, S => n514, Y => 
                           n349);
   U664 : NAND2X1 port map( A => n351, B => n349, Y => n653);
   U665 : MUX2X1 port map( B => opcode_1_1_port, A => n173, S => n514, Y => 
                           n350);
   U666 : NAND2X1 port map( A => n351, B => n350, Y => n652);
   U667 : NAND2X1 port map( A => n102, B => n117, Y => n357);
   U668 : INVX2 port map( A => n125, Y => n354);
   U669 : MUX2X1 port map( B => opcode_0_0_port, A => n170, S => n69, Y => n355
                           );
   U670 : NAND2X1 port map( A => n357, B => n355, Y => n611);
   U671 : MUX2X1 port map( B => opcode_0_1_port, A => n173, S => n69, Y => n356
                           );
   U672 : NAND2X1 port map( A => n357, B => n356, Y => n610);
   U673 : INVX2 port map( A => memory_31_0_port, Y => n358);
   U674 : MUX2X1 port map( B => n358, A => n154, S => n64, Y => n1072);
   U675 : INVX2 port map( A => memory_31_1_port, Y => n359);
   U676 : MUX2X1 port map( B => n359, A => n156, S => n64, Y => n1073);
   U677 : INVX2 port map( A => memory_31_2_port, Y => n360);
   U678 : MUX2X1 port map( B => n360, A => n158, S => n64, Y => n1074);
   U679 : INVX2 port map( A => memory_31_3_port, Y => n361);
   U680 : MUX2X1 port map( B => n361, A => n160, S => n365, Y => n1075);
   U681 : INVX2 port map( A => memory_31_4_port, Y => n362);
   U682 : MUX2X1 port map( B => n362, A => n162, S => n64, Y => n1076);
   U683 : INVX2 port map( A => memory_31_5_port, Y => n363);
   U684 : MUX2X1 port map( B => n363, A => n164, S => n365, Y => n1077);
   U685 : INVX2 port map( A => memory_31_6_port, Y => n364);
   U686 : MUX2X1 port map( B => n364, A => n166, S => n64, Y => n1078);
   U687 : INVX2 port map( A => memory_31_7_port, Y => n366);
   U688 : MUX2X1 port map( B => n366, A => n168, S => n64, Y => n1079);
   U689 : INVX2 port map( A => memory_30_0_port, Y => n367);
   U690 : MUX2X1 port map( B => n367, A => n154, S => n63, Y => n1080);
   U691 : INVX2 port map( A => memory_30_1_port, Y => n368);
   U692 : MUX2X1 port map( B => n368, A => n156, S => n374, Y => n1081);
   U693 : INVX2 port map( A => memory_30_2_port, Y => n369);
   U694 : MUX2X1 port map( B => n369, A => n158, S => n374, Y => n1082);
   U695 : INVX2 port map( A => memory_30_3_port, Y => n370);
   U696 : MUX2X1 port map( B => n370, A => n160, S => n374, Y => n1083);
   U697 : INVX2 port map( A => memory_30_4_port, Y => n371);
   U698 : MUX2X1 port map( B => n371, A => n162, S => n374, Y => n1084);
   U699 : INVX2 port map( A => memory_30_5_port, Y => n372);
   U700 : MUX2X1 port map( B => n372, A => n164, S => n374, Y => n1085);
   U701 : INVX2 port map( A => memory_30_6_port, Y => n373);
   U702 : MUX2X1 port map( B => n373, A => n166, S => n374, Y => n1086);
   U703 : INVX2 port map( A => memory_30_7_port, Y => n375);
   U704 : MUX2X1 port map( B => n375, A => n168, S => n63, Y => n1087);
   U705 : INVX2 port map( A => memory_29_0_port, Y => n376);
   U706 : MUX2X1 port map( B => n376, A => n154, S => n62, Y => n1088);
   U707 : INVX2 port map( A => memory_29_1_port, Y => n377);
   U708 : MUX2X1 port map( B => n377, A => n156, S => n383, Y => n1089);
   U709 : INVX2 port map( A => memory_29_2_port, Y => n378);
   U710 : MUX2X1 port map( B => n378, A => n158, S => n383, Y => n1090);
   U711 : INVX2 port map( A => memory_29_3_port, Y => n379);
   U712 : MUX2X1 port map( B => n379, A => n160, S => n383, Y => n1091);
   U713 : INVX2 port map( A => memory_29_4_port, Y => n380);
   U714 : MUX2X1 port map( B => n380, A => n162, S => n383, Y => n1092);
   U715 : INVX2 port map( A => memory_29_5_port, Y => n381);
   U716 : MUX2X1 port map( B => n381, A => n164, S => n383, Y => n1093);
   U717 : INVX2 port map( A => memory_29_6_port, Y => n382);
   U718 : MUX2X1 port map( B => n382, A => n166, S => n383, Y => n1094);
   U719 : INVX2 port map( A => memory_29_7_port, Y => n384);
   U720 : MUX2X1 port map( B => n384, A => n168, S => n62, Y => n1095);
   U721 : INVX2 port map( A => memory_28_0_port, Y => n385);
   U722 : MUX2X1 port map( B => n385, A => n154, S => n61, Y => n1096);
   U723 : INVX2 port map( A => memory_28_1_port, Y => n386);
   U724 : MUX2X1 port map( B => n386, A => n156, S => n392, Y => n1097);
   U725 : INVX2 port map( A => memory_28_2_port, Y => n387);
   U726 : MUX2X1 port map( B => n387, A => n158, S => n392, Y => n1098);
   U727 : INVX2 port map( A => memory_28_3_port, Y => n388);
   U728 : MUX2X1 port map( B => n388, A => n160, S => n392, Y => n1099);
   U729 : INVX2 port map( A => memory_28_4_port, Y => n389);
   U730 : MUX2X1 port map( B => n389, A => n162, S => n392, Y => n1100);
   U731 : INVX2 port map( A => memory_28_5_port, Y => n390);
   U732 : MUX2X1 port map( B => n390, A => n164, S => n392, Y => n1101);
   U733 : INVX2 port map( A => memory_28_6_port, Y => n391);
   U734 : MUX2X1 port map( B => n391, A => n166, S => n392, Y => n1102);
   U735 : INVX2 port map( A => memory_28_7_port, Y => n393);
   U736 : MUX2X1 port map( B => n393, A => n168, S => n61, Y => n1103);
   U737 : MUX2X1 port map( B => n689, A => n154, S => n24, Y => n1293);
   U738 : MUX2X1 port map( B => n688, A => n156, S => n394, Y => n1292);
   U739 : MUX2X1 port map( B => n687, A => n158, S => n24, Y => n1291);
   U740 : MUX2X1 port map( B => n686, A => n160, S => n24, Y => n1290);
   U741 : MUX2X1 port map( B => n685, A => n162, S => n394, Y => n1289);
   U742 : MUX2X1 port map( B => n684, A => n164, S => n24, Y => n1288);
   U743 : MUX2X1 port map( B => n683, A => n166, S => n24, Y => n1287);
   U744 : MUX2X1 port map( B => n682, A => n168, S => n24, Y => n1286);
   U745 : MUX2X1 port map( B => n697, A => n154, S => n60, Y => n1301);
   U746 : MUX2X1 port map( B => n696, A => n156, S => n395, Y => n1300);
   U747 : MUX2X1 port map( B => n695, A => n158, S => n395, Y => n1299);
   U748 : MUX2X1 port map( B => n694, A => n160, S => n395, Y => n1298);
   U749 : MUX2X1 port map( B => n693, A => n162, S => n395, Y => n1297);
   U750 : MUX2X1 port map( B => n692, A => n164, S => n395, Y => n1296);
   U751 : MUX2X1 port map( B => n691, A => n166, S => n395, Y => n1295);
   U752 : MUX2X1 port map( B => n690, A => n168, S => n60, Y => n1294);
   U753 : MUX2X1 port map( B => n705, A => n154, S => n59, Y => n1309);
   U754 : MUX2X1 port map( B => n704, A => n156, S => n396, Y => n1308);
   U755 : MUX2X1 port map( B => n703, A => n158, S => n396, Y => n1307);
   U756 : MUX2X1 port map( B => n702, A => n160, S => n396, Y => n1306);
   U757 : MUX2X1 port map( B => n701, A => n162, S => n396, Y => n1305);
   U758 : MUX2X1 port map( B => n700, A => n164, S => n396, Y => n1304);
   U759 : MUX2X1 port map( B => n699, A => n166, S => n396, Y => n1303);
   U760 : MUX2X1 port map( B => n698, A => n168, S => n59, Y => n1302);
   U761 : MUX2X1 port map( B => n713, A => n154, S => n93, Y => n1317);
   U762 : MUX2X1 port map( B => n712, A => n156, S => n93, Y => n1316);
   U763 : MUX2X1 port map( B => n711, A => n158, S => n93, Y => n1315);
   U764 : MUX2X1 port map( B => n710, A => n160, S => n93, Y => n1314);
   U765 : MUX2X1 port map( B => n709, A => n162, S => n93, Y => n1313);
   U766 : MUX2X1 port map( B => n708, A => n164, S => n93, Y => n1312);
   U767 : MUX2X1 port map( B => n707, A => n166, S => n93, Y => n1311);
   U768 : MUX2X1 port map( B => n706, A => n168, S => n92, Y => n1310);
   U769 : INVX2 port map( A => memory_23_0_port, Y => n397);
   U770 : MUX2X1 port map( B => n397, A => n154, S => n34, Y => n1325);
   U771 : INVX2 port map( A => memory_23_1_port, Y => n398);
   U772 : MUX2X1 port map( B => n398, A => n156, S => n34, Y => n1324);
   U773 : INVX2 port map( A => memory_23_2_port, Y => n399);
   U774 : MUX2X1 port map( B => n399, A => n158, S => n34, Y => n1323);
   U775 : INVX2 port map( A => memory_23_3_port, Y => n400);
   U776 : MUX2X1 port map( B => n400, A => n160, S => n404, Y => n1322);
   U777 : INVX2 port map( A => memory_23_4_port, Y => n401);
   U778 : MUX2X1 port map( B => n401, A => n162, S => n34, Y => n1321);
   U779 : INVX2 port map( A => memory_23_5_port, Y => n402);
   U780 : MUX2X1 port map( B => n402, A => n164, S => n404, Y => n1320);
   U781 : INVX2 port map( A => memory_23_6_port, Y => n403);
   U782 : MUX2X1 port map( B => n403, A => n166, S => n34, Y => n1319);
   U783 : INVX2 port map( A => memory_23_7_port, Y => n405);
   U784 : MUX2X1 port map( B => n405, A => n168, S => n34, Y => n1318);
   U785 : INVX2 port map( A => memory_22_0_port, Y => n406);
   U786 : MUX2X1 port map( B => n406, A => n154, S => n33, Y => n1333);
   U787 : INVX2 port map( A => memory_22_1_port, Y => n407);
   U788 : MUX2X1 port map( B => n407, A => n156, S => n1, Y => n1332);
   U789 : INVX2 port map( A => memory_22_2_port, Y => n408);
   U790 : MUX2X1 port map( B => n408, A => n158, S => n33, Y => n1331);
   U791 : INVX2 port map( A => memory_22_3_port, Y => n409);
   U792 : MUX2X1 port map( B => n409, A => n160, S => n33, Y => n1330);
   U793 : INVX2 port map( A => memory_22_4_port, Y => n410);
   U794 : MUX2X1 port map( B => n410, A => n162, S => n1, Y => n1329);
   U795 : INVX2 port map( A => memory_22_5_port, Y => n411);
   U796 : MUX2X1 port map( B => n411, A => n164, S => n33, Y => n1328);
   U797 : INVX2 port map( A => memory_22_6_port, Y => n412);
   U798 : MUX2X1 port map( B => n412, A => n166, S => n33, Y => n1327);
   U799 : INVX2 port map( A => memory_22_7_port, Y => n413);
   U800 : MUX2X1 port map( B => n413, A => n168, S => n33, Y => n1326);
   U801 : INVX2 port map( A => memory_21_0_port, Y => n414);
   U802 : MUX2X1 port map( B => n414, A => n154, S => n45, Y => n1341);
   U803 : INVX2 port map( A => memory_21_1_port, Y => n415);
   U804 : MUX2X1 port map( B => n415, A => n156, S => n46, Y => n1340);
   U805 : INVX2 port map( A => memory_21_2_port, Y => n416);
   U806 : MUX2X1 port map( B => n416, A => n158, S => n45, Y => n1339);
   U807 : INVX2 port map( A => memory_21_3_port, Y => n417);
   U808 : MUX2X1 port map( B => n417, A => n160, S => n46, Y => n1338);
   U809 : INVX2 port map( A => memory_21_4_port, Y => n418);
   U810 : MUX2X1 port map( B => n418, A => n162, S => n45, Y => n1337);
   U811 : INVX2 port map( A => memory_21_5_port, Y => n419);
   U812 : MUX2X1 port map( B => n419, A => n164, S => n46, Y => n1336);
   U813 : INVX2 port map( A => memory_21_6_port, Y => n420);
   U814 : MUX2X1 port map( B => n420, A => n166, S => n45, Y => n1335);
   U815 : INVX2 port map( A => memory_21_7_port, Y => n422);
   U816 : MUX2X1 port map( B => n422, A => n168, S => n46, Y => n1334);
   U817 : INVX2 port map( A => memory_20_0_port, Y => n423);
   U818 : MUX2X1 port map( B => n423, A => n154, S => n44, Y => n1349);
   U819 : INVX2 port map( A => memory_20_1_port, Y => n424);
   U820 : MUX2X1 port map( B => n424, A => n156, S => n430, Y => n1348);
   U821 : INVX2 port map( A => memory_20_2_port, Y => n425);
   U822 : MUX2X1 port map( B => n425, A => n158, S => n44, Y => n1347);
   U823 : INVX2 port map( A => memory_20_3_port, Y => n426);
   U824 : MUX2X1 port map( B => n426, A => n160, S => n44, Y => n1346);
   U825 : INVX2 port map( A => memory_20_4_port, Y => n427);
   U826 : MUX2X1 port map( B => n427, A => n162, S => n44, Y => n1345);
   U827 : INVX2 port map( A => memory_20_5_port, Y => n428);
   U828 : MUX2X1 port map( B => n428, A => n164, S => n44, Y => n1344);
   U829 : INVX2 port map( A => memory_20_6_port, Y => n429);
   U830 : MUX2X1 port map( B => n429, A => n166, S => n44, Y => n1343);
   U831 : INVX2 port map( A => memory_20_7_port, Y => n431);
   U832 : MUX2X1 port map( B => n431, A => n168, S => n430, Y => n1342);
   U833 : MUX2X1 port map( B => n811, A => n154, S => n56, Y => n1104);
   U834 : MUX2X1 port map( B => n810, A => n156, S => n56, Y => n1105);
   U835 : MUX2X1 port map( B => n809, A => n159, S => n56, Y => n1106);
   U836 : MUX2X1 port map( B => n808, A => n160, S => n432, Y => n1107);
   U837 : MUX2X1 port map( B => n807, A => n162, S => n56, Y => n1108);
   U838 : MUX2X1 port map( B => n806, A => n164, S => n432, Y => n1109);
   U839 : MUX2X1 port map( B => n805, A => n166, S => n56, Y => n1110);
   U840 : MUX2X1 port map( B => n804, A => n168, S => n56, Y => n1111);
   U841 : MUX2X1 port map( B => n803, A => n154, S => n42, Y => n1112);
   U842 : MUX2X1 port map( B => n802, A => n156, S => n43, Y => n1113);
   U843 : MUX2X1 port map( B => n801, A => n159, S => n42, Y => n1114);
   U844 : MUX2X1 port map( B => n800, A => n160, S => n43, Y => n1115);
   U845 : MUX2X1 port map( B => n799, A => n162, S => n42, Y => n1116);
   U846 : MUX2X1 port map( B => n798, A => n164, S => n43, Y => n1117);
   U847 : MUX2X1 port map( B => n797, A => n166, S => n42, Y => n1118);
   U848 : MUX2X1 port map( B => n796, A => n168, S => n43, Y => n1119);
   U849 : MUX2X1 port map( B => n795, A => n154, S => n73, Y => n1120);
   U850 : MUX2X1 port map( B => n794, A => n156, S => n73, Y => n1121);
   U851 : MUX2X1 port map( B => n793, A => n159, S => n32, Y => n1122);
   U852 : MUX2X1 port map( B => n792, A => n160, S => n32, Y => n1123);
   U853 : MUX2X1 port map( B => n791, A => n162, S => n32, Y => n1124);
   U854 : MUX2X1 port map( B => n790, A => n164, S => n73, Y => n1125);
   U855 : MUX2X1 port map( B => n789, A => n166, S => n32, Y => n1126);
   U856 : MUX2X1 port map( B => n788, A => n168, S => n73, Y => n1127);
   U857 : MUX2X1 port map( B => n787, A => n154, S => n31, Y => n1128);
   U858 : MUX2X1 port map( B => n786, A => n156, S => n31, Y => n1129);
   U859 : MUX2X1 port map( B => n785, A => n159, S => n31, Y => n1130);
   U860 : MUX2X1 port map( B => n784, A => n160, S => n434, Y => n1131);
   U861 : MUX2X1 port map( B => n783, A => n162, S => n31, Y => n1132);
   U862 : MUX2X1 port map( B => n782, A => n164, S => n434, Y => n1133);
   U863 : MUX2X1 port map( B => n781, A => n166, S => n31, Y => n1134);
   U864 : MUX2X1 port map( B => n780, A => n168, S => n31, Y => n1135);
   U865 : INVX2 port map( A => memory_15_0_port, Y => n435);
   U866 : MUX2X1 port map( B => n435, A => n154, S => n67, Y => n1357);
   U867 : INVX2 port map( A => memory_15_1_port, Y => n436);
   U868 : MUX2X1 port map( B => n436, A => n156, S => n67, Y => n1356);
   U869 : INVX2 port map( A => memory_15_2_port, Y => n437);
   U870 : MUX2X1 port map( B => n437, A => n159, S => n67, Y => n1355);
   U871 : INVX2 port map( A => memory_15_3_port, Y => n438);
   U872 : MUX2X1 port map( B => n438, A => n160, S => n442, Y => n1354);
   U873 : INVX2 port map( A => memory_15_4_port, Y => n439);
   U874 : MUX2X1 port map( B => n439, A => n162, S => n67, Y => n1353);
   U875 : INVX2 port map( A => memory_15_5_port, Y => n440);
   U876 : MUX2X1 port map( B => n440, A => n164, S => n442, Y => n1352);
   U877 : INVX2 port map( A => memory_15_6_port, Y => n441);
   U878 : MUX2X1 port map( B => n441, A => n166, S => n67, Y => n1351);
   U879 : INVX2 port map( A => memory_15_7_port, Y => n443);
   U880 : MUX2X1 port map( B => n443, A => n168, S => n67, Y => n1350);
   U881 : INVX2 port map( A => memory_14_0_port, Y => n444);
   U882 : MUX2X1 port map( B => n444, A => n154, S => n65, Y => n1365);
   U883 : INVX2 port map( A => memory_14_1_port, Y => n445);
   U884 : MUX2X1 port map( B => n445, A => n156, S => n451, Y => n1364);
   U885 : INVX2 port map( A => memory_14_2_port, Y => n446);
   U886 : MUX2X1 port map( B => n446, A => n159, S => n65, Y => n1363);
   U887 : INVX2 port map( A => memory_14_3_port, Y => n447);
   U888 : MUX2X1 port map( B => n447, A => n160, S => n65, Y => n1362);
   U889 : INVX2 port map( A => memory_14_4_port, Y => n448);
   U890 : MUX2X1 port map( B => n448, A => n518, S => n65, Y => n1361);
   U891 : INVX2 port map( A => memory_14_5_port, Y => n449);
   U892 : MUX2X1 port map( B => n449, A => n164, S => n65, Y => n1360);
   U893 : INVX2 port map( A => memory_14_6_port, Y => n450);
   U894 : MUX2X1 port map( B => n450, A => n520, S => n65, Y => n1359);
   U895 : INVX2 port map( A => memory_14_7_port, Y => n452);
   U896 : MUX2X1 port map( B => n452, A => n521, S => n65, Y => n1358);
   U897 : INVX2 port map( A => memory_13_0_port, Y => n453);
   U898 : MUX2X1 port map( B => n453, A => n154, S => n460, Y => n1373);
   U899 : INVX2 port map( A => memory_13_1_port, Y => n454);
   U900 : MUX2X1 port map( B => n454, A => n156, S => n460, Y => n1372);
   U901 : INVX2 port map( A => memory_13_2_port, Y => n455);
   U902 : MUX2X1 port map( B => n455, A => n159, S => n460, Y => n1371);
   U903 : INVX2 port map( A => memory_13_3_port, Y => n456);
   U904 : MUX2X1 port map( B => n456, A => n160, S => n460, Y => n1370);
   U905 : INVX2 port map( A => memory_13_4_port, Y => n457);
   U906 : MUX2X1 port map( B => n457, A => n518, S => n460, Y => n1369);
   U907 : INVX2 port map( A => memory_13_5_port, Y => n458);
   U908 : MUX2X1 port map( B => n458, A => n164, S => n460, Y => n1368);
   U909 : INVX2 port map( A => memory_13_6_port, Y => n459);
   U910 : MUX2X1 port map( B => n459, A => n520, S => n460, Y => n1367);
   U911 : INVX2 port map( A => memory_13_7_port, Y => n461);
   U912 : MUX2X1 port map( B => n461, A => n521, S => n460, Y => n1366);
   U913 : INVX2 port map( A => memory_12_0_port, Y => n462);
   U914 : MUX2X1 port map( B => n462, A => n515, S => n469, Y => n1381);
   U915 : INVX2 port map( A => memory_12_1_port, Y => n463);
   U916 : MUX2X1 port map( B => n463, A => n516, S => n469, Y => n1380);
   U917 : INVX2 port map( A => memory_12_2_port, Y => n464);
   U918 : MUX2X1 port map( B => n464, A => n159, S => n469, Y => n1379);
   U919 : INVX2 port map( A => memory_12_3_port, Y => n465);
   U920 : MUX2X1 port map( B => n465, A => n517, S => n469, Y => n1378);
   U921 : INVX2 port map( A => memory_12_4_port, Y => n466);
   U922 : MUX2X1 port map( B => n466, A => n518, S => n469, Y => n1377);
   U923 : INVX2 port map( A => memory_12_5_port, Y => n467);
   U924 : MUX2X1 port map( B => n467, A => n519, S => n469, Y => n1376);
   U925 : INVX2 port map( A => memory_12_6_port, Y => n468);
   U926 : MUX2X1 port map( B => n468, A => n520, S => n469, Y => n1375);
   U927 : INVX2 port map( A => memory_12_7_port, Y => n470);
   U928 : MUX2X1 port map( B => n470, A => n521, S => n469, Y => n1374);
   U929 : MUX2X1 port map( B => n779, A => n515, S => n97, Y => n1136);
   U930 : MUX2X1 port map( B => n778, A => n516, S => n97, Y => n1137);
   U931 : MUX2X1 port map( B => n777, A => n159, S => n97, Y => n1138);
   U932 : MUX2X1 port map( B => n776, A => n517, S => n97, Y => n1139);
   U933 : MUX2X1 port map( B => n775, A => n518, S => n97, Y => n1140);
   U934 : MUX2X1 port map( B => n774, A => n519, S => n97, Y => n1141);
   U935 : MUX2X1 port map( B => n773, A => n520, S => n97, Y => n1142);
   U936 : MUX2X1 port map( B => n772, A => n521, S => n97, Y => n1143);
   U937 : MUX2X1 port map( B => n771, A => n515, S => n473, Y => n1144);
   U938 : MUX2X1 port map( B => n770, A => n516, S => n473, Y => n1145);
   U939 : MUX2X1 port map( B => n769, A => n159, S => n473, Y => n1146);
   U940 : MUX2X1 port map( B => n768, A => n517, S => n473, Y => n1147);
   U941 : MUX2X1 port map( B => n767, A => n518, S => n473, Y => n1148);
   U942 : MUX2X1 port map( B => n766, A => n519, S => n473, Y => n1149);
   U943 : MUX2X1 port map( B => n765, A => n520, S => n473, Y => n1150);
   U944 : MUX2X1 port map( B => n764, A => n521, S => n473, Y => n1151);
   U945 : MUX2X1 port map( B => n763, A => n154, S => n474, Y => n1152);
   U946 : MUX2X1 port map( B => n762, A => n156, S => n474, Y => n1153);
   U947 : MUX2X1 port map( B => n761, A => n159, S => n474, Y => n1154);
   U948 : MUX2X1 port map( B => n760, A => n160, S => n474, Y => n1155);
   U949 : MUX2X1 port map( B => n759, A => n518, S => n474, Y => n1156);
   U950 : MUX2X1 port map( B => n758, A => n164, S => n474, Y => n1157);
   U951 : MUX2X1 port map( B => n757, A => n520, S => n474, Y => n1158);
   U952 : MUX2X1 port map( B => n756, A => n521, S => n474, Y => n1159);
   U953 : MUX2X1 port map( B => n755, A => n154, S => n475, Y => n1160);
   U954 : MUX2X1 port map( B => n754, A => n156, S => n475, Y => n1161);
   U955 : MUX2X1 port map( B => n753, A => n159, S => n475, Y => n1162);
   U956 : MUX2X1 port map( B => n752, A => n160, S => n475, Y => n1163);
   U957 : MUX2X1 port map( B => n751, A => n518, S => n475, Y => n1164);
   U958 : MUX2X1 port map( B => n750, A => n164, S => n475, Y => n1165);
   U959 : MUX2X1 port map( B => n749, A => n520, S => n475, Y => n1166);
   U960 : MUX2X1 port map( B => n748, A => n521, S => n475, Y => n1167);
   U961 : INVX2 port map( A => memory_7_0_port, Y => n476);
   U962 : MUX2X1 port map( B => n476, A => n515, S => n127, Y => n906);
   U963 : INVX2 port map( A => memory_7_1_port, Y => n477);
   U964 : MUX2X1 port map( B => n477, A => n516, S => n127, Y => n905);
   U965 : INVX2 port map( A => memory_7_2_port, Y => n478);
   U966 : MUX2X1 port map( B => n478, A => n159, S => n127, Y => n904);
   U967 : INVX2 port map( A => memory_7_3_port, Y => n479);
   U968 : MUX2X1 port map( B => n479, A => n517, S => n127, Y => n903);
   U969 : INVX2 port map( A => memory_7_4_port, Y => n480);
   U970 : MUX2X1 port map( B => n480, A => n518, S => n127, Y => n902);
   U971 : INVX2 port map( A => memory_7_5_port, Y => n481);
   U972 : MUX2X1 port map( B => n481, A => n519, S => n127, Y => n901);
   U973 : INVX2 port map( A => memory_7_6_port, Y => n482);
   U974 : MUX2X1 port map( B => n482, A => n520, S => n127, Y => n900);
   U975 : INVX2 port map( A => memory_7_7_port, Y => n484);
   U976 : MUX2X1 port map( B => n484, A => n521, S => n127, Y => n899);
   U977 : INVX2 port map( A => memory_6_0_port, Y => n485);
   U978 : MUX2X1 port map( B => n485, A => n515, S => n57, Y => n896);
   U979 : INVX2 port map( A => memory_6_1_port, Y => n486);
   U980 : MUX2X1 port map( B => n486, A => n516, S => n492, Y => n895);
   U981 : INVX2 port map( A => memory_6_2_port, Y => n487);
   U982 : MUX2X1 port map( B => n487, A => n158, S => n58, Y => n894);
   U983 : INVX2 port map( A => memory_6_3_port, Y => n488);
   U984 : MUX2X1 port map( B => n488, A => n517, S => n57, Y => n893);
   U985 : INVX2 port map( A => memory_6_4_port, Y => n489);
   U986 : MUX2X1 port map( B => n489, A => n518, S => n57, Y => n892);
   U987 : INVX2 port map( A => memory_6_5_port, Y => n490);
   U988 : MUX2X1 port map( B => n490, A => n519, S => n58, Y => n891);
   U989 : INVX2 port map( A => memory_6_6_port, Y => n491);
   U990 : MUX2X1 port map( B => n491, A => n520, S => n57, Y => n890);
   U991 : INVX2 port map( A => memory_6_7_port, Y => n493);
   U992 : MUX2X1 port map( B => n493, A => n521, S => n58, Y => n889);
   U993 : INVX2 port map( A => memory_5_0_port, Y => n494);
   U994 : MUX2X1 port map( B => n494, A => n515, S => n66, Y => n886);
   U995 : INVX2 port map( A => memory_5_1_port, Y => n495);
   U996 : MUX2X1 port map( B => n495, A => n516, S => n66, Y => n885);
   U997 : INVX2 port map( A => memory_5_2_port, Y => n496);
   U998 : MUX2X1 port map( B => n496, A => n159, S => n66, Y => n884);
   U999 : INVX2 port map( A => memory_5_3_port, Y => n497);
   U1000 : MUX2X1 port map( B => n497, A => n517, S => n66, Y => n883);
   U1001 : INVX2 port map( A => memory_5_4_port, Y => n498);
   U1002 : MUX2X1 port map( B => n498, A => n518, S => n66, Y => n882);
   U1003 : INVX2 port map( A => memory_5_5_port, Y => n499);
   U1004 : MUX2X1 port map( B => n499, A => n519, S => n66, Y => n881);
   U1005 : INVX2 port map( A => memory_5_6_port, Y => n500);
   U1006 : MUX2X1 port map( B => n500, A => n520, S => n66, Y => n880);
   U1007 : INVX2 port map( A => memory_5_7_port, Y => n502);
   U1008 : MUX2X1 port map( B => n502, A => n521, S => n66, Y => n879);
   U1009 : INVX2 port map( A => memory_4_0_port, Y => n503);
   U1010 : MUX2X1 port map( B => n503, A => n515, S => n39, Y => n876);
   U1011 : INVX2 port map( A => memory_4_1_port, Y => n504);
   U1012 : MUX2X1 port map( B => n504, A => n516, S => n71, Y => n875);
   U1013 : INVX2 port map( A => memory_4_2_port, Y => n505);
   U1014 : MUX2X1 port map( B => n505, A => n158, S => n39, Y => n874);
   U1015 : INVX2 port map( A => memory_4_3_port, Y => n506);
   U1016 : MUX2X1 port map( B => n506, A => n517, S => n71, Y => n873);
   U1017 : INVX2 port map( A => memory_4_4_port, Y => n507);
   U1018 : MUX2X1 port map( B => n507, A => n518, S => n510, Y => n872);
   U1019 : INVX2 port map( A => memory_4_5_port, Y => n508);
   U1020 : MUX2X1 port map( B => n508, A => n519, S => n39, Y => n871);
   U1021 : INVX2 port map( A => memory_4_6_port, Y => n509);
   U1022 : MUX2X1 port map( B => n509, A => n520, S => n71, Y => n870);
   U1023 : INVX2 port map( A => memory_4_7_port, Y => n511);
   U1024 : MUX2X1 port map( B => n511, A => n521, S => n510, Y => n869);
   U1025 : MUX2X1 port map( B => n738, A => n515, S => n47, Y => n1406);
   U1026 : MUX2X1 port map( B => n739, A => n516, S => n3, Y => n1407);
   U1027 : MUX2X1 port map( B => n740, A => n159, S => n3, Y => n1408);
   U1028 : MUX2X1 port map( B => n741, A => n517, S => n3, Y => n1409);
   U1029 : MUX2X1 port map( B => n742, A => n162, S => n47, Y => n1410);
   U1030 : MUX2X1 port map( B => n743, A => n519, S => n3, Y => n1411);
   U1031 : MUX2X1 port map( B => n744, A => n166, S => n47, Y => n1412);
   U1032 : MUX2X1 port map( B => n745, A => n168, S => n3, Y => n1413);
   U1033 : MUX2X1 port map( B => n730, A => n515, S => n513, Y => n1398);
   U1034 : MUX2X1 port map( B => n731, A => n516, S => n513, Y => n1399);
   U1035 : MUX2X1 port map( B => n732, A => n158, S => n40, Y => n1400);
   U1036 : MUX2X1 port map( B => n733, A => n517, S => n40, Y => n1401);
   U1037 : MUX2X1 port map( B => n734, A => n162, S => n513, Y => n1402);
   U1038 : MUX2X1 port map( B => n735, A => n519, S => n40, Y => n1403);
   U1039 : MUX2X1 port map( B => n736, A => n166, S => n513, Y => n1404);
   U1040 : MUX2X1 port map( B => n737, A => n168, S => n40, Y => n1405);
   U1041 : MUX2X1 port map( B => n722, A => n515, S => n48, Y => n1390);
   U1042 : MUX2X1 port map( B => n723, A => n516, S => n4, Y => n1391);
   U1043 : MUX2X1 port map( B => n724, A => n159, S => n4, Y => n1392);
   U1044 : MUX2X1 port map( B => n725, A => n517, S => n4, Y => n1393);
   U1045 : MUX2X1 port map( B => n726, A => n162, S => n48, Y => n1394);
   U1046 : MUX2X1 port map( B => n727, A => n519, S => n4, Y => n1395);
   U1047 : MUX2X1 port map( B => n728, A => n166, S => n48, Y => n1396);
   U1048 : MUX2X1 port map( B => n729, A => n168, S => n4, Y => n1397);
   U1049 : MUX2X1 port map( B => n714, A => n515, S => n79, Y => n1382);
   U1050 : MUX2X1 port map( B => n715, A => n516, S => n80, Y => n1383);
   U1051 : MUX2X1 port map( B => n716, A => n158, S => n70, Y => n1384);
   U1052 : MUX2X1 port map( B => n717, A => n517, S => n80, Y => n1385);
   U1053 : MUX2X1 port map( B => n718, A => n162, S => n79, Y => n1386);
   U1054 : MUX2X1 port map( B => n719, A => n519, S => n70, Y => n1387);
   U1055 : MUX2X1 port map( B => n720, A => n166, S => n70, Y => n1388);
   U1056 : MUX2X1 port map( B => n721, A => n168, S => n80, Y => n1389);
   U1057 : AND2X2 port map( A => state, B => n522, Y => N338);
   U1058 : XOR2X1 port map( A => n524, B => n123, Y => n523);
   U1059 : INVX2 port map( A => state, Y => n598);
   U1060 : NOR2X1 port map( A => n523, B => n598, Y => N339);
   U1061 : NAND2X1 port map( A => n77, B => n594, Y => n526);
   U1062 : OAI21X1 port map( A => n77, B => n594, C => n524, Y => n525);
   U1063 : AND2X2 port map( A => n526, B => n525, Y => n531);
   U1064 : XNOR2X1 port map( A => n531, B => n527, Y => n528);
   U1065 : AND2X2 port map( A => state, B => n528, Y => N340);
   U1066 : NOR2X1 port map( A => n149, B => n663, Y => n530);
   U1067 : NAND2X1 port map( A => n149, B => n663, Y => n529);
   U1068 : OAI21X1 port map( A => n531, B => n530, C => n529, Y => n535);
   U1069 : XNOR2X1 port map( A => n535, B => n532, Y => n533);
   U1070 : NOR2X1 port map( A => n533, B => n598, Y => N341);
   U1071 : NAND2X1 port map( A => n153, B => n568, Y => n536);
   U1072 : NOR2X1 port map( A => n153, B => n568, Y => n534);
   U1073 : AOI21X1 port map( A => n536, B => n535, C => n534, Y => n538);
   U1074 : XNOR2X1 port map( A => n538, B => n28, Y => n539);
   U1075 : AND2X2 port map( A => state, B => n539, Y => N342);
   U1076 : NOR2X1 port map( A => n85, B => n540, Y => n545);
   U1077 : AND2X2 port map( A => n6, B => n541, Y => n543);
   U1078 : NAND3X1 port map( A => n545, B => n544, C => n543, Y => n546);
   U1079 : MUX2X1 port map( B => n546, A => n746, S => RST, Y => n1414);
   U1080 : NAND2X1 port map( A => n89, B => n38, Y => n562);
   U1081 : INVX2 port map( A => n562, Y => n576);
   U1082 : NAND2X1 port map( A => n576, B => n27, Y => n552);
   U1083 : NAND2X1 port map( A => n149, B => n556, Y => n548);
   U1084 : NAND2X1 port map( A => n548, B => n565, Y => n549);
   U1085 : NAND2X1 port map( A => n578, B => n549, Y => n551);
   U1086 : NAND2X1 port map( A => n149, B => n558, Y => n550);
   U1087 : NAND3X1 port map( A => n552, B => n551, C => n550, Y => n854);
   U1088 : NAND2X1 port map( A => n576, B => n554, Y => n561);
   U1089 : NAND2X1 port map( A => n556, B => n72, Y => n557);
   U1090 : NAND2X1 port map( A => n578, B => n557, Y => n560);
   U1091 : NAND2X1 port map( A => n77, B => n558, Y => n559);
   U1092 : NAND3X1 port map( A => n561, B => n560, C => n559, Y => n856);
   U1093 : MUX2X1 port map( B => n564, A => n89, S => n52, Y => n858);
   U1094 : NAND2X1 port map( A => n566, B => n565, Y => n579);
   U1095 : NAND2X1 port map( A => n89, B => n579, Y => n567);
   U1096 : NAND2X1 port map( A => n94, B => n567, Y => n572);
   U1097 : XNOR2X1 port map( A => n569, B => n568, Y => n570);
   U1098 : NAND2X1 port map( A => n570, B => n576, Y => n571);
   U1099 : NAND3X1 port map( A => n572, B => n577, C => n571, Y => n860);
   U1100 : XOR2X1 port map( A => n574, B => n8, Y => n575);
   U1101 : NAND2X1 port map( A => n576, B => n575, Y => n585);
   U1102 : NAND2X1 port map( A => n578, B => n94, Y => n580);
   U1103 : NAND3X1 port map( A => n89, B => n580, C => n579, Y => n582);
   U1104 : MUX2X1 port map( B => n583, A => n582, S => n49, Y => n584);
   U1105 : NAND2X1 port map( A => n585, B => n584, Y => n862);
   U1106 : NAND2X1 port map( A => n81, B => n76, Y => n595);
   U1107 : INVX2 port map( A => n595, Y => n591);
   U1108 : NAND2X1 port map( A => n121, B => n591, Y => n589);
   U1109 : INVX2 port map( A => n589, Y => n586);
   U1110 : NAND2X1 port map( A => n586, B => n153, Y => n587);
   U1111 : XNOR2X1 port map( A => n587, B => n665, Y => n588);
   U1112 : NOR2X1 port map( A => n598, B => n588, Y => N347);
   U1113 : XNOR2X1 port map( A => n589, B => n664, Y => n590);
   U1114 : NOR2X1 port map( A => n598, B => n590, Y => N346);
   U1115 : NAND2X1 port map( A => n120, B => n591, Y => n593);
   U1116 : OAI21X1 port map( A => n595, B => n594, C => n36, Y => n592);
   U1117 : AOI21X1 port map( A => n593, B => n592, C => n598, Y => N345);
   U1118 : XNOR2X1 port map( A => n595, B => n594, Y => n596);
   U1119 : NOR2X1 port map( A => n598, B => n596, Y => N344);
   U1120 : XNOR2X1 port map( A => n597, B => n662, Y => n599);
   U1121 : NOR2X1 port map( A => n599, B => n598, Y => N343);
   U1122 : INVX1 port map( A => FULL_port, Y => n746);
   U1123 : INVX1 port map( A => EMPTY_port, Y => n747);
   U1124 : NAND2X1 port map( A => n829, B => n830, Y => n828);
   U1125 : NOR2X1 port map( A => n831, B => n832, Y => n830);
   U1126 : NAND3X1 port map( A => n833, B => n834, C => n835, Y => n832);
   U1127 : NOR2X1 port map( A => n836, B => n837, Y => n835);
   U1128 : OAI22X1 port map( A => n780, B => n141, C => n788, D => n140, Y => 
                           n837);
   U1129 : OAI22X1 port map( A => n796, B => n128, C => n804, D => n130, Y => 
                           n836);
   U1130 : AOI22X1 port map( A => n114, B => memory_23_7_port, C => n110, D => 
                           memory_22_7_port, Y => n834);
   U1131 : AOI22X1 port map( A => n840, B => memory_21_7_port, C => n841, D => 
                           memory_20_7_port, Y => n833);
   U1132 : NAND3X1 port map( A => n842, B => n843, C => n844, Y => n831);
   U1133 : NOR2X1 port map( A => n845, B => n846, Y => n844);
   U1134 : OAI22X1 port map( A => n706, B => n143, C => n698, D => n142, Y => 
                           n846);
   U1135 : OAI22X1 port map( A => n690, B => n131, C => n682, D => n132, Y => 
                           n845);
   U1136 : AOI22X1 port map( A => n115, B => memory_31_7_port, C => n112, D => 
                           memory_30_7_port, Y => n843);
   U1137 : AOI22X1 port map( A => n852, B => memory_29_7_port, C => n865, D => 
                           memory_28_7_port, Y => n842);
   U1138 : NOR2X1 port map( A => n877, B => n878, Y => n829);
   U1139 : NAND3X1 port map( A => n887, B => n888, C => n897, Y => n878);
   U1140 : NOR2X1 port map( A => n898, B => n907, Y => n897);
   U1141 : OAI22X1 port map( A => n745, B => n133, C => n737, D => n134, Y => 
                           n907);
   U1142 : OAI22X1 port map( A => n729, B => n145, C => n721, D => n144, Y => 
                           n898);
   U1143 : AOI22X1 port map( A => n908, B => memory_4_7_port, C => n909, D => 
                           memory_5_7_port, Y => n888);
   U1144 : AOI22X1 port map( A => n116, B => memory_6_7_port, C => n111, D => 
                           memory_7_7_port, Y => n887);
   U1145 : NAND3X1 port map( A => n910, B => n911, C => n912, Y => n877);
   U1146 : NOR2X1 port map( A => n913, B => n914, Y => n912);
   U1147 : OAI22X1 port map( A => n748, B => n147, C => n756, D => n146, Y => 
                           n914);
   U1148 : OAI22X1 port map( A => n764, B => n135, C => n772, D => n136, Y => 
                           n913);
   U1149 : AOI22X1 port map( A => n113, B => memory_15_7_port, C => n109, D => 
                           memory_14_7_port, Y => n911);
   U1150 : AOI22X1 port map( A => n915, B => memory_13_7_port, C => n916, D => 
                           memory_12_7_port, Y => n910);
   U1151 : NAND2X1 port map( A => n918, B => n919, Y => n917);
   U1152 : NOR2X1 port map( A => n920, B => n921, Y => n919);
   U1153 : NAND3X1 port map( A => n922, B => n923, C => n924, Y => n921);
   U1154 : NOR2X1 port map( A => n925, B => n926, Y => n924);
   U1155 : OAI22X1 port map( A => n781, B => n141, C => n789, D => n140, Y => 
                           n926);
   U1156 : OAI22X1 port map( A => n797, B => n128, C => n805, D => n130, Y => 
                           n925);
   U1157 : AOI22X1 port map( A => n114, B => memory_23_6_port, C => n110, D => 
                           memory_22_6_port, Y => n923);
   U1158 : AOI22X1 port map( A => n840, B => memory_21_6_port, C => n841, D => 
                           memory_20_6_port, Y => n922);
   U1159 : NAND3X1 port map( A => n927, B => n928, C => n929, Y => n920);
   U1160 : NOR2X1 port map( A => n930, B => n931, Y => n929);
   U1161 : OAI22X1 port map( A => n707, B => n143, C => n699, D => n142, Y => 
                           n931);
   U1162 : OAI22X1 port map( A => n691, B => n131, C => n683, D => n132, Y => 
                           n930);
   U1163 : AOI22X1 port map( A => n115, B => memory_31_6_port, C => n112, D => 
                           memory_30_6_port, Y => n928);
   U1164 : AOI22X1 port map( A => n852, B => memory_29_6_port, C => n865, D => 
                           memory_28_6_port, Y => n927);
   U1165 : NOR2X1 port map( A => n932, B => n933, Y => n918);
   U1166 : NAND3X1 port map( A => n934, B => n935, C => n936, Y => n933);
   U1167 : NOR2X1 port map( A => n937, B => n938, Y => n936);
   U1168 : OAI22X1 port map( A => n744, B => n133, C => n736, D => n134, Y => 
                           n938);
   U1169 : OAI22X1 port map( A => n728, B => n145, C => n720, D => n144, Y => 
                           n937);
   U1170 : AOI22X1 port map( A => n908, B => memory_4_6_port, C => n909, D => 
                           memory_5_6_port, Y => n935);
   U1171 : AOI22X1 port map( A => n116, B => memory_6_6_port, C => n111, D => 
                           memory_7_6_port, Y => n934);
   U1172 : NAND3X1 port map( A => n939, B => n940, C => n941, Y => n932);
   U1173 : NOR2X1 port map( A => n942, B => n943, Y => n941);
   U1174 : OAI22X1 port map( A => n749, B => n147, C => n757, D => n146, Y => 
                           n943);
   U1175 : OAI22X1 port map( A => n765, B => n135, C => n773, D => n136, Y => 
                           n942);
   U1176 : AOI22X1 port map( A => n113, B => memory_15_6_port, C => n109, D => 
                           memory_14_6_port, Y => n940);
   U1177 : AOI22X1 port map( A => n915, B => memory_13_6_port, C => n916, D => 
                           memory_12_6_port, Y => n939);
   U1178 : NAND2X1 port map( A => n945, B => n946, Y => n944);
   U1179 : NOR2X1 port map( A => n947, B => n948, Y => n946);
   U1180 : NAND3X1 port map( A => n949, B => n950, C => n951, Y => n948);
   U1181 : NOR2X1 port map( A => n952, B => n953, Y => n951);
   U1182 : OAI22X1 port map( A => n782, B => n141, C => n790, D => n140, Y => 
                           n953);
   U1183 : OAI22X1 port map( A => n798, B => n128, C => n806, D => n130, Y => 
                           n952);
   U1184 : AOI22X1 port map( A => n114, B => memory_23_5_port, C => n110, D => 
                           memory_22_5_port, Y => n950);
   U1185 : AOI22X1 port map( A => n840, B => memory_21_5_port, C => n841, D => 
                           memory_20_5_port, Y => n949);
   U1186 : NAND3X1 port map( A => n954, B => n955, C => n956, Y => n947);
   U1187 : NOR2X1 port map( A => n957, B => n958, Y => n956);
   U1188 : OAI22X1 port map( A => n708, B => n143, C => n700, D => n142, Y => 
                           n958);
   U1189 : OAI22X1 port map( A => n692, B => n131, C => n684, D => n132, Y => 
                           n957);
   U1190 : AOI22X1 port map( A => n115, B => memory_31_5_port, C => n112, D => 
                           memory_30_5_port, Y => n955);
   U1203 : AOI22X1 port map( A => n852, B => memory_29_5_port, C => n865, D => 
                           memory_28_5_port, Y => n954);
   U1207 : NOR2X1 port map( A => n959, B => n960, Y => n945);
   U1208 : NAND3X1 port map( A => n961, B => n962, C => n963, Y => n960);
   U1209 : NOR2X1 port map( A => n964, B => n965, Y => n963);
   U1210 : OAI22X1 port map( A => n743, B => n133, C => n735, D => n134, Y => 
                           n965);
   U1211 : OAI22X1 port map( A => n727, B => n145, C => n719, D => n144, Y => 
                           n964);
   U1212 : AOI22X1 port map( A => n908, B => memory_4_5_port, C => n909, D => 
                           memory_5_5_port, Y => n962);
   U1213 : AOI22X1 port map( A => n116, B => memory_6_5_port, C => n111, D => 
                           memory_7_5_port, Y => n961);
   U1214 : NAND3X1 port map( A => n966, B => n967, C => n968, Y => n959);
   U1215 : NOR2X1 port map( A => n969, B => n970, Y => n968);
   U1216 : OAI22X1 port map( A => n750, B => n147, C => n758, D => n146, Y => 
                           n970);
   U1217 : OAI22X1 port map( A => n766, B => n135, C => n774, D => n136, Y => 
                           n969);
   U1218 : AOI22X1 port map( A => n113, B => memory_15_5_port, C => n109, D => 
                           memory_14_5_port, Y => n967);
   U1219 : AOI22X1 port map( A => n915, B => memory_13_5_port, C => n916, D => 
                           memory_12_5_port, Y => n966);
   U1220 : NAND2X1 port map( A => n972, B => n973, Y => n971);
   U1221 : NOR2X1 port map( A => n974, B => n975, Y => n973);
   U1222 : NAND3X1 port map( A => n976, B => n977, C => n978, Y => n975);
   U1223 : NOR2X1 port map( A => n979, B => n980, Y => n978);
   U1224 : OAI22X1 port map( A => n783, B => n141, C => n791, D => n140, Y => 
                           n980);
   U1225 : OAI22X1 port map( A => n799, B => n128, C => n807, D => n130, Y => 
                           n979);
   U1226 : AOI22X1 port map( A => n114, B => memory_23_4_port, C => n110, D => 
                           memory_22_4_port, Y => n977);
   U1227 : AOI22X1 port map( A => n840, B => memory_21_4_port, C => n841, D => 
                           memory_20_4_port, Y => n976);
   U1228 : NAND3X1 port map( A => n981, B => n982, C => n983, Y => n974);
   U1229 : NOR2X1 port map( A => n984, B => n985, Y => n983);
   U1230 : OAI22X1 port map( A => n709, B => n143, C => n701, D => n142, Y => 
                           n985);
   U1231 : OAI22X1 port map( A => n693, B => n131, C => n685, D => n132, Y => 
                           n984);
   U1232 : AOI22X1 port map( A => n115, B => memory_31_4_port, C => n112, D => 
                           memory_30_4_port, Y => n982);
   U1233 : AOI22X1 port map( A => n852, B => memory_29_4_port, C => n865, D => 
                           memory_28_4_port, Y => n981);
   U1234 : NOR2X1 port map( A => n986, B => n987, Y => n972);
   U1235 : NAND3X1 port map( A => n988, B => n989, C => n990, Y => n987);
   U1236 : NOR2X1 port map( A => n991, B => n992, Y => n990);
   U1237 : OAI22X1 port map( A => n742, B => n133, C => n734, D => n134, Y => 
                           n992);
   U1238 : OAI22X1 port map( A => n726, B => n145, C => n718, D => n144, Y => 
                           n991);
   U1239 : AOI22X1 port map( A => n908, B => memory_4_4_port, C => n909, D => 
                           memory_5_4_port, Y => n989);
   U1240 : AOI22X1 port map( A => n116, B => memory_6_4_port, C => n111, D => 
                           memory_7_4_port, Y => n988);
   U1241 : NAND3X1 port map( A => n993, B => n994, C => n995, Y => n986);
   U1242 : NOR2X1 port map( A => n996, B => n997, Y => n995);
   U1243 : OAI22X1 port map( A => n751, B => n147, C => n759, D => n146, Y => 
                           n997);
   U1244 : OAI22X1 port map( A => n767, B => n135, C => n775, D => n136, Y => 
                           n996);
   U1245 : AOI22X1 port map( A => n113, B => memory_15_4_port, C => n109, D => 
                           memory_14_4_port, Y => n994);
   U1246 : AOI22X1 port map( A => n915, B => memory_13_4_port, C => n916, D => 
                           memory_12_4_port, Y => n993);
   U1247 : NAND2X1 port map( A => n999, B => n1000, Y => n998);
   U1248 : NOR2X1 port map( A => n1001, B => n1002, Y => n1000);
   U1249 : NAND3X1 port map( A => n1003, B => n1004, C => n1005, Y => n1002);
   U1250 : NOR2X1 port map( A => n1006, B => n1007, Y => n1005);
   U1251 : OAI22X1 port map( A => n784, B => n141, C => n792, D => n140, Y => 
                           n1007);
   U1252 : OAI22X1 port map( A => n800, B => n128, C => n808, D => n130, Y => 
                           n1006);
   U1253 : AOI22X1 port map( A => n114, B => memory_23_3_port, C => n110, D => 
                           memory_22_3_port, Y => n1004);
   U1254 : AOI22X1 port map( A => n840, B => memory_21_3_port, C => n841, D => 
                           memory_20_3_port, Y => n1003);
   U1255 : NAND3X1 port map( A => n1008, B => n1009, C => n1010, Y => n1001);
   U1256 : NOR2X1 port map( A => n1011, B => n1012, Y => n1010);
   U1257 : OAI22X1 port map( A => n710, B => n143, C => n702, D => n142, Y => 
                           n1012);
   U1258 : OAI22X1 port map( A => n694, B => n131, C => n686, D => n132, Y => 
                           n1011);
   U1259 : AOI22X1 port map( A => n115, B => memory_31_3_port, C => n112, D => 
                           memory_30_3_port, Y => n1009);
   U1260 : AOI22X1 port map( A => n852, B => memory_29_3_port, C => n865, D => 
                           memory_28_3_port, Y => n1008);
   U1261 : NOR2X1 port map( A => n1013, B => n1014, Y => n999);
   U1262 : NAND3X1 port map( A => n1015, B => n1016, C => n1017, Y => n1014);
   U1263 : NOR2X1 port map( A => n1018, B => n1019, Y => n1017);
   U1264 : OAI22X1 port map( A => n741, B => n133, C => n733, D => n134, Y => 
                           n1019);
   U1265 : OAI22X1 port map( A => n725, B => n145, C => n717, D => n144, Y => 
                           n1018);
   U1266 : AOI22X1 port map( A => n908, B => memory_4_3_port, C => n909, D => 
                           memory_5_3_port, Y => n1016);
   U1267 : AOI22X1 port map( A => n116, B => memory_6_3_port, C => n111, D => 
                           memory_7_3_port, Y => n1015);
   U1268 : NAND3X1 port map( A => n1020, B => n1021, C => n1022, Y => n1013);
   U1269 : NOR2X1 port map( A => n1023, B => n1024, Y => n1022);
   U1270 : OAI22X1 port map( A => n752, B => n147, C => n760, D => n146, Y => 
                           n1024);
   U1271 : OAI22X1 port map( A => n768, B => n135, C => n776, D => n136, Y => 
                           n1023);
   U1272 : AOI22X1 port map( A => n113, B => memory_15_3_port, C => n109, D => 
                           memory_14_3_port, Y => n1021);
   U1273 : AOI22X1 port map( A => n915, B => memory_13_3_port, C => n916, D => 
                           memory_12_3_port, Y => n1020);
   U1274 : NAND2X1 port map( A => n1026, B => n1027, Y => n1025);
   U1275 : NOR2X1 port map( A => n1028, B => n1029, Y => n1027);
   U1276 : NAND3X1 port map( A => n1040, B => n1041, C => n1042, Y => n1029);
   U1277 : NOR2X1 port map( A => n1043, B => n1044, Y => n1042);
   U1278 : OAI22X1 port map( A => n785, B => n141, C => n793, D => n140, Y => 
                           n1044);
   U1279 : OAI22X1 port map( A => n801, B => n128, C => n809, D => n130, Y => 
                           n1043);
   U1280 : AOI22X1 port map( A => n114, B => memory_23_2_port, C => n110, D => 
                           memory_22_2_port, Y => n1041);
   U1281 : AOI22X1 port map( A => n840, B => memory_21_2_port, C => n841, D => 
                           memory_20_2_port, Y => n1040);
   U1282 : NAND3X1 port map( A => n1045, B => n1046, C => n1047, Y => n1028);
   U1283 : NOR2X1 port map( A => n1048, B => n1049, Y => n1047);
   U1284 : OAI22X1 port map( A => n711, B => n143, C => n703, D => n142, Y => 
                           n1049);
   U1285 : OAI22X1 port map( A => n695, B => n131, C => n687, D => n132, Y => 
                           n1048);
   U1286 : AOI22X1 port map( A => n115, B => memory_31_2_port, C => n112, D => 
                           memory_30_2_port, Y => n1046);
   U1287 : AOI22X1 port map( A => n852, B => memory_29_2_port, C => n865, D => 
                           memory_28_2_port, Y => n1045);
   U1288 : NOR2X1 port map( A => n1050, B => n1051, Y => n1026);
   U1289 : NAND3X1 port map( A => n1052, B => n1053, C => n1054, Y => n1051);
   U1290 : NOR2X1 port map( A => n1055, B => n1058, Y => n1054);
   U1291 : OAI22X1 port map( A => n740, B => n133, C => n732, D => n134, Y => 
                           n1058);
   U1292 : OAI22X1 port map( A => n724, B => n145, C => n716, D => n144, Y => 
                           n1055);
   U1293 : AOI22X1 port map( A => n908, B => memory_4_2_port, C => n909, D => 
                           memory_5_2_port, Y => n1053);
   U1294 : AOI22X1 port map( A => n116, B => memory_6_2_port, C => n111, D => 
                           memory_7_2_port, Y => n1052);
   U1295 : NAND3X1 port map( A => n1059, B => n1060, C => n1061, Y => n1050);
   U1296 : NOR2X1 port map( A => n1062, B => n1063, Y => n1061);
   U1297 : OAI22X1 port map( A => n753, B => n147, C => n761, D => n146, Y => 
                           n1063);
   U1298 : OAI22X1 port map( A => n769, B => n135, C => n777, D => n136, Y => 
                           n1062);
   U1299 : AOI22X1 port map( A => n113, B => memory_15_2_port, C => n109, D => 
                           memory_14_2_port, Y => n1060);
   U1300 : AOI22X1 port map( A => n915, B => memory_13_2_port, C => n916, D => 
                           memory_12_2_port, Y => n1059);
   U1301 : NAND2X1 port map( A => n1065, B => n1066, Y => n1064);
   U1302 : NOR2X1 port map( A => n1067, B => n1068, Y => n1066);
   U1303 : NAND3X1 port map( A => n1069, B => n1070, C => n1071, Y => n1068);
   U1304 : NOR2X1 port map( A => n1168, B => n1169, Y => n1071);
   U1305 : OAI22X1 port map( A => n786, B => n141, C => n794, D => n140, Y => 
                           n1169);
   U1306 : OAI22X1 port map( A => n802, B => n128, C => n810, D => n130, Y => 
                           n1168);
   U1307 : AOI22X1 port map( A => n114, B => memory_23_1_port, C => n110, D => 
                           memory_22_1_port, Y => n1070);
   U1308 : AOI22X1 port map( A => n840, B => memory_21_1_port, C => n841, D => 
                           memory_20_1_port, Y => n1069);
   U1309 : NAND3X1 port map( A => n1170, B => n1171, C => n1172, Y => n1067);
   U1310 : NOR2X1 port map( A => n1173, B => n1174, Y => n1172);
   U1311 : OAI22X1 port map( A => n712, B => n143, C => n704, D => n142, Y => 
                           n1174);
   U1312 : OAI22X1 port map( A => n696, B => n131, C => n688, D => n132, Y => 
                           n1173);
   U1313 : AOI22X1 port map( A => n115, B => memory_31_1_port, C => n112, D => 
                           memory_30_1_port, Y => n1171);
   U1314 : AOI22X1 port map( A => n852, B => memory_29_1_port, C => n865, D => 
                           memory_28_1_port, Y => n1170);
   U1315 : NOR2X1 port map( A => n1175, B => n1176, Y => n1065);
   U1316 : NAND3X1 port map( A => n1177, B => n1178, C => n1179, Y => n1176);
   U1317 : NOR2X1 port map( A => n1180, B => n1181, Y => n1179);
   U1318 : OAI22X1 port map( A => n739, B => n133, C => n731, D => n134, Y => 
                           n1181);
   U1319 : OAI22X1 port map( A => n723, B => n145, C => n715, D => n144, Y => 
                           n1180);
   U1320 : AOI22X1 port map( A => n908, B => memory_4_1_port, C => n909, D => 
                           memory_5_1_port, Y => n1178);
   U1321 : AOI22X1 port map( A => n116, B => memory_6_1_port, C => n111, D => 
                           memory_7_1_port, Y => n1177);
   U1322 : NAND3X1 port map( A => n1182, B => n1183, C => n1184, Y => n1175);
   U1323 : NOR2X1 port map( A => n1185, B => n1186, Y => n1184);
   U1324 : OAI22X1 port map( A => n754, B => n147, C => n762, D => n146, Y => 
                           n1186);
   U1325 : OAI22X1 port map( A => n770, B => n135, C => n778, D => n136, Y => 
                           n1185);
   U1326 : AOI22X1 port map( A => n113, B => memory_15_1_port, C => n109, D => 
                           memory_14_1_port, Y => n1183);
   U1327 : AOI22X1 port map( A => n915, B => memory_13_1_port, C => n916, D => 
                           memory_12_1_port, Y => n1182);
   U1328 : NAND2X1 port map( A => n1188, B => n1189, Y => n1187);
   U1329 : NOR2X1 port map( A => n1190, B => n1191, Y => n1189);
   U1330 : NAND3X1 port map( A => n1192, B => n1193, C => n1194, Y => n1191);
   U1331 : NOR2X1 port map( A => n1195, B => n1196, Y => n1194);
   U1332 : OAI22X1 port map( A => n787, B => n141, C => n795, D => n140, Y => 
                           n1196);
   U1333 : OAI22X1 port map( A => n803, B => n128, C => n811, D => n130, Y => 
                           n1195);
   U1334 : AOI22X1 port map( A => n114, B => memory_23_0_port, C => n110, D => 
                           memory_22_0_port, Y => n1193);
   U1335 : AOI22X1 port map( A => n840, B => memory_21_0_port, C => n841, D => 
                           memory_20_0_port, Y => n1192);
   U1336 : NAND3X1 port map( A => n1197, B => n1198, C => n1199, Y => n1190);
   U1337 : NOR2X1 port map( A => n1200, B => n1201, Y => n1199);
   U1338 : OAI22X1 port map( A => n713, B => n143, C => n705, D => n142, Y => 
                           n1201);
   U1339 : OAI22X1 port map( A => n697, B => n131, C => n689, D => n132, Y => 
                           n1200);
   U1340 : AOI22X1 port map( A => n115, B => memory_31_0_port, C => n112, D => 
                           memory_30_0_port, Y => n1198);
   U1341 : AOI22X1 port map( A => n852, B => memory_29_0_port, C => n865, D => 
                           memory_28_0_port, Y => n1197);
   U1342 : NOR2X1 port map( A => n1202, B => n1203, Y => n1188);
   U1343 : NAND3X1 port map( A => n1204, B => n1205, C => n1206, Y => n1203);
   U1344 : NOR2X1 port map( A => n1207, B => n1208, Y => n1206);
   U1345 : OAI22X1 port map( A => n738, B => n133, C => n730, D => n134, Y => 
                           n1208);
   U1346 : OAI22X1 port map( A => n722, B => n145, C => n714, D => n144, Y => 
                           n1207);
   U1347 : AOI22X1 port map( A => n908, B => memory_4_0_port, C => n909, D => 
                           memory_5_0_port, Y => n1205);
   U1348 : AOI22X1 port map( A => n116, B => memory_6_0_port, C => n111, D => 
                           memory_7_0_port, Y => n1204);
   U1349 : NAND3X1 port map( A => n1209, B => n1210, C => n1211, Y => n1202);
   U1350 : NOR2X1 port map( A => n1212, B => n1213, Y => n1211);
   U1351 : OAI22X1 port map( A => n755, B => n147, C => n763, D => n146, Y => 
                           n1213);
   U1352 : OAI22X1 port map( A => n771, B => n135, C => n779, D => n136, Y => 
                           n1212);
   U1353 : AOI22X1 port map( A => n113, B => memory_15_0_port, C => n109, D => 
                           memory_14_0_port, Y => n1210);
   U1354 : AOI22X1 port map( A => n915, B => memory_13_0_port, C => n916, D => 
                           memory_12_0_port, Y => n1209);
   U1355 : NAND2X1 port map( A => n1215, B => n1216, Y => n1214);
   U1356 : NOR2X1 port map( A => n1217, B => n1218, Y => n1216);
   U1357 : NAND3X1 port map( A => n1219, B => n1220, C => n1221, Y => n1218);
   U1358 : NOR2X1 port map( A => n1222, B => n1223, Y => n1221);
   U1359 : OAI22X1 port map( A => n820, B => n141, C => n822, D => n140, Y => 
                           n1223);
   U1360 : OAI22X1 port map( A => n824, B => n128, C => n826, D => n130, Y => 
                           n1222);
   U1361 : AOI22X1 port map( A => n114, B => opcode_23_1_port, C => n110, D => 
                           opcode_22_1_port, Y => n1220);
   U1362 : AOI22X1 port map( A => n840, B => opcode_21_1_port, C => n841, D => 
                           opcode_20_1_port, Y => n1219);
   U1363 : NAND3X1 port map( A => n1224, B => n1225, C => n1226, Y => n1217);
   U1364 : NOR2X1 port map( A => n1227, B => n1228, Y => n1226);
   U1365 : OAI22X1 port map( A => n672, B => n143, C => n670, D => n142, Y => 
                           n1228);
   U1366 : OAI22X1 port map( A => n668, B => n131, C => n666, D => n132, Y => 
                           n1227);
   U1367 : AOI22X1 port map( A => n115, B => opcode_31_1_port, C => n112, D => 
                           opcode_30_1_port, Y => n1225);
   U1368 : AOI22X1 port map( A => n852, B => opcode_29_1_port, C => n865, D => 
                           opcode_28_1_port, Y => n1224);
   U1369 : NOR2X1 port map( A => n1229, B => n1230, Y => n1215);
   U1370 : NAND3X1 port map( A => n1231, B => n1232, C => n1233, Y => n1230);
   U1371 : NOR2X1 port map( A => n1234, B => n1235, Y => n1233);
   U1372 : OAI22X1 port map( A => n681, B => n133, C => n679, D => n134, Y => 
                           n1235);
   U1373 : OAI22X1 port map( A => n677, B => n145, C => n675, D => n144, Y => 
                           n1234);
   U1374 : AOI22X1 port map( A => n908, B => opcode_4_1_port, C => n909, D => 
                           opcode_5_1_port, Y => n1232);
   U1375 : AOI22X1 port map( A => n116, B => opcode_6_1_port, C => n111, D => 
                           opcode_7_1_port, Y => n1231);
   U1376 : NAND3X1 port map( A => n1236, B => n1237, C => n1238, Y => n1229);
   U1377 : NOR2X1 port map( A => n1239, B => n1240, Y => n1238);
   U1378 : OAI22X1 port map( A => n812, B => n147, C => n814, D => n146, Y => 
                           n1240);
   U1379 : OAI22X1 port map( A => n816, B => n135, C => n818, D => n136, Y => 
                           n1239);
   U1380 : AOI22X1 port map( A => n113, B => opcode_15_1_port, C => n109, D => 
                           opcode_14_1_port, Y => n1237);
   U1381 : AOI22X1 port map( A => n915, B => opcode_13_1_port, C => n916, D => 
                           opcode_12_1_port, Y => n1236);
   U1382 : NAND2X1 port map( A => n1242, B => n1243, Y => n1241);
   U1383 : NOR2X1 port map( A => n1244, B => n1245, Y => n1243);
   U1384 : NAND3X1 port map( A => n1246, B => n1247, C => n1248, Y => n1245);
   U1385 : NOR2X1 port map( A => n1249, B => n1250, Y => n1248);
   U1386 : OAI22X1 port map( A => n821, B => n141, C => n823, D => n140, Y => 
                           n1250);
   U1387 : NAND2X1 port map( A => n1251, B => n1252, Y => n838);
   U1388 : OAI22X1 port map( A => n825, B => n128, C => n827, D => n130, Y => 
                           n1249);
   U1389 : AOI22X1 port map( A => n114, B => opcode_23_0_port, C => n110, D => 
                           opcode_22_0_port, Y => n1247);
   U1390 : AOI22X1 port map( A => n840, B => opcode_21_0_port, C => n841, D => 
                           opcode_20_0_port, Y => n1246);
   U1391 : INVX1 port map( A => n1255, Y => n1253);
   U1392 : NAND3X1 port map( A => n662, B => n664, C => n84, Y => n1255);
   U1393 : INVX1 port map( A => n1256, Y => n1251);
   U1394 : NAND3X1 port map( A => n76, B => n664, C => n84, Y => n1256);
   U1395 : NAND3X1 port map( A => n1257, B => n1258, C => n1259, Y => n1244);
   U1396 : NOR2X1 port map( A => n1260, B => n1261, Y => n1259);
   U1397 : OAI22X1 port map( A => n673, B => n143, C => n671, D => n142, Y => 
                           n1261);
   U1398 : OAI22X1 port map( A => n669, B => n131, C => n667, D => n132, Y => 
                           n1260);
   U1399 : AOI22X1 port map( A => n115, B => opcode_31_0_port, C => n112, D => 
                           opcode_30_0_port, Y => n1258);
   U1400 : AOI22X1 port map( A => n852, B => opcode_29_0_port, C => n865, D => 
                           opcode_28_0_port, Y => n1257);
   U1401 : INVX1 port map( A => n1264, Y => n1263);
   U1402 : NAND3X1 port map( A => n153, B => n662, C => n84, Y => n1264);
   U1403 : INVX1 port map( A => n1265, Y => n1262);
   U1404 : NAND3X1 port map( A => n153, B => n76, C => n84, Y => n1265);
   U1405 : NOR2X1 port map( A => n1266, B => n1267, Y => n1242);
   U1406 : NAND3X1 port map( A => n1268, B => n1269, C => n1270, Y => n1267);
   U1407 : NOR2X1 port map( A => n1271, B => n1272, Y => n1270);
   U1408 : OAI22X1 port map( A => n680, B => n133, C => n678, D => n134, Y => 
                           n1272);
   U1409 : OAI22X1 port map( A => n676, B => n145, C => n674, D => n144, Y => 
                           n1271);
   U1410 : AOI22X1 port map( A => n908, B => opcode_4_0_port, C => n909, D => 
                           opcode_5_0_port, Y => n1269);
   U1411 : AOI22X1 port map( A => n116, B => opcode_6_0_port, C => n111, D => 
                           opcode_7_0_port, Y => n1268);
   U1412 : INVX1 port map( A => n1275, Y => n1274);
   U1413 : NAND3X1 port map( A => n664, B => n665, C => n76, Y => n1275);
   U1414 : INVX1 port map( A => n1276, Y => n1273);
   U1415 : NAND3X1 port map( A => n664, B => n665, C => n662, Y => n1276);
   U1416 : NAND3X1 port map( A => n1277, B => n1278, C => n1279, Y => n1266);
   U1417 : NOR2X1 port map( A => n1280, B => n1281, Y => n1279);
   U1418 : OAI22X1 port map( A => n813, B => n147, C => n815, D => n146, Y => 
                           n1281);
   U1419 : NOR2X1 port map( A => n51, B => readptr_2_port, Y => n1252);
   U1420 : OAI22X1 port map( A => n817, B => n135, C => n819, D => n136, Y => 
                           n1280);
   U1421 : AOI22X1 port map( A => n113, B => opcode_15_0_port, C => n109, D => 
                           opcode_14_0_port, Y => n1278);
   U1422 : AOI22X1 port map( A => n915, B => opcode_13_0_port, C => n916, D => 
                           opcode_12_0_port, Y => n1277);
   U1423 : INVX1 port map( A => n1284, Y => n1283);
   U1424 : NAND3X1 port map( A => n662, B => n665, C => n153, Y => n1284);
   U1425 : NOR2X1 port map( A => n663, B => n51, Y => n1254);
   U1426 : INVX1 port map( A => n1285, Y => n1282);
   U1427 : NAND3X1 port map( A => n76, B => n665, C => n153, Y => n1285);

end SYN_BRFIFO;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RBUFFER_1 is

   port( CLK, RST, NEXT_BYTE : in std_logic;  DATA : in std_logic_vector (7 
         downto 0);  OPCODE : in std_logic_vector (1 downto 0);  BYTE_COUNT : 
         in std_logic_vector (4 downto 0);  EOP : in std_logic;  B_READY, 
         R_ENABLE : out std_logic;  PRGA_IN : out std_logic_vector (7 downto 0)
         ;  PRGA_OPCODE : out std_logic_vector (1 downto 0));

end RBUFFER_1;

architecture SYN_brbuffer of RBUFFER_1 is

   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal B_READY_port, R_ENABLE_port, PRGA_IN_7_port, PRGA_IN_6_port, 
      PRGA_IN_5_port, PRGA_IN_4_port, PRGA_IN_3_port, PRGA_IN_2_port, 
      PRGA_IN_1_port, PRGA_IN_0_port, PRGA_OPCODE_1_port, PRGA_OPCODE_0_port, 
      state_2_port, state_1_port, state_0_port, nextState_2_port, 
      nextState_1_port, nextState_0_port, tempData_7_port, tempData_6_port, 
      tempData_5_port, tempData_4_port, tempData_3_port, tempData_2_port, 
      tempData_1_port, tempData_0_port, tempOpcode_1_port, tempOpcode_0_port, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n97, n98, n99, 
      n100, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n86, n88 : std_logic;

begin
   B_READY <= B_READY_port;
   R_ENABLE <= R_ENABLE_port;
   PRGA_IN <= ( PRGA_IN_7_port, PRGA_IN_6_port, PRGA_IN_5_port, PRGA_IN_4_port,
      PRGA_IN_3_port, PRGA_IN_2_port, PRGA_IN_1_port, PRGA_IN_0_port );
   PRGA_OPCODE <= ( PRGA_OPCODE_1_port, PRGA_OPCODE_0_port );
   
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n1, S => n100, Q => state_0_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n1, S => n99, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n1, S => n98, Q => state_1_port);
   B_READY_reg : DFFPOSX1 port map( D => n97, CLK => CLK, Q => B_READY_port);
   tempData_reg_7_inst : DFFPOSX1 port map( D => n68, CLK => CLK, Q => 
                           tempData_7_port);
   tempData_reg_6_inst : DFFPOSX1 port map( D => n69, CLK => CLK, Q => 
                           tempData_6_port);
   tempData_reg_5_inst : DFFPOSX1 port map( D => n70, CLK => CLK, Q => 
                           tempData_5_port);
   tempData_reg_4_inst : DFFPOSX1 port map( D => n71, CLK => CLK, Q => 
                           tempData_4_port);
   tempData_reg_3_inst : DFFPOSX1 port map( D => n72, CLK => CLK, Q => 
                           tempData_3_port);
   tempData_reg_2_inst : DFFPOSX1 port map( D => n73, CLK => CLK, Q => 
                           tempData_2_port);
   tempData_reg_1_inst : DFFPOSX1 port map( D => n74, CLK => CLK, Q => 
                           tempData_1_port);
   tempData_reg_0_inst : DFFPOSX1 port map( D => n75, CLK => CLK, Q => 
                           tempData_0_port);
   tempOpcode_reg_1_inst : DFFPOSX1 port map( D => n86, CLK => CLK, Q => 
                           tempOpcode_1_port);
   PRGA_OPCODE_reg_1_inst : DFFPOSX1 port map( D => n87, CLK => CLK, Q => 
                           PRGA_OPCODE_1_port);
   tempOpcode_reg_0_inst : DFFPOSX1 port map( D => n88, CLK => CLK, Q => 
                           tempOpcode_0_port);
   PRGA_OPCODE_reg_0_inst : DFFPOSX1 port map( D => n85, CLK => CLK, Q => 
                           PRGA_OPCODE_0_port);
   R_ENABLE_reg : DFFPOSX1 port map( D => n84, CLK => CLK, Q => R_ENABLE_port);
   PRGA_IN_reg_7_inst : DFFPOSX1 port map( D => n83, CLK => CLK, Q => 
                           PRGA_IN_7_port);
   PRGA_IN_reg_6_inst : DFFPOSX1 port map( D => n82, CLK => CLK, Q => 
                           PRGA_IN_6_port);
   PRGA_IN_reg_5_inst : DFFPOSX1 port map( D => n81, CLK => CLK, Q => 
                           PRGA_IN_5_port);
   PRGA_IN_reg_4_inst : DFFPOSX1 port map( D => n80, CLK => CLK, Q => 
                           PRGA_IN_4_port);
   PRGA_IN_reg_3_inst : DFFPOSX1 port map( D => n79, CLK => CLK, Q => 
                           PRGA_IN_3_port);
   PRGA_IN_reg_2_inst : DFFPOSX1 port map( D => n78, CLK => CLK, Q => 
                           PRGA_IN_2_port);
   PRGA_IN_reg_1_inst : DFFPOSX1 port map( D => n77, CLK => CLK, Q => 
                           PRGA_IN_1_port);
   PRGA_IN_reg_0_inst : DFFPOSX1 port map( D => n76, CLK => CLK, Q => 
                           PRGA_IN_0_port);
   n98 <= '1';
   n99 <= '1';
   n100 <= '1';
   U3 : INVX2 port map( A => n41, Y => n28);
   U4 : INVX2 port map( A => RST, Y => n1);
   U5 : OR2X2 port map( A => n39, B => RST, Y => n29);
   U6 : AND2X2 port map( A => n39, B => n1, Y => n44);
   U7 : OAI21X1 port map( A => n2, B => n3, C => n4, Y => nextState_2_port);
   U8 : MUX2X1 port map( B => n5, A => n6, S => state_0_port, Y => n4);
   U9 : NOR2X1 port map( A => state_2_port, B => n7, Y => n6);
   U10 : AND2X1 port map( A => state_2_port, B => n8, Y => n5);
   U11 : OAI21X1 port map( A => NEXT_BYTE, B => n9, C => state_1_port, Y => n8)
                           ;
   U12 : AND2X1 port map( A => n10, B => NEXT_BYTE, Y => n2);
   U13 : OAI21X1 port map( A => state_2_port, B => n11, C => n12, Y => 
                           nextState_1_port);
   U14 : OAI21X1 port map( A => n13, B => n14, C => n15, Y => n12);
   U15 : INVX1 port map( A => n3, Y => n14);
   U16 : OAI21X1 port map( A => state_2_port, B => n16, C => n17, Y => 
                           nextState_0_port);
   U17 : AOI22X1 port map( A => n18, B => n19, C => NEXT_BYTE, D => n20, Y => 
                           n17);
   U18 : OAI21X1 port map( A => n10, B => n3, C => n21, Y => n20);
   U19 : INVX1 port map( A => n13, Y => n21);
   U20 : NOR2X1 port map( A => n16, B => n9, Y => n13);
   U21 : NOR2X1 port map( A => n22, B => BYTE_COUNT(4), Y => n9);
   U22 : NAND3X1 port map( A => state_0_port, B => n7, C => state_2_port, Y => 
                           n3);
   U23 : AND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n10);
   U24 : OAI21X1 port map( A => n23, B => n15, C => n24, Y => n19);
   U25 : INVX1 port map( A => NEXT_BYTE, Y => n15);
   U26 : AOI21X1 port map( A => EOP, B => n22, C => BYTE_COUNT(4), Y => n23);
   U27 : NAND2X1 port map( A => n25, B => n26, Y => n22);
   U28 : NOR2X1 port map( A => BYTE_COUNT(3), B => BYTE_COUNT(2), Y => n26);
   U29 : NOR2X1 port map( A => BYTE_COUNT(1), B => BYTE_COUNT(0), Y => n25);
   U30 : NOR2X1 port map( A => state_1_port, B => state_0_port, Y => n18);
   U31 : INVX1 port map( A => n27, Y => n68);
   U32 : AOI22X1 port map( A => n28, B => DATA(7), C => n29, D => 
                           tempData_7_port, Y => n27);
   U33 : INVX1 port map( A => n30, Y => n69);
   U34 : AOI22X1 port map( A => n28, B => DATA(6), C => n29, D => 
                           tempData_6_port, Y => n30);
   U35 : INVX1 port map( A => n31, Y => n70);
   U36 : AOI22X1 port map( A => n28, B => DATA(5), C => n29, D => 
                           tempData_5_port, Y => n31);
   U37 : INVX1 port map( A => n32, Y => n71);
   U38 : AOI22X1 port map( A => n28, B => DATA(4), C => n29, D => 
                           tempData_4_port, Y => n32);
   U39 : INVX1 port map( A => n33, Y => n72);
   U40 : AOI22X1 port map( A => n28, B => DATA(3), C => n29, D => 
                           tempData_3_port, Y => n33);
   U41 : INVX1 port map( A => n34, Y => n73);
   U42 : AOI22X1 port map( A => n28, B => DATA(2), C => n29, D => 
                           tempData_2_port, Y => n34);
   U43 : INVX1 port map( A => n35, Y => n74);
   U44 : AOI22X1 port map( A => n28, B => DATA(1), C => n29, D => 
                           tempData_1_port, Y => n35);
   U45 : INVX1 port map( A => n36, Y => n75);
   U46 : AOI22X1 port map( A => n28, B => DATA(0), C => n29, D => 
                           tempData_0_port, Y => n36);
   U47 : INVX1 port map( A => n37, Y => n86);
   U48 : AOI22X1 port map( A => OPCODE(1), B => n28, C => n29, D => 
                           tempOpcode_1_port, Y => n37);
   U49 : INVX1 port map( A => n38, Y => n88);
   U50 : AOI22X1 port map( A => OPCODE(0), B => n28, C => n29, D => 
                           tempOpcode_0_port, Y => n38);
   U51 : OAI21X1 port map( A => n1, B => n40, C => n41, Y => n97);
   U52 : INVX1 port map( A => B_READY_port, Y => n40);
   U53 : OAI21X1 port map( A => n1, B => n42, C => n43, Y => n87);
   U54 : AOI22X1 port map( A => n28, B => OPCODE(1), C => n44, D => 
                           tempOpcode_1_port, Y => n43);
   U55 : INVX1 port map( A => PRGA_OPCODE_1_port, Y => n42);
   U56 : OAI21X1 port map( A => n1, B => n45, C => n46, Y => n85);
   U57 : AOI22X1 port map( A => n28, B => OPCODE(0), C => n44, D => 
                           tempOpcode_0_port, Y => n46);
   U58 : INVX1 port map( A => PRGA_OPCODE_0_port, Y => n45);
   U59 : MUX2X1 port map( B => n47, A => n48, S => RST, Y => n84);
   U60 : INVX1 port map( A => R_ENABLE_port, Y => n48);
   U61 : NAND3X1 port map( A => n7, B => n24, C => state_0_port, Y => n47);
   U62 : OAI21X1 port map( A => n1, B => n49, C => n50, Y => n83);
   U63 : AOI22X1 port map( A => DATA(7), B => n28, C => n44, D => 
                           tempData_7_port, Y => n50);
   U64 : INVX1 port map( A => PRGA_IN_7_port, Y => n49);
   U65 : OAI21X1 port map( A => n1, B => n51, C => n52, Y => n82);
   U66 : AOI22X1 port map( A => DATA(6), B => n28, C => n44, D => 
                           tempData_6_port, Y => n52);
   U67 : INVX1 port map( A => PRGA_IN_6_port, Y => n51);
   U68 : OAI21X1 port map( A => n1, B => n53, C => n54, Y => n81);
   U69 : AOI22X1 port map( A => DATA(5), B => n28, C => n44, D => 
                           tempData_5_port, Y => n54);
   U70 : INVX1 port map( A => PRGA_IN_5_port, Y => n53);
   U71 : OAI21X1 port map( A => n1, B => n55, C => n56, Y => n80);
   U72 : AOI22X1 port map( A => DATA(4), B => n28, C => n44, D => 
                           tempData_4_port, Y => n56);
   U73 : INVX1 port map( A => PRGA_IN_4_port, Y => n55);
   U74 : OAI21X1 port map( A => n1, B => n57, C => n58, Y => n79);
   U75 : AOI22X1 port map( A => DATA(3), B => n28, C => n44, D => 
                           tempData_3_port, Y => n58);
   U76 : INVX1 port map( A => PRGA_IN_3_port, Y => n57);
   U77 : OAI21X1 port map( A => n1, B => n59, C => n60, Y => n78);
   U78 : AOI22X1 port map( A => DATA(2), B => n28, C => n44, D => 
                           tempData_2_port, Y => n60);
   U79 : INVX1 port map( A => PRGA_IN_2_port, Y => n59);
   U80 : OAI21X1 port map( A => n1, B => n61, C => n62, Y => n77);
   U81 : AOI22X1 port map( A => DATA(1), B => n28, C => n44, D => 
                           tempData_1_port, Y => n62);
   U82 : INVX1 port map( A => PRGA_IN_1_port, Y => n61);
   U83 : OAI21X1 port map( A => n1, B => n63, C => n64, Y => n76);
   U84 : AOI22X1 port map( A => DATA(0), B => n28, C => n44, D => 
                           tempData_0_port, Y => n64);
   U85 : NAND2X1 port map( A => n11, B => state_2_port, Y => n39);
   U86 : INVX1 port map( A => n65, Y => n11);
   U87 : OAI21X1 port map( A => state_1_port, B => n66, C => n16, Y => n65);
   U88 : NAND2X1 port map( A => state_1_port, B => n66, Y => n16);
   U89 : NAND3X1 port map( A => n66, B => n7, C => n67, Y => n41);
   U90 : NOR2X1 port map( A => RST, B => n24, Y => n67);
   U91 : INVX1 port map( A => state_2_port, Y => n24);
   U92 : INVX1 port map( A => state_1_port, Y => n7);
   U93 : INVX1 port map( A => state_0_port, Y => n66);
   U94 : INVX1 port map( A => PRGA_IN_0_port, Y => n63);

end SYN_brbuffer;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_block_1 is

   port( CLK, RST, SERIAL_IN : in std_logic;  KEY_ERROR, PROG_ERROR : out 
         std_logic;  PLAINKEY : out std_logic_vector (63 downto 0);  RBUF_FULL,
         PARITY_ERROR : out std_logic);

end uart_rcv_block_1;

architecture SYN_struct1 of uart_rcv_block_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component uart_timer_1
      port( CLK, RST, TIMER_TRIG : in std_logic;  STOP_RCVING, SHIFT_STROBE : 
            out std_logic);
   end component;
   
   component keyreg_1
      port( CLK, RST, SBE, OE, RBUF_FULL : in std_logic;  RCV_DATA : in 
            std_logic_vector (7 downto 0);  PLAINKEY : out std_logic_vector (63
            downto 0);  KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR : out 
            std_logic);
   end component;
   
   component uart_sr_10bit_1
      port( CLK, RST, SHIFT_STROBE, SERIAL_IN : in std_logic;  LOAD_DATA : out 
            std_logic_vector (7 downto 0);  STOP_DATA : out std_logic_vector (1
            downto 0));
   end component;
   
   component uart_sb_check_1
      port( RST, CLK, SBC_CLR, SBC_EN : in std_logic;  STOP_DATA : in 
            std_logic_vector (1 downto 0);  SB_DETECT, SBE : out std_logic);
   end component;
   
   component uart_rcv_buf_full_1
      port( CLK, RST, CLR_RBUF, SET_RBUF_FULL : in std_logic;  RBUF_FULL : out 
            std_logic);
   end component;
   
   component uart_rcv_buf_1
      port( CLK, RST, LOAD_RBUF : in std_logic;  LOAD_DATA : in 
            std_logic_vector (7 downto 0);  RCV_DATA : out std_logic_vector (7 
            downto 0));
   end component;
   
   component uart_rcu_1
      port( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT : in std_logic;  
            RBUF_LOAD, TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR : 
            out std_logic);
   end component;
   
   component uart_error_1
      port( RST, CLK, RBUF_FULL, CHK_ERROR : in std_logic;  OE : out std_logic
            );
   end component;
   
   component uart_edge_detector_1
      port( CLK, RST, SERIAL_IN : in std_logic;  START_BIT : out std_logic);
   end component;
   
   signal RBUF_FULL_port, START_BIT, CHK_ERROR, OE, SB_DETECT, STOP_RCVING, 
      RBUF_LOAD, SBC_CLR, SBC_EN, SET_RBUF_FULL, TIMER_TRIG, LOAD_DATA_7_port, 
      LOAD_DATA_6_port, LOAD_DATA_5_port, LOAD_DATA_4_port, LOAD_DATA_3_port, 
      LOAD_DATA_2_port, LOAD_DATA_1_port, LOAD_DATA_0_port, RCV_DATA_7_port, 
      RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, RCV_DATA_3_port, 
      RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, CLR_RBUF, 
      STOP_DATA_1_port, STOP_DATA_0_port, SBE, SHIFT_STROBE, n1, n2 : std_logic
      ;

begin
   RBUF_FULL <= RBUF_FULL_port;
   
   U_0 : uart_edge_detector_1 port map( CLK => CLK, RST => n1, SERIAL_IN => 
                           SERIAL_IN, START_BIT => START_BIT);
   U_1 : uart_error_1 port map( RST => n1, CLK => CLK, RBUF_FULL => 
                           RBUF_FULL_port, CHK_ERROR => CHK_ERROR, OE => OE);
   U_2 : uart_rcu_1 port map( CLK => CLK, RST => n1, START_BIT => START_BIT, 
                           STOP_RCVING => STOP_RCVING, SB_DETECT => SB_DETECT, 
                           RBUF_LOAD => RBUF_LOAD, TIMER_TRIG => TIMER_TRIG, 
                           CHK_ERROR => CHK_ERROR, SET_RBUF_FULL => 
                           SET_RBUF_FULL, SBC_EN => SBC_EN, SBC_CLR => SBC_CLR)
                           ;
   U_3 : uart_rcv_buf_1 port map( CLK => CLK, RST => n1, LOAD_RBUF => RBUF_LOAD
                           , LOAD_DATA(7) => LOAD_DATA_7_port, LOAD_DATA(6) => 
                           LOAD_DATA_6_port, LOAD_DATA(5) => LOAD_DATA_5_port, 
                           LOAD_DATA(4) => LOAD_DATA_4_port, LOAD_DATA(3) => 
                           LOAD_DATA_3_port, LOAD_DATA(2) => LOAD_DATA_2_port, 
                           LOAD_DATA(1) => LOAD_DATA_1_port, LOAD_DATA(0) => 
                           LOAD_DATA_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port);
   U_4 : uart_rcv_buf_full_1 port map( CLK => CLK, RST => n1, CLR_RBUF => 
                           CLR_RBUF, SET_RBUF_FULL => SET_RBUF_FULL, RBUF_FULL 
                           => RBUF_FULL_port);
   U_5 : uart_sb_check_1 port map( RST => n1, CLK => CLK, SBC_CLR => SBC_CLR, 
                           SBC_EN => SBC_EN, STOP_DATA(1) => STOP_DATA_1_port, 
                           STOP_DATA(0) => STOP_DATA_0_port, SB_DETECT => 
                           SB_DETECT, SBE => SBE);
   U_6 : uart_sr_10bit_1 port map( CLK => CLK, RST => n1, SHIFT_STROBE => 
                           SHIFT_STROBE, SERIAL_IN => SERIAL_IN, LOAD_DATA(7) 
                           => LOAD_DATA_7_port, LOAD_DATA(6) => 
                           LOAD_DATA_6_port, LOAD_DATA(5) => LOAD_DATA_5_port, 
                           LOAD_DATA(4) => LOAD_DATA_4_port, LOAD_DATA(3) => 
                           LOAD_DATA_3_port, LOAD_DATA(2) => LOAD_DATA_2_port, 
                           LOAD_DATA(1) => LOAD_DATA_1_port, LOAD_DATA(0) => 
                           LOAD_DATA_0_port, STOP_DATA(1) => STOP_DATA_1_port, 
                           STOP_DATA(0) => STOP_DATA_0_port);
   U_8 : keyreg_1 port map( CLK => CLK, RST => n1, SBE => SBE, OE => OE, 
                           RBUF_FULL => RBUF_FULL_port, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           PLAINKEY(63) => PLAINKEY(63), PLAINKEY(62) => 
                           PLAINKEY(62), PLAINKEY(61) => PLAINKEY(61), 
                           PLAINKEY(60) => PLAINKEY(60), PLAINKEY(59) => 
                           PLAINKEY(59), PLAINKEY(58) => PLAINKEY(58), 
                           PLAINKEY(57) => PLAINKEY(57), PLAINKEY(56) => 
                           PLAINKEY(56), PLAINKEY(55) => PLAINKEY(55), 
                           PLAINKEY(54) => PLAINKEY(54), PLAINKEY(53) => 
                           PLAINKEY(53), PLAINKEY(52) => PLAINKEY(52), 
                           PLAINKEY(51) => PLAINKEY(51), PLAINKEY(50) => 
                           PLAINKEY(50), PLAINKEY(49) => PLAINKEY(49), 
                           PLAINKEY(48) => PLAINKEY(48), PLAINKEY(47) => 
                           PLAINKEY(47), PLAINKEY(46) => PLAINKEY(46), 
                           PLAINKEY(45) => PLAINKEY(45), PLAINKEY(44) => 
                           PLAINKEY(44), PLAINKEY(43) => PLAINKEY(43), 
                           PLAINKEY(42) => PLAINKEY(42), PLAINKEY(41) => 
                           PLAINKEY(41), PLAINKEY(40) => PLAINKEY(40), 
                           PLAINKEY(39) => PLAINKEY(39), PLAINKEY(38) => 
                           PLAINKEY(38), PLAINKEY(37) => PLAINKEY(37), 
                           PLAINKEY(36) => PLAINKEY(36), PLAINKEY(35) => 
                           PLAINKEY(35), PLAINKEY(34) => PLAINKEY(34), 
                           PLAINKEY(33) => PLAINKEY(33), PLAINKEY(32) => 
                           PLAINKEY(32), PLAINKEY(31) => PLAINKEY(31), 
                           PLAINKEY(30) => PLAINKEY(30), PLAINKEY(29) => 
                           PLAINKEY(29), PLAINKEY(28) => PLAINKEY(28), 
                           PLAINKEY(27) => PLAINKEY(27), PLAINKEY(26) => 
                           PLAINKEY(26), PLAINKEY(25) => PLAINKEY(25), 
                           PLAINKEY(24) => PLAINKEY(24), PLAINKEY(23) => 
                           PLAINKEY(23), PLAINKEY(22) => PLAINKEY(22), 
                           PLAINKEY(21) => PLAINKEY(21), PLAINKEY(20) => 
                           PLAINKEY(20), PLAINKEY(19) => PLAINKEY(19), 
                           PLAINKEY(18) => PLAINKEY(18), PLAINKEY(17) => 
                           PLAINKEY(17), PLAINKEY(16) => PLAINKEY(16), 
                           PLAINKEY(15) => PLAINKEY(15), PLAINKEY(14) => 
                           PLAINKEY(14), PLAINKEY(13) => PLAINKEY(13), 
                           PLAINKEY(12) => PLAINKEY(12), PLAINKEY(11) => 
                           PLAINKEY(11), PLAINKEY(10) => PLAINKEY(10), 
                           PLAINKEY(9) => PLAINKEY(9), PLAINKEY(8) => 
                           PLAINKEY(8), PLAINKEY(7) => PLAINKEY(7), PLAINKEY(6)
                           => PLAINKEY(6), PLAINKEY(5) => PLAINKEY(5), 
                           PLAINKEY(4) => PLAINKEY(4), PLAINKEY(3) => 
                           PLAINKEY(3), PLAINKEY(2) => PLAINKEY(2), PLAINKEY(1)
                           => PLAINKEY(1), PLAINKEY(0) => PLAINKEY(0), 
                           KEY_ERROR => KEY_ERROR, PROG_ERROR => PROG_ERROR, 
                           CLR_RBUFF => CLR_RBUF, PARITY_ERROR => PARITY_ERROR)
                           ;
   U_7 : uart_timer_1 port map( CLK => CLK, RST => n1, TIMER_TRIG => TIMER_TRIG
                           , STOP_RCVING => STOP_RCVING, SHIFT_STROBE => 
                           SHIFT_STROBE);
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct1;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1 is

   port( KEY : in std_logic_vector (63 downto 0);  CLK, RST, KEY_ERROR, 
         BYTE_READY : in std_logic;  BYTE : in std_logic_vector (7 downto 0);  
         OPCODE : in std_logic_vector (1 downto 0);  DATA_IN : in 
         std_logic_vector (7 downto 0);  PROCESSED_DATA : out std_logic_vector 
         (7 downto 0);  PDATA_READY, W_ENABLE, R_ENABLE : out std_logic;  ADDR,
         DATA : out std_logic_vector (7 downto 0));

end KSA_1;

architecture SYN_bksa of KSA_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUFX1
      port( A, EN : in std_logic;  Y : out std_logic);
   end component;
   
   component TBUFX2
      port( A, EN : in std_logic;  Y : out std_logic);
   end component;
   
   component KSA_1_DW01_inc_3
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_1_DW01_add_9
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_1_DW01_add_8
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_1_DW01_add_7
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_1_DW01_add_6
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_1_DW01_inc_1
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_1_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, PROCESSED_DATA_5_port, 
      PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, PROCESSED_DATA_2_port, 
      PROCESSED_DATA_1_port, PROCESSED_DATA_0_port, W_ENABLE_port, 
      R_ENABLE_port, ADDR_7_port, ADDR_6_port, ADDR_5_port, ADDR_4_port, 
      ADDR_3_port, ADDR_2_port, ADDR_1_port, ADDR_0_port, DATA_7_port, 
      DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, DATA_2_port, 
      DATA_1_port, DATA_0_port, state_4_port, state_3_port, state_2_port, 
      state_1_port, state_0_port, si_7_port, si_6_port, si_5_port, si_4_port, 
      si_3_port, si_2_port, si_1_port, si_0_port, sj_7_port, sj_6_port, 
      sj_5_port, sj_4_port, sj_3_port, sj_2_port, sj_1_port, sj_0_port, 
      currentProcessedData_7_port, currentProcessedData_6_port, 
      currentProcessedData_5_port, currentProcessedData_4_port, 
      currentProcessedData_3_port, currentProcessedData_2_port, 
      currentProcessedData_1_port, currentProcessedData_0_port, 
      nextState_4_port, nextState_3_port, nextState_2_port, nextState_1_port, 
      nextState_0_port, inti_7_port, inti_6_port, inti_5_port, inti_4_port, 
      inti_3_port, inti_2_port, inti_1_port, inti_0_port, intj_7_port, 
      intj_6_port, intj_5_port, intj_4_port, intj_3_port, intj_2_port, 
      intj_1_port, intj_0_port, keyi_2_port, keyi_1_port, keyi_0_port, 
      permuteComplete, temp_7_port, temp_6_port, temp_5_port, temp_4_port, 
      temp_3_port, temp_2_port, temp_1_port, temp_0_port, extratemp_7_port, 
      extratemp_6_port, extratemp_5_port, extratemp_4_port, extratemp_3_port, 
      extratemp_2_port, extratemp_1_port, extratemp_0_port, 
      nextProcessedData_7_port, nextProcessedData_6_port, 
      nextProcessedData_5_port, nextProcessedData_4_port, 
      nextProcessedData_3_port, nextProcessedData_2_port, 
      nextProcessedData_1_port, nextProcessedData_0_port, keyTable_0_7_port, 
      keyTable_0_6_port, keyTable_0_5_port, keyTable_0_4_port, 
      keyTable_0_3_port, keyTable_0_2_port, keyTable_0_1_port, 
      keyTable_0_0_port, keyTable_1_7_port, keyTable_1_6_port, 
      keyTable_1_5_port, keyTable_1_4_port, keyTable_1_3_port, 
      keyTable_1_2_port, keyTable_1_1_port, keyTable_1_0_port, 
      keyTable_2_7_port, keyTable_2_6_port, keyTable_2_5_port, 
      keyTable_2_4_port, keyTable_2_3_port, keyTable_2_2_port, 
      keyTable_2_1_port, keyTable_2_0_port, keyTable_3_7_port, 
      keyTable_3_6_port, keyTable_3_5_port, keyTable_3_4_port, 
      keyTable_3_3_port, keyTable_3_2_port, keyTable_3_1_port, 
      keyTable_3_0_port, keyTable_4_7_port, keyTable_4_6_port, 
      keyTable_4_5_port, keyTable_4_4_port, keyTable_4_3_port, 
      keyTable_4_2_port, keyTable_4_1_port, keyTable_4_0_port, 
      keyTable_5_7_port, keyTable_5_6_port, keyTable_5_5_port, 
      keyTable_5_4_port, keyTable_5_3_port, keyTable_5_2_port, 
      keyTable_5_1_port, keyTable_5_0_port, keyTable_6_7_port, 
      keyTable_6_6_port, keyTable_6_5_port, keyTable_6_4_port, 
      keyTable_6_3_port, keyTable_6_2_port, keyTable_6_1_port, 
      keyTable_6_0_port, keyTable_7_7_port, keyTable_7_6_port, 
      keyTable_7_5_port, keyTable_7_4_port, keyTable_7_3_port, 
      keyTable_7_2_port, keyTable_7_1_port, keyTable_7_0_port, delaydata_7_port
      , delaydata_6_port, delaydata_5_port, delaydata_4_port, delaydata_3_port,
      delaydata_2_port, delaydata_1_port, delaydata_0_port, 
      prefillCounter_7_port, prefillCounter_6_port, prefillCounter_5_port, 
      prefillCounter_4_port, prefillCounter_3_port, prefillCounter_2_port, 
      prefillCounter_1_port, prefillCounter_0_port, faddr_7_port, faddr_6_port,
      faddr_5_port, faddr_4_port, faddr_3_port, faddr_2_port, faddr_1_port, 
      faddr_0_port, nfaddr_7_port, nfaddr_6_port, nfaddr_5_port, nfaddr_4_port,
      nfaddr_3_port, nfaddr_2_port, nfaddr_1_port, nfaddr_0_port, fdata_7_port,
      fdata_6_port, fdata_5_port, fdata_4_port, fdata_3_port, fdata_2_port, 
      fdata_1_port, fdata_0_port, nfdata_7_port, nfdata_6_port, nfdata_5_port, 
      nfdata_4_port, nfdata_3_port, nfdata_2_port, nfdata_1_port, nfdata_0_port
      , fw_enable, fr_enable, N407, N408, N409, N410, N411, N412, N413, N414, 
      N424, N425, N426, N427, N428, N429, N430, N431, N472, N473, N474, N475, 
      N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, 
      N496, N497, N498, N499, N500, N501, N502, N503, N512, N513, N514, N515, 
      N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, 
      n1, n2, n124, n126, n128, n130, n155, n158, n159, n163, n165, n168, n173,
      n174, n176, n186, n204, n588, n589, n691, n693, n694, n695, n696, n697, 
      n698, n699, n700, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n767, n768, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n891, n892, n893, n894, n895, 
      n896, n897, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
      n909, n910, n911, n912, n913, n914, n915, N456, N455, N454, N453, N452, 
      N451, N450, N449, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n125, n127, 
      n129, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n156, n157, n160, n161, n162, n164, n166, n167, n169, n170, n171, 
      n172, n175, n177, n178, n179, n180, n181, n182, n183, n184, n185, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, 
      n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n406, n407_port, n408_port, n409_port, n410_port, n411_port, 
      n412_port, n413_port, n414_port, n415, n416, n417, n418, n419, n420, n421
      , n422, n423, n424_port, n425_port, n426_port, n427_port, n428_port, 
      n429_port, n430_port, n431_port, n432, n433, n434, n435, n436, n437, n438
      , n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449_port, 
      n450_port, n451_port, n452_port, n453_port, n454_port, n455_port, 
      n456_port, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, 
      n467, n468, n469, n470, n471, n472_port, n473_port, n474_port, n475_port,
      n476_port, n477_port, n478_port, n479_port, n480_port, n481_port, 
      n482_port, n483_port, n484_port, n485_port, n486_port, n487_port, n488, 
      n489, n490, n491, n492, n493, n494, n495, n496_port, n497_port, n498_port
      , n499_port, n500_port, n501_port, n502_port, n503_port, n504, n505, n506
      , n507, n508, n509, n510, n511, n512_port, n513_port, n514_port, 
      n515_port, n516_port, n517_port, n518_port, n519_port, n520_port, 
      n521_port, n522_port, n523_port, n524_port, n525_port, n526_port, 
      n527_port, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n692, n701, n765, n766, n769, 
      n770, n783, n784, n785, n786, n787, n788, n789, n790, n791, n864, n865, 
      n866, n867, n868, n869, n870, n871, n883, n884, n885, n886, n887, n888, 
      n889, n890, n898, n916, n917, n918, n919, n920, n921, n922, n923, n924, 
      n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, 
      n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, 
      n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, 
      n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, 
      n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, 
      n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
      n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, 
      n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
      n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, 
      n1138, n_1032, n_1033, n_1034, n_1035 : std_logic;

begin
   PROCESSED_DATA <= ( PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, 
      PROCESSED_DATA_5_port, PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, 
      PROCESSED_DATA_2_port, PROCESSED_DATA_1_port, PROCESSED_DATA_0_port );
   W_ENABLE <= W_ENABLE_port;
   R_ENABLE <= R_ENABLE_port;
   ADDR <= ( ADDR_7_port, ADDR_6_port, ADDR_5_port, ADDR_4_port, ADDR_3_port, 
      ADDR_2_port, ADDR_1_port, ADDR_0_port );
   DATA <= ( DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, 
      DATA_2_port, DATA_1_port, DATA_0_port );
   
   n1 <= '0';
   n2 <= '0';
   prefillCounter_reg_0_inst : DFFPOSX1 port map( D => n915, CLK => CLK, Q => 
                           prefillCounter_0_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n212, S => n782, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n212, S => n781, Q => state_2_port);
   state_reg_4_inst : DFFSR port map( D => nextState_4_port, CLK => CLK, R => 
                           n211, S => n780, Q => state_4_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n211, S => n779, Q => state_0_port);
   permuteComplete_reg : DFFPOSX1 port map( D => n899, CLK => CLK, Q => 
                           permuteComplete);
   state_reg_3_inst : DFFSR port map( D => nextState_3_port, CLK => CLK, R => 
                           n211, S => n778, Q => state_3_port);
   PDATA_READY_reg : DFFSR port map( D => n1135, CLK => CLK, R => n211, S => 
                           n777, Q => PDATA_READY);
   extratemp_reg_7_inst : DFFPOSX1 port map( D => n1134, CLK => CLK, Q => 
                           extratemp_7_port);
   extratemp_reg_6_inst : DFFPOSX1 port map( D => n1133, CLK => CLK, Q => 
                           extratemp_6_port);
   extratemp_reg_5_inst : DFFPOSX1 port map( D => n1132, CLK => CLK, Q => 
                           extratemp_5_port);
   extratemp_reg_4_inst : DFFPOSX1 port map( D => n1131, CLK => CLK, Q => 
                           extratemp_4_port);
   extratemp_reg_3_inst : DFFPOSX1 port map( D => n1130, CLK => CLK, Q => 
                           extratemp_3_port);
   extratemp_reg_2_inst : DFFPOSX1 port map( D => n1129, CLK => CLK, Q => 
                           extratemp_2_port);
   extratemp_reg_1_inst : DFFPOSX1 port map( D => n1128, CLK => CLK, Q => 
                           extratemp_1_port);
   extratemp_reg_0_inst : DFFPOSX1 port map( D => n1127, CLK => CLK, Q => 
                           extratemp_0_port);
   keyTable_reg_7_0_inst : DFFPOSX1 port map( D => n792, CLK => CLK, Q => 
                           keyTable_7_0_port);
   keyTable_reg_7_1_inst : DFFPOSX1 port map( D => n793, CLK => CLK, Q => 
                           keyTable_7_1_port);
   keyTable_reg_7_2_inst : DFFPOSX1 port map( D => n794, CLK => CLK, Q => 
                           keyTable_7_2_port);
   keyTable_reg_7_3_inst : DFFPOSX1 port map( D => n795, CLK => CLK, Q => 
                           keyTable_7_3_port);
   keyTable_reg_7_4_inst : DFFPOSX1 port map( D => n796, CLK => CLK, Q => 
                           keyTable_7_4_port);
   keyTable_reg_7_5_inst : DFFPOSX1 port map( D => n797, CLK => CLK, Q => 
                           keyTable_7_5_port);
   keyTable_reg_7_6_inst : DFFPOSX1 port map( D => n798, CLK => CLK, Q => 
                           keyTable_7_6_port);
   keyTable_reg_7_7_inst : DFFPOSX1 port map( D => n799, CLK => CLK, Q => 
                           keyTable_7_7_port);
   keyTable_reg_6_0_inst : DFFPOSX1 port map( D => n800, CLK => CLK, Q => 
                           keyTable_6_0_port);
   keyTable_reg_6_1_inst : DFFPOSX1 port map( D => n801, CLK => CLK, Q => 
                           keyTable_6_1_port);
   keyTable_reg_6_2_inst : DFFPOSX1 port map( D => n802, CLK => CLK, Q => 
                           keyTable_6_2_port);
   keyTable_reg_6_3_inst : DFFPOSX1 port map( D => n803, CLK => CLK, Q => 
                           keyTable_6_3_port);
   keyTable_reg_6_4_inst : DFFPOSX1 port map( D => n804, CLK => CLK, Q => 
                           keyTable_6_4_port);
   keyTable_reg_6_5_inst : DFFPOSX1 port map( D => n805, CLK => CLK, Q => 
                           keyTable_6_5_port);
   keyTable_reg_6_6_inst : DFFPOSX1 port map( D => n806, CLK => CLK, Q => 
                           keyTable_6_6_port);
   keyTable_reg_6_7_inst : DFFPOSX1 port map( D => n807, CLK => CLK, Q => 
                           keyTable_6_7_port);
   keyTable_reg_5_0_inst : DFFPOSX1 port map( D => n808, CLK => CLK, Q => 
                           keyTable_5_0_port);
   keyTable_reg_5_1_inst : DFFPOSX1 port map( D => n809, CLK => CLK, Q => 
                           keyTable_5_1_port);
   keyTable_reg_5_2_inst : DFFPOSX1 port map( D => n810, CLK => CLK, Q => 
                           keyTable_5_2_port);
   keyTable_reg_5_3_inst : DFFPOSX1 port map( D => n811, CLK => CLK, Q => 
                           keyTable_5_3_port);
   keyTable_reg_5_4_inst : DFFPOSX1 port map( D => n812, CLK => CLK, Q => 
                           keyTable_5_4_port);
   keyTable_reg_5_5_inst : DFFPOSX1 port map( D => n813, CLK => CLK, Q => 
                           keyTable_5_5_port);
   keyTable_reg_5_6_inst : DFFPOSX1 port map( D => n814, CLK => CLK, Q => 
                           keyTable_5_6_port);
   keyTable_reg_5_7_inst : DFFPOSX1 port map( D => n815, CLK => CLK, Q => 
                           keyTable_5_7_port);
   keyTable_reg_4_0_inst : DFFPOSX1 port map( D => n816, CLK => CLK, Q => 
                           keyTable_4_0_port);
   keyTable_reg_4_1_inst : DFFPOSX1 port map( D => n817, CLK => CLK, Q => 
                           keyTable_4_1_port);
   keyTable_reg_4_2_inst : DFFPOSX1 port map( D => n818, CLK => CLK, Q => 
                           keyTable_4_2_port);
   keyTable_reg_4_3_inst : DFFPOSX1 port map( D => n819, CLK => CLK, Q => 
                           keyTable_4_3_port);
   keyTable_reg_4_4_inst : DFFPOSX1 port map( D => n820, CLK => CLK, Q => 
                           keyTable_4_4_port);
   keyTable_reg_4_5_inst : DFFPOSX1 port map( D => n821, CLK => CLK, Q => 
                           keyTable_4_5_port);
   keyTable_reg_4_6_inst : DFFPOSX1 port map( D => n822, CLK => CLK, Q => 
                           keyTable_4_6_port);
   keyTable_reg_4_7_inst : DFFPOSX1 port map( D => n823, CLK => CLK, Q => 
                           keyTable_4_7_port);
   keyTable_reg_3_0_inst : DFFPOSX1 port map( D => n824, CLK => CLK, Q => 
                           keyTable_3_0_port);
   keyTable_reg_3_1_inst : DFFPOSX1 port map( D => n825, CLK => CLK, Q => 
                           keyTable_3_1_port);
   keyTable_reg_3_2_inst : DFFPOSX1 port map( D => n826, CLK => CLK, Q => 
                           keyTable_3_2_port);
   keyTable_reg_3_3_inst : DFFPOSX1 port map( D => n827, CLK => CLK, Q => 
                           keyTable_3_3_port);
   keyTable_reg_3_4_inst : DFFPOSX1 port map( D => n828, CLK => CLK, Q => 
                           keyTable_3_4_port);
   keyTable_reg_3_5_inst : DFFPOSX1 port map( D => n829, CLK => CLK, Q => 
                           keyTable_3_5_port);
   keyTable_reg_3_6_inst : DFFPOSX1 port map( D => n830, CLK => CLK, Q => 
                           keyTable_3_6_port);
   keyTable_reg_3_7_inst : DFFPOSX1 port map( D => n831, CLK => CLK, Q => 
                           keyTable_3_7_port);
   keyTable_reg_2_0_inst : DFFPOSX1 port map( D => n832, CLK => CLK, Q => 
                           keyTable_2_0_port);
   keyTable_reg_2_1_inst : DFFPOSX1 port map( D => n833, CLK => CLK, Q => 
                           keyTable_2_1_port);
   keyTable_reg_2_2_inst : DFFPOSX1 port map( D => n834, CLK => CLK, Q => 
                           keyTable_2_2_port);
   keyTable_reg_2_3_inst : DFFPOSX1 port map( D => n835, CLK => CLK, Q => 
                           keyTable_2_3_port);
   keyTable_reg_2_4_inst : DFFPOSX1 port map( D => n836, CLK => CLK, Q => 
                           keyTable_2_4_port);
   keyTable_reg_2_5_inst : DFFPOSX1 port map( D => n837, CLK => CLK, Q => 
                           keyTable_2_5_port);
   keyTable_reg_2_6_inst : DFFPOSX1 port map( D => n838, CLK => CLK, Q => 
                           keyTable_2_6_port);
   keyTable_reg_2_7_inst : DFFPOSX1 port map( D => n839, CLK => CLK, Q => 
                           keyTable_2_7_port);
   keyTable_reg_1_0_inst : DFFPOSX1 port map( D => n840, CLK => CLK, Q => 
                           keyTable_1_0_port);
   keyTable_reg_1_1_inst : DFFPOSX1 port map( D => n841, CLK => CLK, Q => 
                           keyTable_1_1_port);
   keyTable_reg_1_2_inst : DFFPOSX1 port map( D => n842, CLK => CLK, Q => 
                           keyTable_1_2_port);
   keyTable_reg_1_3_inst : DFFPOSX1 port map( D => n843, CLK => CLK, Q => 
                           keyTable_1_3_port);
   keyTable_reg_1_4_inst : DFFPOSX1 port map( D => n844, CLK => CLK, Q => 
                           keyTable_1_4_port);
   keyTable_reg_1_5_inst : DFFPOSX1 port map( D => n845, CLK => CLK, Q => 
                           keyTable_1_5_port);
   keyTable_reg_1_6_inst : DFFPOSX1 port map( D => n846, CLK => CLK, Q => 
                           keyTable_1_6_port);
   keyTable_reg_0_6_inst : DFFPOSX1 port map( D => n847, CLK => CLK, Q => 
                           keyTable_0_6_port);
   keyTable_reg_0_5_inst : DFFPOSX1 port map( D => n848, CLK => CLK, Q => 
                           keyTable_0_5_port);
   keyTable_reg_0_4_inst : DFFPOSX1 port map( D => n849, CLK => CLK, Q => 
                           keyTable_0_4_port);
   keyTable_reg_0_3_inst : DFFPOSX1 port map( D => n850, CLK => CLK, Q => 
                           keyTable_0_3_port);
   keyTable_reg_0_2_inst : DFFPOSX1 port map( D => n851, CLK => CLK, Q => 
                           keyTable_0_2_port);
   keyTable_reg_0_1_inst : DFFPOSX1 port map( D => n852, CLK => CLK, Q => 
                           keyTable_0_1_port);
   keyTable_reg_0_0_inst : DFFPOSX1 port map( D => n853, CLK => CLK, Q => 
                           keyTable_0_0_port);
   keyTable_reg_1_7_inst : DFFPOSX1 port map( D => n854, CLK => CLK, Q => 
                           keyTable_1_7_port);
   keyTable_reg_0_7_inst : DFFPOSX1 port map( D => n855, CLK => CLK, Q => 
                           keyTable_0_7_port);
   prefillCounter_reg_7_inst : DFFPOSX1 port map( D => n914, CLK => CLK, Q => 
                           prefillCounter_7_port);
   prefillCounter_reg_1_inst : DFFPOSX1 port map( D => n913, CLK => CLK, Q => 
                           prefillCounter_1_port);
   prefillCounter_reg_2_inst : DFFPOSX1 port map( D => n912, CLK => CLK, Q => 
                           prefillCounter_2_port);
   prefillCounter_reg_3_inst : DFFPOSX1 port map( D => n911, CLK => CLK, Q => 
                           prefillCounter_3_port);
   prefillCounter_reg_4_inst : DFFPOSX1 port map( D => n910, CLK => CLK, Q => 
                           prefillCounter_4_port);
   prefillCounter_reg_5_inst : DFFPOSX1 port map( D => n909, CLK => CLK, Q => 
                           prefillCounter_5_port);
   prefillCounter_reg_6_inst : DFFPOSX1 port map( D => n908, CLK => CLK, Q => 
                           prefillCounter_6_port);
   temp_reg_7_inst : DFFPOSX1 port map( D => n856, CLK => CLK, Q => temp_7_port
                           );
   temp_reg_0_inst : DFFPOSX1 port map( D => n863, CLK => CLK, Q => temp_0_port
                           );
   temp_reg_1_inst : DFFPOSX1 port map( D => n862, CLK => CLK, Q => temp_1_port
                           );
   temp_reg_2_inst : DFFPOSX1 port map( D => n861, CLK => CLK, Q => temp_2_port
                           );
   temp_reg_3_inst : DFFPOSX1 port map( D => n860, CLK => CLK, Q => temp_3_port
                           );
   temp_reg_4_inst : DFFPOSX1 port map( D => n859, CLK => CLK, Q => temp_4_port
                           );
   temp_reg_5_inst : DFFPOSX1 port map( D => n858, CLK => CLK, Q => temp_5_port
                           );
   temp_reg_6_inst : DFFPOSX1 port map( D => n857, CLK => CLK, Q => temp_6_port
                           );
   si_reg_0_inst : DFFSR port map( D => n907, CLK => CLK, R => n211, S => n776,
                           Q => si_0_port);
   si_reg_1_inst : DFFSR port map( D => n906, CLK => CLK, R => n210, S => n775,
                           Q => si_1_port);
   si_reg_2_inst : DFFSR port map( D => n905, CLK => CLK, R => n210, S => n774,
                           Q => si_2_port);
   si_reg_3_inst : DFFSR port map( D => n904, CLK => CLK, R => n210, S => n773,
                           Q => si_3_port);
   si_reg_4_inst : DFFSR port map( D => n903, CLK => CLK, R => n209, S => n772,
                           Q => si_4_port);
   si_reg_5_inst : DFFSR port map( D => n902, CLK => CLK, R => n210, S => n771,
                           Q => si_5_port);
   delaydata_reg_7_inst : DFFPOSX1 port map( D => n1111, CLK => CLK, Q => 
                           delaydata_7_port);
   delaydata_reg_0_inst : DFFPOSX1 port map( D => n1118, CLK => CLK, Q => 
                           delaydata_0_port);
   delaydata_reg_1_inst : DFFPOSX1 port map( D => n1117, CLK => CLK, Q => 
                           delaydata_1_port);
   delaydata_reg_2_inst : DFFPOSX1 port map( D => n1116, CLK => CLK, Q => 
                           delaydata_2_port);
   delaydata_reg_3_inst : DFFPOSX1 port map( D => n1115, CLK => CLK, Q => 
                           delaydata_3_port);
   delaydata_reg_4_inst : DFFPOSX1 port map( D => n1114, CLK => CLK, Q => 
                           delaydata_4_port);
   delaydata_reg_5_inst : DFFPOSX1 port map( D => n1113, CLK => CLK, Q => 
                           delaydata_5_port);
   delaydata_reg_6_inst : DFFPOSX1 port map( D => n1112, CLK => CLK, Q => 
                           delaydata_6_port);
   intj_reg_7_inst : DFFPOSX1 port map( D => n875, CLK => CLK, Q => intj_7_port
                           );
   intj_reg_0_inst : DFFPOSX1 port map( D => n882, CLK => CLK, Q => intj_0_port
                           );
   intj_reg_1_inst : DFFPOSX1 port map( D => n881, CLK => CLK, Q => intj_1_port
                           );
   intj_reg_2_inst : DFFPOSX1 port map( D => n880, CLK => CLK, Q => intj_2_port
                           );
   intj_reg_3_inst : DFFPOSX1 port map( D => n879, CLK => CLK, Q => intj_3_port
                           );
   intj_reg_4_inst : DFFPOSX1 port map( D => n878, CLK => CLK, Q => intj_4_port
                           );
   intj_reg_5_inst : DFFPOSX1 port map( D => n877, CLK => CLK, Q => intj_5_port
                           );
   intj_reg_6_inst : DFFPOSX1 port map( D => n876, CLK => CLK, Q => intj_6_port
                           );
   sj_reg_7_inst : DFFSR port map( D => n1099, CLK => CLK, R => n209, S => n768
                           , Q => sj_7_port);
   sj_reg_6_inst : DFFSR port map( D => n897, CLK => CLK, R => n209, S => n767,
                           Q => sj_6_port);
   sj_reg_3_inst : DFFSR port map( D => n894, CLK => CLK, R => n208, S => n764,
                           Q => sj_3_port);
   sj_reg_2_inst : DFFSR port map( D => n893, CLK => CLK, R => n208, S => n763,
                           Q => sj_2_port);
   sj_reg_1_inst : DFFSR port map( D => n892, CLK => CLK, R => n208, S => n762,
                           Q => sj_1_port);
   sj_reg_0_inst : DFFSR port map( D => n891, CLK => CLK, R => n207, S => n761,
                           Q => sj_0_port);
   keyi_reg_2_inst : DFFPOSX1 port map( D => n874, CLK => CLK, Q => keyi_2_port
                           );
   keyi_reg_1_inst : DFFPOSX1 port map( D => n873, CLK => CLK, Q => keyi_1_port
                           );
   keyi_reg_0_inst : DFFPOSX1 port map( D => n872, CLK => CLK, Q => keyi_0_port
                           );
   inti_reg_7_inst : DFFPOSX1 port map( D => n1126, CLK => CLK, Q => 
                           inti_7_port);
   inti_reg_0_inst : DFFPOSX1 port map( D => n1119, CLK => CLK, Q => 
                           inti_0_port);
   inti_reg_1_inst : DFFPOSX1 port map( D => n1120, CLK => CLK, Q => 
                           inti_1_port);
   inti_reg_2_inst : DFFPOSX1 port map( D => n1121, CLK => CLK, Q => 
                           inti_2_port);
   inti_reg_3_inst : DFFPOSX1 port map( D => n1122, CLK => CLK, Q => 
                           inti_3_port);
   inti_reg_4_inst : DFFPOSX1 port map( D => n1123, CLK => CLK, Q => 
                           inti_4_port);
   inti_reg_5_inst : DFFPOSX1 port map( D => n1124, CLK => CLK, Q => 
                           inti_5_port);
   inti_reg_6_inst : DFFPOSX1 port map( D => n1125, CLK => CLK, Q => 
                           inti_6_port);
   currentProcessedData_reg_0_inst : DFFSR port map( D => 
                           nextProcessedData_0_port, CLK => CLK, R => n207, S 
                           => n760, Q => currentProcessedData_0_port);
   PROCESSED_DATA_reg_0_inst : DFFPOSX1 port map( D => n759, CLK => CLK, Q => 
                           PROCESSED_DATA_0_port);
   currentProcessedData_reg_1_inst : DFFSR port map( D => 
                           nextProcessedData_1_port, CLK => CLK, R => n206, S 
                           => n758, Q => currentProcessedData_1_port);
   PROCESSED_DATA_reg_1_inst : DFFPOSX1 port map( D => n757, CLK => CLK, Q => 
                           PROCESSED_DATA_1_port);
   currentProcessedData_reg_2_inst : DFFSR port map( D => n37, CLK => CLK, R =>
                           n206, S => n756, Q => currentProcessedData_2_port);
   PROCESSED_DATA_reg_2_inst : DFFPOSX1 port map( D => n755, CLK => CLK, Q => 
                           PROCESSED_DATA_2_port);
   currentProcessedData_reg_3_inst : DFFSR port map( D => n38, CLK => CLK, R =>
                           n205, S => n754, Q => currentProcessedData_3_port);
   PROCESSED_DATA_reg_3_inst : DFFPOSX1 port map( D => n753, CLK => CLK, Q => 
                           PROCESSED_DATA_3_port);
   currentProcessedData_reg_4_inst : DFFSR port map( D => n39, CLK => CLK, R =>
                           n205, S => n752, Q => currentProcessedData_4_port);
   PROCESSED_DATA_reg_4_inst : DFFPOSX1 port map( D => n751, CLK => CLK, Q => 
                           PROCESSED_DATA_4_port);
   currentProcessedData_reg_5_inst : DFFSR port map( D => n40, CLK => CLK, R =>
                           n203, S => n750, Q => currentProcessedData_5_port);
   PROCESSED_DATA_reg_5_inst : DFFPOSX1 port map( D => n749, CLK => CLK, Q => 
                           PROCESSED_DATA_5_port);
   currentProcessedData_reg_6_inst : DFFSR port map( D => n95, CLK => CLK, R =>
                           n203, S => n748, Q => currentProcessedData_6_port);
   PROCESSED_DATA_reg_6_inst : DFFPOSX1 port map( D => n747, CLK => CLK, Q => 
                           PROCESSED_DATA_6_port);
   currentProcessedData_reg_7_inst : DFFSR port map( D => 
                           nextProcessedData_7_port, CLK => CLK, R => n210, S 
                           => n746, Q => currentProcessedData_7_port);
   PROCESSED_DATA_reg_7_inst : DFFPOSX1 port map( D => n745, CLK => CLK, Q => 
                           PROCESSED_DATA_7_port);
   faddr_reg_7_inst : DFFPOSX1 port map( D => n744, CLK => CLK, Q => 
                           faddr_7_port);
   ADDR_reg_7_inst : DFFPOSX1 port map( D => n743, CLK => CLK, Q => ADDR_7_port
                           );
   faddr_reg_6_inst : DFFPOSX1 port map( D => n742, CLK => CLK, Q => 
                           faddr_6_port);
   ADDR_reg_6_inst : DFFPOSX1 port map( D => n741, CLK => CLK, Q => ADDR_6_port
                           );
   faddr_reg_5_inst : DFFPOSX1 port map( D => n740, CLK => CLK, Q => 
                           faddr_5_port);
   ADDR_reg_5_inst : DFFPOSX1 port map( D => n739, CLK => CLK, Q => ADDR_5_port
                           );
   faddr_reg_4_inst : DFFPOSX1 port map( D => n738, CLK => CLK, Q => 
                           faddr_4_port);
   ADDR_reg_4_inst : DFFPOSX1 port map( D => n737, CLK => CLK, Q => ADDR_4_port
                           );
   faddr_reg_3_inst : DFFPOSX1 port map( D => n736, CLK => CLK, Q => 
                           faddr_3_port);
   ADDR_reg_3_inst : DFFPOSX1 port map( D => n735, CLK => CLK, Q => ADDR_3_port
                           );
   faddr_reg_2_inst : DFFPOSX1 port map( D => n734, CLK => CLK, Q => 
                           faddr_2_port);
   ADDR_reg_2_inst : DFFPOSX1 port map( D => n733, CLK => CLK, Q => ADDR_2_port
                           );
   faddr_reg_1_inst : DFFPOSX1 port map( D => n732, CLK => CLK, Q => 
                           faddr_1_port);
   ADDR_reg_1_inst : DFFPOSX1 port map( D => n731, CLK => CLK, Q => ADDR_1_port
                           );
   faddr_reg_0_inst : DFFPOSX1 port map( D => n730, CLK => CLK, Q => 
                           faddr_0_port);
   ADDR_reg_0_inst : DFFPOSX1 port map( D => n729, CLK => CLK, Q => ADDR_0_port
                           );
   fdata_reg_7_inst : DFFPOSX1 port map( D => n728, CLK => CLK, Q => 
                           fdata_7_port);
   fdata_reg_6_inst : DFFPOSX1 port map( D => n727, CLK => CLK, Q => 
                           fdata_6_port);
   fdata_reg_5_inst : DFFPOSX1 port map( D => n726, CLK => CLK, Q => 
                           fdata_5_port);
   fdata_reg_4_inst : DFFPOSX1 port map( D => n725, CLK => CLK, Q => 
                           fdata_4_port);
   fdata_reg_3_inst : DFFPOSX1 port map( D => n724, CLK => CLK, Q => 
                           fdata_3_port);
   fdata_reg_2_inst : DFFPOSX1 port map( D => n723, CLK => CLK, Q => 
                           fdata_2_port);
   fdata_reg_1_inst : DFFPOSX1 port map( D => n722, CLK => CLK, Q => 
                           fdata_1_port);
   fdata_reg_0_inst : DFFPOSX1 port map( D => n721, CLK => CLK, Q => 
                           fdata_0_port);
   fw_enable_reg : DFFPOSX1 port map( D => n720, CLK => CLK, Q => fw_enable);
   fr_enable_reg : DFFPOSX1 port map( D => n719, CLK => CLK, Q => fr_enable);
   W_ENABLE_reg : DFFPOSX1 port map( D => n718, CLK => CLK, Q => W_ENABLE_port)
                           ;
   R_ENABLE_reg : DFFPOSX1 port map( D => n717, CLK => CLK, Q => R_ENABLE_port)
                           ;
   DATA_reg_7_inst : DFFPOSX1 port map( D => n716, CLK => CLK, Q => DATA_7_port
                           );
   DATA_reg_6_inst : DFFPOSX1 port map( D => n715, CLK => CLK, Q => DATA_6_port
                           );
   DATA_reg_5_inst : DFFPOSX1 port map( D => n714, CLK => CLK, Q => DATA_5_port
                           );
   DATA_reg_4_inst : DFFPOSX1 port map( D => n713, CLK => CLK, Q => DATA_4_port
                           );
   DATA_reg_3_inst : DFFPOSX1 port map( D => n712, CLK => CLK, Q => DATA_3_port
                           );
   DATA_reg_2_inst : DFFPOSX1 port map( D => n711, CLK => CLK, Q => DATA_2_port
                           );
   DATA_reg_1_inst : DFFPOSX1 port map( D => n710, CLK => CLK, Q => DATA_1_port
                           );
   DATA_reg_0_inst : DFFPOSX1 port map( D => n709, CLK => CLK, Q => DATA_0_port
                           );
   U110 : NOR2X1 port map( A => KEY_ERROR, B => n128, Y => n126);
   U111 : OAI21X1 port map( A => n1107, B => n130, C => n1106, Y => n124);
   U123 : NOR2X1 port map( A => n159, B => n1107, Y => n155);
   U126 : NAND3X1 port map( A => n163, B => n1101, C => n165, Y => 
                           nextState_1_port);
   U130 : NOR2X1 port map( A => prefillCounter_2_port, B => 
                           prefillCounter_1_port, Y => n173);
   U131 : NAND3X1 port map( A => n174, B => n1136, C => n176, Y => n168);
   U132 : NOR2X1 port map( A => prefillCounter_4_port, B => 
                           prefillCounter_3_port, Y => n176);
   U133 : NOR2X1 port map( A => prefillCounter_7_port, B => 
                           prefillCounter_6_port, Y => n174);
   U143 : NAND3X1 port map( A => n1110, B => n1109, C => BYTE_READY, Y => n158)
                           ;
   U156 : NAND2X1 port map( A => OPCODE(0), B => n1109, Y => n130);
   U158 : NAND2X1 port map( A => BYTE_READY, B => n204, Y => n128);
   U159 : OAI21X1 port map( A => OPCODE(0), B => OPCODE(1), C => n186, Y => 
                           n204);
   U160 : NAND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n186);
   U669 : NOR2X1 port map( A => n1104, B => n1105, Y => n588);
   U673 : NOR2X1 port map( A => n1102, B => n1103, Y => n589);
   n746 <= '1';
   n748 <= '1';
   n750 <= '1';
   n752 <= '1';
   n754 <= '1';
   n756 <= '1';
   n758 <= '1';
   n760 <= '1';
   n761 <= '1';
   n762 <= '1';
   n763 <= '1';
   n764 <= '1';
   n767 <= '1';
   n768 <= '1';
   n771 <= '1';
   n772 <= '1';
   n773 <= '1';
   n774 <= '1';
   n775 <= '1';
   n776 <= '1';
   n777 <= '1';
   n778 <= '1';
   n779 <= '1';
   n780 <= '1';
   n781 <= '1';
   n782 <= '1';
   U142 : AND2X2 port map( A => n130, B => n186, Y => n159);
   add_289 : KSA_1_DW01_inc_0 port map( A(7) => si_7_port, A(6) => si_6_port, 
                           A(5) => si_5_port, A(4) => si_4_port, A(3) => 
                           si_3_port, A(2) => si_2_port, A(1) => si_1_port, 
                           A(0) => n24, SUM(7) => N431, SUM(6) => N430, SUM(5) 
                           => N429, SUM(4) => N428, SUM(3) => N427, SUM(2) => 
                           N426, SUM(1) => N425, SUM(0) => N424);
   add_263 : KSA_1_DW01_inc_1 port map( A(7) => prefillCounter_7_port, A(6) => 
                           prefillCounter_6_port, A(5) => prefillCounter_5_port
                           , A(4) => prefillCounter_4_port, A(3) => 
                           prefillCounter_3_port, A(2) => prefillCounter_2_port
                           , A(1) => prefillCounter_1_port, A(0) => 
                           prefillCounter_0_port, SUM(7) => N414, SUM(6) => 
                           N413, SUM(5) => N412, SUM(4) => N411, SUM(3) => N410
                           , SUM(2) => N409, SUM(1) => N408, SUM(0) => N407);
   add_377 : KSA_1_DW01_add_6 port map( A(7) => temp_7_port, A(6) => 
                           temp_6_port, A(5) => temp_5_port, A(4) => 
                           temp_4_port, A(3) => temp_3_port, A(2) => 
                           temp_2_port, A(1) => temp_1_port, A(0) => 
                           temp_0_port, B(7) => extratemp_7_port, B(6) => 
                           extratemp_6_port, B(5) => extratemp_5_port, B(4) => 
                           extratemp_4_port, B(3) => extratemp_3_port, B(2) => 
                           extratemp_2_port, B(1) => extratemp_1_port, B(0) => 
                           extratemp_0_port, CI => n1, SUM(7) => N527, SUM(6) 
                           => N526, SUM(5) => N525, SUM(4) => N524, SUM(3) => 
                           N523, SUM(2) => N522, SUM(1) => N521, SUM(0) => N520
                           , CO => n_1032);
   add_337 : KSA_1_DW01_add_7 port map( A(7) => intj_7_port, A(6) => 
                           intj_6_port, A(5) => intj_5_port, A(4) => 
                           intj_4_port, A(3) => intj_3_port, A(2) => 
                           intj_2_port, A(1) => intj_1_port, A(0) => 
                           intj_0_port, B(7) => DATA_IN(7), B(6) => DATA_IN(6),
                           B(5) => DATA_IN(5), B(4) => DATA_IN(4), B(3) => 
                           DATA_IN(3), B(2) => DATA_IN(2), B(1) => DATA_IN(1), 
                           B(0) => DATA_IN(0), CI => n2, SUM(7) => N519, SUM(6)
                           => N518, SUM(5) => N517, SUM(4) => N516, SUM(3) => 
                           N515, SUM(2) => N514, SUM(1) => N513, SUM(0) => N512
                           , CO => n_1033);
   add_1_root_add_0_root_add_302_2 : KSA_1_DW01_add_8 port map( A(7) => 
                           DATA_IN(7), A(6) => DATA_IN(6), A(5) => DATA_IN(5), 
                           A(4) => DATA_IN(4), A(3) => DATA_IN(3), A(2) => 
                           DATA_IN(2), A(1) => DATA_IN(1), A(0) => DATA_IN(0), 
                           B(7) => sj_7_port, B(6) => sj_6_port, B(5) => 
                           sj_5_port, B(4) => sj_4_port, B(3) => sj_3_port, 
                           B(2) => sj_2_port, B(1) => sj_1_port, B(0) => n48, 
                           CI => n1137, SUM(7) => N456, SUM(6) => N455, SUM(5) 
                           => N454, SUM(4) => N453, SUM(3) => N452, SUM(2) => 
                           N451, SUM(1) => N450, SUM(0) => N449, CO => n_1034);
   add_0_root_add_0_root_add_302_2 : KSA_1_DW01_add_9 port map( A(7) => N472, 
                           A(6) => N473, A(5) => N474, A(4) => N475, A(3) => 
                           N476, A(2) => N477, A(1) => N478, A(0) => N479, B(7)
                           => N456, B(6) => N455, B(5) => N454, B(4) => N453, 
                           B(3) => N452, B(2) => N451, B(1) => N450, B(0) => 
                           N449, CI => n1138, SUM(7) => N487, SUM(6) => N486, 
                           SUM(5) => N485, SUM(4) => N484, SUM(3) => N483, 
                           SUM(2) => N482, SUM(1) => N481, SUM(0) => N480, CO 
                           => n_1035);
   r126 : KSA_1_DW01_inc_3 port map( A(7) => inti_7_port, A(6) => inti_6_port, 
                           A(5) => inti_5_port, A(4) => inti_4_port, A(3) => 
                           inti_3_port, A(2) => inti_2_port, A(1) => 
                           inti_1_port, A(0) => inti_0_port, SUM(7) => N503, 
                           SUM(6) => N502, SUM(5) => N501, SUM(4) => N500, 
                           SUM(3) => N499, SUM(2) => N498, SUM(1) => N497, 
                           SUM(0) => N496);
   nfaddr_tri_0_inst : TBUFX1 port map( A => n708, EN => n1100, Y => 
                           nfaddr_0_port);
   nfaddr_tri_1_inst : TBUFX1 port map( A => n707, EN => n1100, Y => 
                           nfaddr_1_port);
   nfaddr_tri_2_inst : TBUFX1 port map( A => n706, EN => n1100, Y => 
                           nfaddr_2_port);
   nfaddr_tri_3_inst : TBUFX1 port map( A => n705, EN => n1100, Y => 
                           nfaddr_3_port);
   nfaddr_tri_4_inst : TBUFX1 port map( A => n704, EN => n1100, Y => 
                           nfaddr_4_port);
   nfaddr_tri_5_inst : TBUFX1 port map( A => n703, EN => n1100, Y => 
                           nfaddr_5_port);
   nfdata_tri_1_inst : TBUFX1 port map( A => n698, EN => n29, Y => 
                           nfdata_1_port);
   nfdata_tri_2_inst : TBUFX1 port map( A => n697, EN => n29, Y => 
                           nfdata_2_port);
   nfdata_tri_3_inst : TBUFX1 port map( A => n696, EN => n29, Y => 
                           nfdata_3_port);
   nfdata_tri_4_inst : TBUFX1 port map( A => n695, EN => n29, Y => 
                           nfdata_4_port);
   nfdata_tri_5_inst : TBUFX1 port map( A => n694, EN => n29, Y => 
                           nfdata_5_port);
   nfdata_tri_6_inst : TBUFX1 port map( A => n693, EN => n29, Y => 
                           nfdata_6_port);
   nfdata_tri_7_inst : TBUFX1 port map( A => n691, EN => n29, Y => 
                           nfdata_7_port);
   nfaddr_tri_7_inst : TBUFX2 port map( A => n700, EN => n1100, Y => 
                           nfaddr_7_port);
   nfaddr_tri_6_inst : TBUFX1 port map( A => n702, EN => n1100, Y => 
                           nfaddr_6_port);
   nfdata_tri_0_inst : TBUFX1 port map( A => n699, EN => n29, Y => 
                           nfdata_0_port);
   si_reg_6_inst : DFFSR port map( D => n901, CLK => CLK, R => n199, S => n16, 
                           Q => si_6_port);
   si_reg_7_inst : DFFSR port map( D => n900, CLK => CLK, R => n199, S => n15, 
                           Q => si_7_port);
   sj_reg_5_inst : DFFSR port map( D => n896, CLK => CLK, R => n199, S => n14, 
                           Q => sj_5_port);
   sj_reg_4_inst : DFFSR port map( D => n895, CLK => CLK, R => n199, S => n13, 
                           Q => sj_4_port);
   U3 : INVX8 port map( A => n63, Y => n136);
   U4 : NAND2X1 port map( A => n54, B => n1090, Y => n3);
   U7 : AND2X1 port map( A => n70, B => n58, Y => n4);
   U8 : AND2X2 port map( A => n591, B => n590, Y => n5);
   U9 : BUFX4 port map( A => n154, Y => n143);
   U10 : INVX2 port map( A => n31, Y => n552);
   U11 : INVX2 port map( A => n47, Y => n563);
   U12 : INVX2 port map( A => n183, Y => n1081);
   U13 : INVX2 port map( A => n269, Y => n30);
   U14 : INVX2 port map( A => n188, Y => n189);
   U15 : INVX2 port map( A => n89, Y => n67);
   U16 : INVX2 port map( A => n89, Y => n70);
   U17 : OR2X2 port map( A => n1025, B => n1024, Y => n6);
   U18 : INVX2 port map( A => n682, Y => n429_port);
   U19 : NAND2X1 port map( A => n135, B => n1082, Y => n7);
   U20 : OR2X1 port map( A => n119, B => n120, Y => n8);
   U21 : AND2X2 port map( A => n481_port, B => n482_port, Y => n9);
   U22 : AND2X2 port map( A => n473_port, B => n474_port, Y => n10);
   U23 : AND2X2 port map( A => n437, B => n438, Y => n11);
   U24 : AND2X2 port map( A => n107, B => n76, Y => n12);
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   U29 : NAND3X1 port map( A => n162, B => n70, C => n238, Y => n17);
   U30 : INVX2 port map( A => n244, Y => n18);
   U31 : BUFX2 port map( A => n242, Y => n142);
   U32 : BUFX2 port map( A => n72, Y => n19);
   U33 : AOI21X1 port map( A => n177, B => n18, C => n88, Y => n20);
   U34 : BUFX4 port map( A => n1026, Y => n21);
   U35 : NOR2X1 port map( A => n75, B => n74, Y => n22);
   U36 : AND2X2 port map( A => n433, B => n432, Y => n23);
   U37 : BUFX2 port map( A => si_0_port, Y => n24);
   U38 : AND2X2 port map( A => n49, B => n32, Y => n25);
   U39 : INVX2 port map( A => n25, Y => n240);
   U40 : INVX2 port map( A => n240, Y => n1046);
   U41 : AND2X2 port map( A => n64, B => n237, Y => n26);
   U42 : INVX1 port map( A => n1060, Y => n1084);
   U43 : INVX1 port map( A => n66, Y => n27);
   U44 : INVX2 port map( A => n49, Y => n243);
   U45 : INVX1 port map( A => n119, Y => n28);
   U46 : INVX2 port map( A => n135, Y => n119);
   U47 : INVX4 port map( A => n76, Y => n223);
   U48 : INVX1 port map( A => n645, Y => n29);
   U49 : NOR3X1 port map( A => n510, B => n512_port, C => keyi_2_port, Y => n31
                           );
   U50 : INVX4 port map( A => keyi_1_port, Y => n510);
   U51 : INVX4 port map( A => keyi_0_port, Y => n512_port);
   U52 : INVX4 port map( A => keyi_2_port, Y => n511);
   U53 : BUFX2 port map( A => n161, Y => n32);
   U54 : NAND2X1 port map( A => n644, B => n115, Y => n33);
   U55 : INVX2 port map( A => n114, Y => n115);
   U56 : INVX1 port map( A => n18, Y => n34);
   U57 : INVX1 port map( A => n7, Y => n645);
   U58 : MUX2X1 port map( B => n640, A => n511, S => n35, Y => n874);
   U59 : NAND2X1 port map( A => n92, B => n563, Y => n35);
   U60 : INVX1 port map( A => n429_port, Y => n36);
   U61 : INVX1 port map( A => n471, Y => n37);
   U62 : INVX1 port map( A => n465, Y => n38);
   U63 : INVX1 port map( A => n459, Y => n39);
   U64 : INVX1 port map( A => n453_port, Y => n40);
   U65 : NAND2X1 port map( A => n41, B => n432, Y => n297);
   U66 : NOR2X1 port map( A => n47, B => n1135, Y => n41);
   U67 : INVX2 port map( A => n101, Y => n432);
   U68 : AND2X2 port map( A => n183, B => n161, Y => n62);
   U69 : AND2X1 port map( A => n680, B => n681, Y => n42);
   U70 : NAND2X1 port map( A => n644, B => n115, Y => n43);
   U71 : NAND2X1 port map( A => n644, B => n115, Y => n44);
   U72 : INVX1 port map( A => n487_port, Y => n45);
   U73 : INVX1 port map( A => n45, Y => n46);
   U74 : NAND2X1 port map( A => n188, B => n273, Y => n242);
   U75 : BUFX2 port map( A => state_2_port, Y => n179);
   U76 : AND2X2 port map( A => n178, B => n1082, Y => n47);
   U77 : BUFX4 port map( A => sj_0_port, Y => n48);
   U78 : AND2X2 port map( A => n189, B => n273, Y => n49);
   U79 : NAND3X1 port map( A => n96, B => n110, C => n223, Y => n50);
   U80 : NOR2X1 port map( A => n562, B => n47, Y => n51);
   U81 : INVX2 port map( A => n57, Y => n562);
   U82 : BUFX2 port map( A => n562, Y => n52);
   U83 : BUFX4 port map( A => n185, Y => n53);
   U84 : AND2X2 port map( A => n585, B => n1048, Y => n54);
   U85 : INVX4 port map( A => n5, Y => n55);
   U86 : MUX2X1 port map( B => n1102, A => n512_port, S => n56, Y => n872);
   U87 : NAND2X1 port map( A => n563, B => n92, Y => n56);
   U88 : AND2X2 port map( A => n670, B => n646, Y => n57);
   U89 : INVX2 port map( A => n1077, Y => n58);
   U90 : AND2X2 port map( A => n90, B => n638, Y => n59);
   U91 : INVX1 port map( A => n59, Y => n328);
   U92 : INVX1 port map( A => n434, Y => n479_port);
   U93 : AND2X2 port map( A => n7, B => n42, Y => n60);
   U94 : INVX1 port map( A => n60, Y => n1025);
   U95 : MUX2X1 port map( B => fdata_7_port, A => nfdata_7_port, S => n206, Y 
                           => n412_port);
   U96 : MUX2X1 port map( B => fdata_6_port, A => nfdata_6_port, S => n205, Y 
                           => n411_port);
   U97 : MUX2X1 port map( B => fdata_5_port, A => nfdata_5_port, S => n205, Y 
                           => n410_port);
   U98 : MUX2X1 port map( B => fdata_4_port, A => nfdata_4_port, S => n205, Y 
                           => n409_port);
   U99 : MUX2X1 port map( B => fdata_3_port, A => nfdata_3_port, S => n205, Y 
                           => n408_port);
   U100 : MUX2X1 port map( B => fdata_2_port, A => nfdata_2_port, S => n205, Y 
                           => n407_port);
   U101 : MUX2X1 port map( B => fdata_1_port, A => nfdata_1_port, S => n205, Y 
                           => n406);
   U102 : MUX2X1 port map( B => fdata_0_port, A => nfdata_0_port, S => n205, Y 
                           => n405);
   U103 : MUX2X1 port map( B => DATA_7_port, A => nfdata_7_port, S => n205, Y 
                           => n386);
   U104 : MUX2X1 port map( B => DATA_6_port, A => nfdata_6_port, S => n205, Y 
                           => n385);
   U105 : MUX2X1 port map( B => DATA_5_port, A => nfdata_5_port, S => n205, Y 
                           => n384);
   U106 : MUX2X1 port map( B => DATA_4_port, A => nfdata_4_port, S => n203, Y 
                           => n383);
   U107 : MUX2X1 port map( B => DATA_3_port, A => nfdata_3_port, S => n203, Y 
                           => n382);
   U108 : MUX2X1 port map( B => DATA_2_port, A => nfdata_2_port, S => n203, Y 
                           => n381);
   U109 : MUX2X1 port map( B => DATA_1_port, A => nfdata_1_port, S => n205, Y 
                           => n380);
   U112 : AND2X2 port map( A => n682, B => n153, Y => n430_port);
   U113 : MUX2X1 port map( B => DATA_0_port, A => nfdata_0_port, S => n199, Y 
                           => n379);
   U114 : MUX2X1 port map( B => n1103, A => n510, S => n61, Y => n873);
   U115 : NAND2X1 port map( A => n563, B => n92, Y => n61);
   U116 : INVX1 port map( A => n62, Y => n274);
   U117 : INVX2 port map( A => n108, Y => n63);
   U118 : INVX2 port map( A => n108, Y => n154);
   U119 : BUFX4 port map( A => state_4_port, Y => n197);
   U120 : AND2X2 port map( A => n182, B => n139, Y => n64);
   U121 : INVX1 port map( A => n64, Y => n220);
   U122 : INVX1 port map( A => n66, Y => n111);
   U124 : NAND2X1 port map( A => n246, B => n1082, Y => n65);
   U125 : BUFX2 port map( A => state_1_port, Y => n66);
   U127 : NAND2X1 port map( A => n684, B => n141, Y => n68);
   U128 : INVX4 port map( A => n237, Y => n105);
   U129 : NAND2X1 port map( A => n237, B => n169, Y => n69);
   U134 : INVX2 port map( A => n69, Y => n135);
   U135 : INVX1 port map( A => n194, Y => n131);
   U136 : BUFX2 port map( A => state_0_port, Y => n182);
   U137 : INVX1 port map( A => sj_2_port, Y => n572);
   U138 : INVX2 port map( A => n297, Y => n71);
   U139 : AND2X2 port map( A => n96, B => n64, Y => n72);
   U140 : NOR2X1 port map( A => n47, B => n156, Y => n73);
   U141 : NOR2X1 port map( A => n75, B => n74, Y => n565);
   U144 : INVX1 port map( A => n73, Y => n74);
   U145 : BUFX4 port map( A => n564, Y => n75);
   U146 : NOR2X1 port map( A => n94, B => n486_port, Y => n629);
   U147 : INVX1 port map( A => n486_port, Y => n1100);
   U148 : INVX4 port map( A => n133, Y => n1135);
   U149 : BUFX4 port map( A => state_0_port, Y => n76);
   U150 : NAND2X1 port map( A => n190, B => n51, Y => n1026);
   U151 : AND2X2 port map( A => n18, B => n1071, Y => n156);
   U152 : INVX4 port map( A => n195, Y => n196);
   U153 : INVX8 port map( A => n136, Y => n77);
   U154 : INVX8 port map( A => n136, Y => n78);
   U155 : INVX4 port map( A => n148, Y => n79);
   U157 : INVX8 port map( A => n79, Y => n80);
   U161 : INVX4 port map( A => n198, Y => n81);
   U162 : INVX8 port map( A => n81, Y => n82);
   U163 : NOR2X1 port map( A => n245, B => n25, Y => n83);
   U164 : AND2X2 port map( A => n83, B => n84, Y => n289);
   U165 : AND2X1 port map( A => n8, B => n670, Y => n84);
   U166 : INVX1 port map( A => n50, Y => n85);
   U167 : INVX1 port map( A => n50, Y => n246);
   U168 : AND2X2 port map( A => n566, B => n86, Y => n152);
   U169 : AND2X1 port map( A => n565, B => n591, Y => n86);
   U170 : BUFX2 port map( A => n169, Y => n87);
   U171 : INVX1 port map( A => n436, Y => n480_port);
   U172 : INVX4 port map( A => n297, Y => n650);
   U173 : INVX2 port map( A => n139, Y => n184);
   U174 : AND2X2 port map( A => n32, B => n1082, Y => n88);
   U175 : INVX2 port map( A => n88, Y => n560);
   U176 : AND2X1 port map( A => n193, B => n123, Y => n649);
   U177 : INVX2 port map( A => n131, Y => n132);
   U178 : AND2X2 port map( A => n167, B => n26, Y => n89);
   U179 : NOR2X1 port map( A => n354, B => si_2_port, Y => n90);
   U180 : INVX1 port map( A => n90, Y => n341);
   U181 : INVX1 port map( A => si_2_port, Y => n640);
   U182 : NOR2X1 port map( A => n1046, B => n245, Y => n91);
   U183 : AND2X2 port map( A => n507, B => n4, Y => n92);
   U184 : INVX1 port map( A => n92, Y => n1057);
   U185 : BUFX2 port map( A => n1089, Y => n93);
   U186 : INVX1 port map( A => si_1_port, Y => n1103);
   U187 : NAND2X1 port map( A => n70, B => n563, Y => n94);
   U188 : NAND2X1 port map( A => n483_port, B => n9, Y => 
                           nextProcessedData_0_port);
   U189 : INVX1 port map( A => nextProcessedData_0_port, Y => n485_port);
   U190 : NAND2X1 port map( A => n475_port, B => n10, Y => 
                           nextProcessedData_1_port);
   U191 : INVX1 port map( A => nextProcessedData_1_port, Y => n477_port);
   U192 : INVX1 port map( A => n447, Y => n95);
   U193 : BUFX4 port map( A => state_4_port, Y => n96);
   U194 : OR2X1 port map( A => n562, B => n561, Y => n97);
   U195 : NAND2X1 port map( A => n1090, B => n157, Y => n98);
   U196 : INVX4 port map( A => n195, Y => n99);
   U197 : INVX1 port map( A => n223, Y => n100);
   U198 : NAND2X1 port map( A => n121, B => n20, Y => n101);
   U199 : NAND2X1 port map( A => n23, B => n629, Y => n102);
   U200 : NAND2X1 port map( A => n23, B => n629, Y => n103);
   U201 : NAND2X1 port map( A => n289, B => n54, Y => n104);
   U202 : INVX2 port map( A => n195, Y => n122);
   U203 : INVX1 port map( A => n785, Y => n683);
   U204 : BUFX2 port map( A => n585, Y => n106);
   U205 : AND2X1 port map( A => n328, B => si_4_port, Y => n316);
   U206 : INVX1 port map( A => n24, Y => n1102);
   U207 : OR2X2 port map( A => n213, B => n181, Y => n1065);
   U208 : INVX1 port map( A => n144, Y => n107);
   U209 : INVX4 port map( A => n674, Y => n195);
   U210 : INVX1 port map( A => n412_port, Y => n728);
   U211 : INVX1 port map( A => n411_port, Y => n727);
   U212 : INVX1 port map( A => n410_port, Y => n726);
   U213 : INVX1 port map( A => n409_port, Y => n725);
   U214 : INVX1 port map( A => n408_port, Y => n724);
   U215 : INVX1 port map( A => n407_port, Y => n723);
   U216 : INVX1 port map( A => n406, Y => n722);
   U217 : INVX1 port map( A => n386, Y => n716);
   U218 : INVX1 port map( A => n385, Y => n715);
   U219 : INVX1 port map( A => n384, Y => n714);
   U220 : INVX1 port map( A => n383, Y => n713);
   U221 : INVX1 port map( A => n382, Y => n712);
   U222 : INVX1 port map( A => n381, Y => n711);
   U223 : INVX1 port map( A => n380, Y => n710);
   U224 : NAND2X1 port map( A => n786, B => n190, Y => n108);
   U225 : INVX2 port map( A => n122, Y => n151);
   U226 : BUFX2 port map( A => n160, Y => n109);
   U227 : INVX1 port map( A => n66, Y => n110);
   U228 : INVX1 port map( A => n66, Y => n144);
   U229 : BUFX2 port map( A => n190, Y => n112);
   U230 : BUFX2 port map( A => n305, Y => n113);
   U231 : INVX1 port map( A => n507, Y => n114);
   U232 : AND2X2 port map( A => n305, B => n275, Y => n116);
   U233 : AND2X1 port map( A => n113, B => n275, Y => n171);
   U234 : NAND2X1 port map( A => n23, B => n629, Y => n117);
   U235 : NAND2X1 port map( A => n23, B => n629, Y => n118);
   U236 : INVX8 port map( A => n99, Y => n675);
   U237 : INVX1 port map( A => n428_port, Y => n744);
   U238 : AND2X1 port map( A => n303, B => si_5_port, Y => n304);
   U239 : INVX1 port map( A => n427_port, Y => n743);
   U240 : INVX2 port map( A => n1071, Y => n120);
   U241 : NOR2X1 port map( A => n194, B => n97, Y => n566);
   U242 : AND2X2 port map( A => n146, B => n1060, Y => n121);
   U243 : INVX1 port map( A => n121, Y => n1050);
   U244 : INVX4 port map( A => n125, Y => n608);
   U245 : NOR2X1 port map( A => n648, B => n684, Y => n123);
   U246 : AND2X2 port map( A => n224, B => n152, Y => n125);
   U247 : INVX1 port map( A => n187, Y => n127);
   U248 : INVX1 port map( A => n187, Y => n129);
   U249 : NOR2X1 port map( A => n197, B => n1045, Y => n161);
   U250 : AND2X2 port map( A => n434, B => n436, Y => n133);
   U251 : BUFX2 port map( A => n49, Y => n134);
   U252 : NAND2X1 port map( A => n439, B => n11, Y => nextProcessedData_7_port)
                           ;
   U253 : INVX1 port map( A => nextProcessedData_7_port, Y => n441);
   U254 : INVX1 port map( A => state_2_port, Y => n273);
   U255 : INVX8 port map( A => n136, Y => n137);
   U256 : INVX2 port map( A => state_1_port, Y => n139);
   U257 : NOR3X1 port map( A => n75, B => n156, C => n194, Y => n138);
   U258 : INVX4 port map( A => n193, Y => n194);
   U259 : NOR2X1 port map( A => n144, B => n76, Y => n140);
   U260 : AND2X2 port map( A => n683, B => n112, Y => n141);
   U261 : INVX4 port map( A => n141, Y => n149);
   U262 : BUFX2 port map( A => n154, Y => n148);
   U263 : NOR2X1 port map( A => n1135, B => n431_port, Y => n145);
   U264 : INVX1 port map( A => n145, Y => n387);
   U265 : AND2X2 port map( A => n487_port, B => n1074, Y => n146);
   U266 : INVX1 port map( A => n146, Y => n1085);
   U267 : INVX2 port map( A => n67, Y => n644);
   U268 : NAND2X1 port map( A => n167, B => n28, Y => n147);
   U269 : NOR2X1 port map( A => n27, B => n76, Y => n169);
   U270 : AND2X1 port map( A => n88, B => n1055, Y => n166);
   U271 : AND2X1 port map( A => keyi_2_port, B => keyi_1_port, Y => n172);
   U272 : INVX1 port map( A => n19, Y => n150);
   U273 : INVX2 port map( A => n205, Y => n202);
   U274 : INVX2 port map( A => n206, Y => n201);
   U275 : INVX2 port map( A => n207, Y => n200);
   U276 : BUFX2 port map( A => n154, Y => n198);
   U277 : INVX4 port map( A => n1027, Y => n1042);
   U278 : BUFX2 port map( A => n199, Y => n203);
   U279 : BUFX2 port map( A => n212, Y => n205);
   U280 : BUFX2 port map( A => n199, Y => n206);
   U281 : BUFX2 port map( A => n212, Y => n207);
   U282 : BUFX2 port map( A => n199, Y => n208);
   U283 : BUFX2 port map( A => n199, Y => n209);
   U284 : BUFX2 port map( A => n199, Y => n210);
   U285 : BUFX2 port map( A => n199, Y => n211);
   U286 : BUFX2 port map( A => n199, Y => n212);
   U287 : AND2X2 port map( A => n278, B => n1065, Y => n153);
   U288 : AND2X2 port map( A => n585, B => n1048, Y => n157);
   U289 : INVX2 port map( A => n1081, Y => n177);
   U290 : AND2X2 port map( A => n183, B => n140, Y => n160);
   U291 : AND2X2 port map( A => n1089, B => n236, Y => n162);
   U292 : INVX2 port map( A => RST, Y => n199);
   U293 : AND2X2 port map( A => n172, B => n512_port, Y => n164);
   U294 : AND2X2 port map( A => n189, B => n179, Y => n167);
   U295 : AND2X2 port map( A => n172, B => keyi_0_port, Y => n170);
   U296 : INVX1 port map( A => n405, Y => n721);
   U297 : INVX1 port map( A => n379, Y => n709);
   U298 : INVX4 port map( A => n242, Y => n1082);
   U299 : INVX1 port map( A => n189, Y => n1071);
   U300 : INVX4 port map( A => n197, Y => n237);
   U301 : NOR2X1 port map( A => n182, B => n184, Y => n175);
   U302 : AND2X2 port map( A => n175, B => n237, Y => n178);
   U303 : AND2X1 port map( A => n175, B => n237, Y => n180);
   U304 : INVX2 port map( A => n181, Y => n183);
   U305 : NAND2X1 port map( A => n188, B => n179, Y => n181);
   U306 : INVX1 port map( A => n147, Y => n224);
   U307 : INVX1 port map( A => n1074, Y => n1077);
   U308 : OR2X2 port map( A => n6, B => n1026, Y => n1027);
   U309 : INVX1 port map( A => n153, Y => n185);
   U310 : INVX1 port map( A => n681, Y => n268);
   U311 : INVX1 port map( A => n53, Y => n1075);
   U312 : INVX1 port map( A => n670, Y => n676);
   U313 : AND2X2 port map( A => n276, B => n681, Y => n187);
   U314 : INVX2 port map( A => state_3_port, Y => n188);
   U315 : AND2X2 port map( A => n239, B => n145, Y => n190);
   U316 : INVX1 port map( A => n112, Y => n401);
   U317 : AND2X2 port map( A => n152, B => n58, Y => n191);
   U318 : AND2X2 port map( A => n152, B => n58, Y => n192);
   U319 : INVX1 port map( A => n1065, Y => n269);
   U320 : AND2X1 port map( A => n1065, B => n208, Y => n680);
   U321 : INVX2 port map( A => n647, Y => n193);
   U322 : INVX4 port map( A => n1022, Y => n684);
   U323 : INVX2 port map( A => si_4_port, Y => n1104);
   U324 : INVX2 port map( A => si_5_port, Y => n1105);
   U325 : INVX2 port map( A => prefillCounter_5_port, Y => n1136);
   U326 : NAND3X1 port map( A => n167, B => n175, C => n237, Y => n1074);
   U327 : NAND3X1 port map( A => n111, B => n96, C => n223, Y => n213);
   U328 : NAND2X1 port map( A => n85, B => n167, Y => n487_port);
   U329 : INVX2 port map( A => n158, Y => n214);
   U330 : NAND2X1 port map( A => n1085, B => n214, Y => n219);
   U331 : NAND2X1 port map( A => n105, B => n64, Y => n232);
   U332 : NAND3X1 port map( A => n96, B => n184, C => n76, Y => n241);
   U333 : INVX2 port map( A => n241, Y => n215);
   U334 : OAI21X1 port map( A => n159, B => n1107, C => n215, Y => n216);
   U335 : OAI21X1 port map( A => n158, B => n150, C => n216, Y => n217);
   U336 : NAND2X1 port map( A => n134, B => n217, Y => n218);
   U337 : NAND2X1 port map( A => n219, B => n218, Y => n222);
   U338 : NOR2X1 port map( A => n220, B => n142, Y => n221);
   U339 : AOI21X1 port map( A => n1106, B => n222, C => n221, Y => n163);
   U340 : NAND2X1 port map( A => n160, B => n237, Y => n1090);
   U341 : NAND2X1 port map( A => n184, B => n182, Y => n1045);
   U342 : INVX2 port map( A => permuteComplete, Y => n1054);
   U343 : NAND2X1 port map( A => n167, B => n135, Y => n1048);
   U344 : AOI21X1 port map( A => n1046, B => n1054, C => n224, Y => n227);
   U345 : NAND2X1 port map( A => n160, B => n105, Y => n1089);
   U346 : XOR2X1 port map( A => n189, B => n96, Y => n225);
   U347 : NAND3X1 port map( A => n87, B => n225, C => n273, Y => n682);
   U348 : AND2X2 port map( A => n93, B => n36, Y => n226);
   U349 : NAND3X1 port map( A => n1090, B => n227, C => n226, Y => n1067);
   U350 : INVX2 port map( A => n1067, Y => n1101);
   U351 : NOR2X1 port map( A => prefillCounter_0_port, B => n168, Y => n228);
   U352 : NAND3X1 port map( A => n173, B => n645, C => n228, Y => n229);
   U353 : NAND3X1 port map( A => n49, B => n140, C => n105, Y => n436);
   U354 : NAND2X1 port map( A => n229, B => n436, Y => n231);
   U355 : NAND2X1 port map( A => n177, B => n72, Y => n670);
   U356 : NAND2X1 port map( A => n64, B => n237, Y => n244);
   U357 : NAND2X1 port map( A => n670, B => n34, Y => n230);
   U358 : NOR2X1 port map( A => n231, B => n230, Y => n165);
   U359 : NAND2X1 port map( A => n246, B => n49, Y => n434);
   U360 : AOI21X1 port map( A => n177, B => n26, C => n88, Y => n234);
   U361 : NAND2X1 port map( A => n241, B => n232, Y => n233);
   U362 : NAND2X1 port map( A => n49, B => n233, Y => n1060);
   U363 : NAND2X1 port map( A => n234, B => n121, Y => n431_port);
   U364 : NAND2X1 port map( A => n246, B => n1082, Y => n1070);
   U365 : OAI21X1 port map( A => n1081, B => n241, C => n1070, Y => n235);
   U366 : INVX2 port map( A => n235, Y => n585);
   U367 : AOI21X1 port map( A => n72, B => n1082, C => n62, Y => n236);
   U368 : NAND2X1 port map( A => n178, B => n183, Y => n276);
   U369 : NAND2X1 port map( A => n167, B => n32, Y => n278);
   U370 : AND2X2 port map( A => n276, B => n278, Y => n238);
   U371 : NAND3X1 port map( A => n162, B => n67, C => n238, Y => n398);
   U372 : NOR2X1 port map( A => n398, B => n98, Y => n239);
   U373 : OAI22X1 port map( A => n244, B => n243, C => n142, D => n241, Y => 
                           n245);
   U374 : NOR2X1 port map( A => n25, B => n245, Y => n646);
   U375 : NAND2X1 port map( A => n180, B => n49, Y => n681);
   U376 : NAND2X1 port map( A => n268, B => DATA_IN(7), Y => n248);
   U377 : NAND2X1 port map( A => n1082, B => n26, Y => n1022);
   U378 : NAND2X1 port map( A => prefillCounter_7_port, B => n684, Y => n282);
   U379 : AOI22X1 port map( A => extratemp_7_port, B => n269, C => n429_port, D
                           => temp_7_port, Y => n247);
   U380 : NAND3X1 port map( A => n248, B => n282, C => n247, Y => n249);
   U381 : AOI21X1 port map( A => n21, B => fdata_7_port, C => n249, Y => n691);
   U382 : NAND2X1 port map( A => n268, B => DATA_IN(6), Y => n251);
   U383 : NAND2X1 port map( A => prefillCounter_6_port, B => n684, Y => n295);
   U384 : AOI22X1 port map( A => extratemp_6_port, B => n269, C => n429_port, D
                           => temp_6_port, Y => n250);
   U385 : NAND3X1 port map( A => n251, B => n295, C => n250, Y => n252);
   U386 : AOI21X1 port map( A => n21, B => fdata_6_port, C => n252, Y => n693);
   U387 : NAND2X1 port map( A => n268, B => DATA_IN(5), Y => n254);
   U388 : NAND2X1 port map( A => n684, B => prefillCounter_5_port, Y => n309);
   U389 : AOI22X1 port map( A => extratemp_5_port, B => n269, C => n429_port, D
                           => temp_5_port, Y => n253);
   U390 : NAND3X1 port map( A => n254, B => n309, C => n253, Y => n255);
   U391 : AOI21X1 port map( A => n21, B => fdata_5_port, C => n255, Y => n694);
   U392 : NAND2X1 port map( A => n268, B => DATA_IN(4), Y => n257);
   U393 : NAND2X1 port map( A => prefillCounter_4_port, B => n684, Y => n321);
   U394 : AOI22X1 port map( A => extratemp_4_port, B => n269, C => n429_port, D
                           => temp_4_port, Y => n256);
   U395 : NAND3X1 port map( A => n257, B => n321, C => n256, Y => n258);
   U396 : AOI21X1 port map( A => n21, B => fdata_4_port, C => n258, Y => n695);
   U397 : NAND2X1 port map( A => n268, B => DATA_IN(3), Y => n260);
   U398 : NAND2X1 port map( A => prefillCounter_3_port, B => n684, Y => n334);
   U399 : AOI22X1 port map( A => extratemp_3_port, B => n269, C => n429_port, D
                           => temp_3_port, Y => n259);
   U400 : NAND3X1 port map( A => n260, B => n334, C => n259, Y => n261);
   U401 : AOI21X1 port map( A => n21, B => fdata_3_port, C => n261, Y => n696);
   U402 : NAND2X1 port map( A => n268, B => DATA_IN(2), Y => n263);
   U403 : NAND2X1 port map( A => prefillCounter_2_port, B => n684, Y => n347);
   U404 : AOI22X1 port map( A => extratemp_2_port, B => n269, C => n429_port, D
                           => temp_2_port, Y => n262);
   U405 : NAND3X1 port map( A => n263, B => n347, C => n262, Y => n264);
   U406 : AOI21X1 port map( A => n21, B => fdata_2_port, C => n264, Y => n697);
   U407 : NAND2X1 port map( A => n268, B => DATA_IN(1), Y => n266);
   U408 : NAND2X1 port map( A => prefillCounter_1_port, B => n684, Y => n360);
   U409 : AOI22X1 port map( A => extratemp_1_port, B => n269, C => n429_port, D
                           => temp_1_port, Y => n265);
   U410 : NAND3X1 port map( A => n266, B => n360, C => n265, Y => n267);
   U411 : AOI21X1 port map( A => n21, B => fdata_1_port, C => n267, Y => n698);
   U412 : NAND2X1 port map( A => n268, B => DATA_IN(0), Y => n271);
   U413 : NAND2X1 port map( A => prefillCounter_0_port, B => n684, Y => n371);
   U414 : AOI22X1 port map( A => extratemp_0_port, B => n269, C => n429_port, D
                           => temp_0_port, Y => n270);
   U415 : NAND3X1 port map( A => n271, B => n371, C => n270, Y => n272);
   U416 : AOI21X1 port map( A => n21, B => fdata_0_port, C => n272, Y => n699);
   U417 : NAND2X1 port map( A => n135, B => n273, Y => n388);
   U418 : NAND2X1 port map( A => n388, B => n274, Y => n367);
   U419 : OR2X2 port map( A => si_1_port, B => si_0_port, Y => n354);
   U420 : INVX2 port map( A => si_3_port, Y => n638);
   U421 : NAND2X1 port map( A => n59, B => n1104, Y => n303);
   U422 : INVX2 port map( A => n303, Y => n317);
   U423 : NAND2X1 port map( A => n317, B => n1105, Y => n290);
   U424 : INVX2 port map( A => n290, Y => n305);
   U425 : INVX2 port map( A => si_6_port, Y => n275);
   U426 : XOR2X1 port map( A => n116, B => si_7_port, Y => n277);
   U427 : AOI22X1 port map( A => sj_7_port, B => n367, C => n277, D => n127, Y 
                           => n287);
   U428 : AOI22X1 port map( A => N503, B => n644, C => intj_7_port, D => n53, Y
                           => n286);
   U429 : AND2X2 port map( A => faddr_7_port, B => n297, Y => n284);
   U430 : NAND2X1 port map( A => temp_7_port, B => n109, Y => n281);
   U431 : OAI21X1 port map( A => n87, B => n19, C => n1082, Y => n279);
   U432 : INVX2 port map( A => n279, Y => n373);
   U433 : NAND2X1 port map( A => n373, B => inti_7_port, Y => n280);
   U434 : NAND3X1 port map( A => n282, B => n281, C => n280, Y => n283);
   U435 : NOR2X1 port map( A => n284, B => n283, Y => n285);
   U436 : NAND3X1 port map( A => n287, B => n286, C => n285, Y => n288);
   U437 : INVX2 port map( A => n288, Y => n700);
   U438 : NAND2X1 port map( A => n54, B => n289, Y => n486_port);
   U439 : NAND2X1 port map( A => sj_6_port, B => n367, Y => n294);
   U440 : AND2X2 port map( A => si_6_port, B => n290, Y => n291);
   U441 : OAI21X1 port map( A => n171, B => n291, C => n127, Y => n293);
   U442 : AOI22X1 port map( A => intj_6_port, B => n53, C => N502, D => n644, Y
                           => n292);
   U443 : NAND3X1 port map( A => n294, B => n293, C => n292, Y => n302);
   U444 : NAND2X1 port map( A => temp_6_port, B => n109, Y => n296);
   U445 : NAND2X1 port map( A => n296, B => n295, Y => n301);
   U446 : INVX2 port map( A => faddr_6_port, Y => n299);
   U447 : NAND2X1 port map( A => n373, B => inti_6_port, Y => n298);
   U448 : OAI21X1 port map( A => n650, B => n299, C => n298, Y => n300);
   U449 : NOR3X1 port map( A => n302, B => n301, C => n300, Y => n702);
   U450 : NAND2X1 port map( A => sj_5_port, B => n367, Y => n308);
   U451 : OAI21X1 port map( A => n113, B => n304, C => n129, Y => n307);
   U452 : AOI22X1 port map( A => intj_5_port, B => n53, C => N501, D => n644, Y
                           => n306);
   U453 : NAND3X1 port map( A => n308, B => n307, C => n306, Y => n315);
   U454 : NAND2X1 port map( A => temp_5_port, B => n109, Y => n310);
   U455 : NAND2X1 port map( A => n310, B => n309, Y => n314);
   U456 : INVX2 port map( A => faddr_5_port, Y => n312);
   U457 : NAND2X1 port map( A => n373, B => inti_5_port, Y => n311);
   U458 : OAI21X1 port map( A => n650, B => n312, C => n311, Y => n313);
   U459 : NOR3X1 port map( A => n315, B => n314, C => n313, Y => n703);
   U460 : NAND2X1 port map( A => sj_4_port, B => n367, Y => n320);
   U461 : OAI21X1 port map( A => n317, B => n316, C => n127, Y => n319);
   U462 : AOI22X1 port map( A => intj_4_port, B => n53, C => N500, D => n644, Y
                           => n318);
   U463 : NAND3X1 port map( A => n320, B => n319, C => n318, Y => n327);
   U464 : NAND2X1 port map( A => temp_4_port, B => n109, Y => n322);
   U465 : NAND2X1 port map( A => n322, B => n321, Y => n326);
   U466 : INVX2 port map( A => faddr_4_port, Y => n324);
   U467 : NAND2X1 port map( A => n373, B => inti_4_port, Y => n323);
   U468 : OAI21X1 port map( A => n650, B => n324, C => n323, Y => n325);
   U469 : NOR3X1 port map( A => n327, B => n326, C => n325, Y => n704);
   U470 : NAND2X1 port map( A => sj_3_port, B => n367, Y => n333);
   U471 : NAND2X1 port map( A => si_3_port, B => n341, Y => n329);
   U472 : NAND2X1 port map( A => n329, B => n328, Y => n330);
   U473 : NAND2X1 port map( A => n330, B => n129, Y => n332);
   U474 : AOI22X1 port map( A => intj_3_port, B => n53, C => N499, D => n644, Y
                           => n331);
   U475 : NAND3X1 port map( A => n333, B => n332, C => n331, Y => n340);
   U476 : NAND2X1 port map( A => temp_3_port, B => n109, Y => n335);
   U477 : NAND2X1 port map( A => n335, B => n334, Y => n339);
   U478 : INVX2 port map( A => faddr_3_port, Y => n337);
   U479 : NAND2X1 port map( A => n373, B => inti_3_port, Y => n336);
   U480 : OAI21X1 port map( A => n650, B => n337, C => n336, Y => n338);
   U481 : NOR3X1 port map( A => n340, B => n339, C => n338, Y => n705);
   U482 : NAND2X1 port map( A => sj_2_port, B => n367, Y => n346);
   U483 : NAND2X1 port map( A => si_2_port, B => n354, Y => n342);
   U484 : NAND2X1 port map( A => n342, B => n341, Y => n343);
   U485 : NAND2X1 port map( A => n343, B => n127, Y => n345);
   U486 : AOI22X1 port map( A => intj_2_port, B => n53, C => N498, D => n644, Y
                           => n344);
   U487 : NAND3X1 port map( A => n346, B => n345, C => n344, Y => n353);
   U488 : NAND2X1 port map( A => temp_2_port, B => n109, Y => n348);
   U489 : NAND2X1 port map( A => n348, B => n347, Y => n352);
   U490 : INVX2 port map( A => faddr_2_port, Y => n350);
   U491 : NAND2X1 port map( A => n373, B => inti_2_port, Y => n349);
   U492 : OAI21X1 port map( A => n650, B => n350, C => n349, Y => n351);
   U493 : NOR3X1 port map( A => n353, B => n352, C => n351, Y => n706);
   U494 : NAND2X1 port map( A => sj_1_port, B => n367, Y => n359);
   U495 : NAND2X1 port map( A => n24, B => si_1_port, Y => n355);
   U496 : NAND2X1 port map( A => n355, B => n354, Y => n356);
   U497 : NAND2X1 port map( A => n356, B => n129, Y => n358);
   U498 : AOI22X1 port map( A => intj_1_port, B => n53, C => N497, D => n644, Y
                           => n357);
   U499 : NAND3X1 port map( A => n359, B => n358, C => n357, Y => n366);
   U500 : NAND2X1 port map( A => temp_1_port, B => n109, Y => n361);
   U501 : NAND2X1 port map( A => n361, B => n360, Y => n365);
   U502 : INVX2 port map( A => faddr_1_port, Y => n363);
   U503 : NAND2X1 port map( A => n373, B => inti_1_port, Y => n362);
   U504 : OAI21X1 port map( A => n650, B => n363, C => n362, Y => n364);
   U505 : NOR3X1 port map( A => n366, B => n365, C => n364, Y => n707);
   U506 : NAND2X1 port map( A => n48, B => n367, Y => n370);
   U507 : NAND2X1 port map( A => n129, B => n1102, Y => n369);
   U508 : AOI22X1 port map( A => intj_0_port, B => n53, C => N496, D => n644, Y
                           => n368);
   U509 : NAND3X1 port map( A => n370, B => n369, C => n368, Y => n378);
   U510 : NAND2X1 port map( A => temp_0_port, B => n109, Y => n372);
   U511 : NAND2X1 port map( A => n372, B => n371, Y => n377);
   U512 : INVX2 port map( A => faddr_0_port, Y => n375);
   U513 : NAND2X1 port map( A => n373, B => inti_0_port, Y => n374);
   U514 : OAI21X1 port map( A => n650, B => n375, C => n374, Y => n376);
   U515 : NOR3X1 port map( A => n378, B => n377, C => n376, Y => n708);
   U516 : NOR2X1 port map( A => n684, B => n52, Y => n391);
   U517 : INVX2 port map( A => n387, Y => n390);
   U518 : AND2X2 port map( A => n388, B => n30, Y => n389);
   U519 : NAND3X1 port map( A => n391, B => n390, C => n389, Y => n397);
   U520 : AOI21X1 port map( A => fr_enable, B => n397, C => n17, Y => n393);
   U521 : INVX2 port map( A => R_ENABLE_port, Y => n392);
   U522 : MUX2X1 port map( B => n393, A => n392, S => n202, Y => n717);
   U523 : AND2X2 port map( A => n681, B => n30, Y => n394);
   U524 : NAND3X1 port map( A => n36, B => n1022, C => n394, Y => n402);
   U525 : AOI21X1 port map( A => fw_enable, B => n401, C => n402, Y => n396);
   U526 : INVX2 port map( A => W_ENABLE_port, Y => n395);
   U527 : MUX2X1 port map( B => n396, A => n395, S => n202, Y => n718);
   U528 : OAI21X1 port map( A => n202, B => n397, C => fr_enable, Y => n400);
   U529 : NAND2X1 port map( A => n17, B => n207, Y => n399);
   U530 : NAND2X1 port map( A => n400, B => n399, Y => n719);
   U531 : OAI21X1 port map( A => n202, B => n401, C => fw_enable, Y => n404);
   U532 : NAND2X1 port map( A => n402, B => n206, Y => n403);
   U533 : NAND2X1 port map( A => n404, B => n403, Y => n720);
   U534 : MUX2X1 port map( B => nfaddr_0_port, A => ADDR_0_port, S => n201, Y 
                           => n413_port);
   U535 : INVX2 port map( A => n413_port, Y => n729);
   U536 : MUX2X1 port map( B => nfaddr_0_port, A => faddr_0_port, S => n201, Y 
                           => n414_port);
   U537 : INVX2 port map( A => n414_port, Y => n730);
   U538 : MUX2X1 port map( B => nfaddr_1_port, A => ADDR_1_port, S => n201, Y 
                           => n415);
   U539 : INVX2 port map( A => n415, Y => n731);
   U540 : MUX2X1 port map( B => nfaddr_1_port, A => faddr_1_port, S => n201, Y 
                           => n416);
   U541 : INVX2 port map( A => n416, Y => n732);
   U542 : MUX2X1 port map( B => nfaddr_2_port, A => ADDR_2_port, S => n201, Y 
                           => n417);
   U543 : INVX2 port map( A => n417, Y => n733);
   U544 : MUX2X1 port map( B => nfaddr_2_port, A => faddr_2_port, S => n201, Y 
                           => n418);
   U545 : INVX2 port map( A => n418, Y => n734);
   U546 : MUX2X1 port map( B => nfaddr_3_port, A => ADDR_3_port, S => n201, Y 
                           => n419);
   U547 : INVX2 port map( A => n419, Y => n735);
   U548 : MUX2X1 port map( B => nfaddr_3_port, A => faddr_3_port, S => n201, Y 
                           => n420);
   U549 : INVX2 port map( A => n420, Y => n736);
   U550 : MUX2X1 port map( B => nfaddr_4_port, A => ADDR_4_port, S => n201, Y 
                           => n421);
   U551 : INVX2 port map( A => n421, Y => n737);
   U552 : MUX2X1 port map( B => nfaddr_4_port, A => faddr_4_port, S => n201, Y 
                           => n422);
   U553 : INVX2 port map( A => n422, Y => n738);
   U554 : MUX2X1 port map( B => nfaddr_5_port, A => ADDR_5_port, S => n201, Y 
                           => n423);
   U555 : INVX2 port map( A => n423, Y => n739);
   U556 : MUX2X1 port map( B => nfaddr_5_port, A => faddr_5_port, S => n200, Y 
                           => n424_port);
   U557 : INVX2 port map( A => n424_port, Y => n740);
   U558 : MUX2X1 port map( B => nfaddr_6_port, A => ADDR_6_port, S => n200, Y 
                           => n425_port);
   U559 : INVX2 port map( A => n425_port, Y => n741);
   U560 : MUX2X1 port map( B => nfaddr_6_port, A => faddr_6_port, S => n200, Y 
                           => n426_port);
   U561 : INVX2 port map( A => n426_port, Y => n742);
   U562 : MUX2X1 port map( B => nfaddr_7_port, A => ADDR_7_port, S => n201, Y 
                           => n427_port);
   U563 : MUX2X1 port map( B => nfaddr_7_port, A => faddr_7_port, S => n200, Y 
                           => n428_port);
   U564 : NAND3X1 port map( A => n187, B => n162, C => n430_port, Y => n647);
   U565 : NOR2X1 port map( A => n194, B => n684, Y => n433);
   U566 : NAND2X1 port map( A => n103, B => currentProcessedData_7_port, Y => 
                           n439);
   U567 : XOR2X1 port map( A => delaydata_7_port, B => temp_7_port, Y => n435);
   U568 : NAND2X1 port map( A => n479_port, B => n435, Y => n438);
   U569 : NAND2X1 port map( A => BYTE(7), B => n480_port, Y => n437);
   U570 : INVX2 port map( A => PROCESSED_DATA_7_port, Y => n440);
   U571 : MUX2X1 port map( B => n441, A => n440, S => n200, Y => n745);
   U572 : NAND2X1 port map( A => n118, B => currentProcessedData_6_port, Y => 
                           n445);
   U573 : XOR2X1 port map( A => delaydata_6_port, B => temp_6_port, Y => n442);
   U574 : NAND2X1 port map( A => n479_port, B => n442, Y => n444);
   U575 : NAND2X1 port map( A => BYTE(6), B => n480_port, Y => n443);
   U576 : NAND3X1 port map( A => n445, B => n444, C => n443, Y => 
                           nextProcessedData_6_port);
   U577 : INVX2 port map( A => nextProcessedData_6_port, Y => n447);
   U578 : INVX2 port map( A => PROCESSED_DATA_6_port, Y => n446);
   U579 : MUX2X1 port map( B => n447, A => n446, S => n200, Y => n747);
   U580 : NAND2X1 port map( A => n117, B => currentProcessedData_5_port, Y => 
                           n451_port);
   U581 : XOR2X1 port map( A => delaydata_5_port, B => temp_5_port, Y => n448);
   U582 : NAND2X1 port map( A => n479_port, B => n448, Y => n450_port);
   U583 : NAND2X1 port map( A => BYTE(5), B => n480_port, Y => n449_port);
   U584 : NAND3X1 port map( A => n451_port, B => n450_port, C => n449_port, Y 
                           => nextProcessedData_5_port);
   U585 : INVX2 port map( A => nextProcessedData_5_port, Y => n453_port);
   U586 : INVX2 port map( A => PROCESSED_DATA_5_port, Y => n452_port);
   U587 : MUX2X1 port map( B => n453_port, A => n452_port, S => n200, Y => n749
                           );
   U588 : NAND2X1 port map( A => n103, B => currentProcessedData_4_port, Y => 
                           n457);
   U589 : XOR2X1 port map( A => delaydata_4_port, B => temp_4_port, Y => 
                           n454_port);
   U590 : NAND2X1 port map( A => n479_port, B => n454_port, Y => n456_port);
   U591 : NAND2X1 port map( A => BYTE(4), B => n480_port, Y => n455_port);
   U592 : NAND3X1 port map( A => n457, B => n456_port, C => n455_port, Y => 
                           nextProcessedData_4_port);
   U593 : INVX2 port map( A => nextProcessedData_4_port, Y => n459);
   U594 : INVX2 port map( A => PROCESSED_DATA_4_port, Y => n458);
   U595 : MUX2X1 port map( B => n459, A => n458, S => n200, Y => n751);
   U596 : NAND2X1 port map( A => n102, B => currentProcessedData_3_port, Y => 
                           n463);
   U597 : XOR2X1 port map( A => delaydata_3_port, B => temp_3_port, Y => n460);
   U598 : NAND2X1 port map( A => n479_port, B => n460, Y => n462);
   U599 : NAND2X1 port map( A => BYTE(3), B => n480_port, Y => n461);
   U600 : NAND3X1 port map( A => n463, B => n462, C => n461, Y => 
                           nextProcessedData_3_port);
   U601 : INVX2 port map( A => nextProcessedData_3_port, Y => n465);
   U602 : INVX2 port map( A => PROCESSED_DATA_3_port, Y => n464);
   U603 : MUX2X1 port map( B => n465, A => n464, S => n200, Y => n753);
   U604 : NAND2X1 port map( A => n118, B => currentProcessedData_2_port, Y => 
                           n469);
   U605 : XOR2X1 port map( A => delaydata_2_port, B => temp_2_port, Y => n466);
   U606 : NAND2X1 port map( A => n479_port, B => n466, Y => n468);
   U607 : NAND2X1 port map( A => BYTE(2), B => n480_port, Y => n467);
   U608 : NAND3X1 port map( A => n469, B => n468, C => n467, Y => 
                           nextProcessedData_2_port);
   U609 : INVX2 port map( A => nextProcessedData_2_port, Y => n471);
   U610 : INVX2 port map( A => PROCESSED_DATA_2_port, Y => n470);
   U611 : MUX2X1 port map( B => n471, A => n470, S => n200, Y => n755);
   U612 : NAND2X1 port map( A => n102, B => currentProcessedData_1_port, Y => 
                           n475_port);
   U613 : XOR2X1 port map( A => delaydata_1_port, B => temp_1_port, Y => 
                           n472_port);
   U614 : NAND2X1 port map( A => n479_port, B => n472_port, Y => n474_port);
   U615 : NAND2X1 port map( A => BYTE(1), B => n480_port, Y => n473_port);
   U616 : INVX2 port map( A => PROCESSED_DATA_1_port, Y => n476_port);
   U617 : MUX2X1 port map( B => n477_port, A => n476_port, S => n200, Y => n757
                           );
   U618 : NAND2X1 port map( A => n117, B => currentProcessedData_0_port, Y => 
                           n483_port);
   U619 : XOR2X1 port map( A => delaydata_0_port, B => temp_0_port, Y => 
                           n478_port);
   U620 : NAND2X1 port map( A => n479_port, B => n478_port, Y => n482_port);
   U621 : NAND2X1 port map( A => BYTE(0), B => n480_port, Y => n481_port);
   U622 : INVX2 port map( A => PROCESSED_DATA_0_port, Y => n484_port);
   U623 : MUX2X1 port map( B => n485_port, A => n484_port, S => n200, Y => n759
                           );
   U624 : NOR2X1 port map( A => n202, B => n104, Y => n489);
   U625 : NAND2X1 port map( A => n46, B => n1060, Y => n1073);
   U626 : INVX2 port map( A => n1073, Y => n488);
   U627 : NAND2X1 port map( A => n488, B => n133, Y => n564);
   U628 : NOR3X1 port map( A => n75, B => n156, C => n132, Y => n628);
   U629 : AND2X2 port map( A => n138, B => n489, Y => n507);
   U630 : INVX2 port map( A => N502, Y => n491);
   U631 : NAND3X1 port map( A => n560, B => n507, C => n563, Y => n504);
   U632 : NAND2X1 port map( A => inti_6_port, B => n504, Y => n490);
   U633 : OAI21X1 port map( A => n44, B => n491, C => n490, Y => n1125);
   U634 : INVX2 port map( A => N501, Y => n493);
   U635 : NAND2X1 port map( A => inti_5_port, B => n504, Y => n492);
   U636 : OAI21X1 port map( A => n44, B => n493, C => n492, Y => n1124);
   U637 : INVX2 port map( A => N500, Y => n495);
   U638 : NAND2X1 port map( A => inti_4_port, B => n504, Y => n494);
   U639 : OAI21X1 port map( A => n43, B => n495, C => n494, Y => n1123);
   U640 : INVX2 port map( A => N499, Y => n497_port);
   U641 : NAND2X1 port map( A => inti_3_port, B => n504, Y => n496_port);
   U642 : OAI21X1 port map( A => n33, B => n497_port, C => n496_port, Y => 
                           n1122);
   U643 : INVX2 port map( A => N498, Y => n499_port);
   U644 : NAND2X1 port map( A => inti_2_port, B => n504, Y => n498_port);
   U645 : OAI21X1 port map( A => n43, B => n499_port, C => n498_port, Y => 
                           n1121);
   U646 : INVX2 port map( A => N497, Y => n501_port);
   U647 : NAND2X1 port map( A => inti_1_port, B => n504, Y => n500_port);
   U648 : OAI21X1 port map( A => n44, B => n501_port, C => n500_port, Y => 
                           n1120);
   U649 : INVX2 port map( A => N496, Y => n503_port);
   U650 : NAND2X1 port map( A => inti_0_port, B => n504, Y => n502_port);
   U651 : OAI21X1 port map( A => n43, B => n503_port, C => n502_port, Y => 
                           n1119);
   U652 : INVX2 port map( A => N503, Y => n506);
   U653 : NAND2X1 port map( A => inti_7_port, B => n504, Y => n505);
   U654 : OAI21X1 port map( A => n33, B => n506, C => n505, Y => n1126);
   U655 : NAND3X1 port map( A => keyi_2_port, B => n510, C => n512_port, Y => 
                           n508);
   U656 : INVX2 port map( A => n508, Y => n550);
   U657 : NAND3X1 port map( A => keyi_2_port, B => keyi_0_port, C => n510, Y =>
                           n509);
   U658 : INVX2 port map( A => n509, Y => n549);
   U659 : AOI22X1 port map( A => keyTable_4_7_port, B => n550, C => 
                           keyTable_5_7_port, D => n549, Y => n518_port);
   U660 : AOI22X1 port map( A => keyTable_6_7_port, B => n164, C => 
                           keyTable_7_7_port, D => n170, Y => n517_port);
   U661 : INVX2 port map( A => keyTable_3_7_port, Y => n943);
   U662 : NAND3X1 port map( A => keyi_1_port, B => n511, C => n512_port, Y => 
                           n551);
   U663 : INVX2 port map( A => keyTable_2_7_port, Y => n927);
   U664 : OAI22X1 port map( A => n552, B => n943, C => n551, D => n927, Y => 
                           n515_port);
   U665 : NAND3X1 port map( A => keyi_0_port, B => n511, C => n510, Y => n554);
   U666 : INVX2 port map( A => keyTable_1_7_port, Y => n790);
   U667 : NOR2X1 port map( A => keyi_2_port, B => keyi_1_port, Y => n513_port);
   U668 : NAND2X1 port map( A => n513_port, B => n512_port, Y => n553);
   U670 : INVX2 port map( A => keyTable_0_7_port, Y => n788);
   U671 : OAI22X1 port map( A => n554, B => n790, C => n553, D => n788, Y => 
                           n514_port);
   U672 : NOR2X1 port map( A => n515_port, B => n514_port, Y => n516_port);
   U674 : NAND3X1 port map( A => n518_port, B => n517_port, C => n516_port, Y 
                           => N472);
   U675 : AOI22X1 port map( A => keyTable_4_6_port, B => n550, C => 
                           keyTable_5_6_port, D => n549, Y => n523_port);
   U676 : AOI22X1 port map( A => keyTable_6_6_port, B => n164, C => 
                           keyTable_7_6_port, D => n170, Y => n522_port);
   U677 : INVX2 port map( A => keyTable_3_6_port, Y => n945);
   U678 : INVX2 port map( A => keyTable_2_6_port, Y => n929);
   U679 : OAI22X1 port map( A => n552, B => n945, C => n551, D => n929, Y => 
                           n520_port);
   U680 : INVX2 port map( A => keyTable_1_6_port, Y => n889);
   U681 : INVX2 port map( A => keyTable_0_6_port, Y => n887);
   U682 : OAI22X1 port map( A => n554, B => n889, C => n553, D => n887, Y => 
                           n519_port);
   U683 : NOR2X1 port map( A => n520_port, B => n519_port, Y => n521_port);
   U684 : NAND3X1 port map( A => n523_port, B => n522_port, C => n521_port, Y 
                           => N473);
   U685 : AOI22X1 port map( A => keyTable_4_5_port, B => n550, C => 
                           keyTable_5_5_port, D => n549, Y => n528);
   U686 : AOI22X1 port map( A => keyTable_6_5_port, B => n164, C => 
                           keyTable_7_5_port, D => n170, Y => n527_port);
   U687 : INVX2 port map( A => keyTable_3_5_port, Y => n947);
   U688 : INVX2 port map( A => keyTable_2_5_port, Y => n931);
   U689 : OAI22X1 port map( A => n552, B => n947, C => n551, D => n931, Y => 
                           n525_port);
   U690 : INVX2 port map( A => keyTable_1_5_port, Y => n898);
   U691 : INVX2 port map( A => keyTable_0_5_port, Y => n885);
   U692 : OAI22X1 port map( A => n554, B => n898, C => n553, D => n885, Y => 
                           n524_port);
   U693 : NOR2X1 port map( A => n525_port, B => n524_port, Y => n526_port);
   U694 : NAND3X1 port map( A => n528, B => n527_port, C => n526_port, Y => 
                           N474);
   U695 : AOI22X1 port map( A => keyTable_4_4_port, B => n550, C => 
                           keyTable_5_4_port, D => n549, Y => n533);
   U696 : AOI22X1 port map( A => keyTable_6_4_port, B => n164, C => 
                           keyTable_7_4_port, D => n170, Y => n532);
   U697 : INVX2 port map( A => keyTable_3_4_port, Y => n949);
   U698 : INVX2 port map( A => keyTable_2_4_port, Y => n933);
   U699 : OAI22X1 port map( A => n552, B => n949, C => n551, D => n933, Y => 
                           n530);
   U700 : INVX2 port map( A => keyTable_1_4_port, Y => n917);
   U701 : INVX2 port map( A => keyTable_0_4_port, Y => n883);
   U702 : OAI22X1 port map( A => n554, B => n917, C => n553, D => n883, Y => 
                           n529);
   U703 : NOR2X1 port map( A => n530, B => n529, Y => n531);
   U704 : NAND3X1 port map( A => n533, B => n532, C => n531, Y => N475);
   U705 : AOI22X1 port map( A => keyTable_4_3_port, B => n550, C => 
                           keyTable_5_3_port, D => n549, Y => n538);
   U706 : AOI22X1 port map( A => keyTable_6_3_port, B => n164, C => 
                           keyTable_7_3_port, D => n170, Y => n537);
   U707 : INVX2 port map( A => keyTable_3_3_port, Y => n951);
   U708 : INVX2 port map( A => keyTable_2_3_port, Y => n935);
   U709 : OAI22X1 port map( A => n552, B => n951, C => n551, D => n935, Y => 
                           n535);
   U710 : INVX2 port map( A => keyTable_1_3_port, Y => n919);
   U711 : INVX2 port map( A => keyTable_0_3_port, Y => n870);
   U712 : OAI22X1 port map( A => n554, B => n919, C => n553, D => n870, Y => 
                           n534);
   U713 : NOR2X1 port map( A => n535, B => n534, Y => n536);
   U714 : NAND3X1 port map( A => n538, B => n537, C => n536, Y => N476);
   U715 : AOI22X1 port map( A => keyTable_4_2_port, B => n550, C => 
                           keyTable_5_2_port, D => n549, Y => n543);
   U716 : AOI22X1 port map( A => keyTable_6_2_port, B => n164, C => 
                           keyTable_7_2_port, D => n170, Y => n542);
   U717 : INVX2 port map( A => keyTable_3_2_port, Y => n953);
   U718 : INVX2 port map( A => keyTable_2_2_port, Y => n937);
   U719 : OAI22X1 port map( A => n552, B => n953, C => n551, D => n937, Y => 
                           n540);
   U720 : INVX2 port map( A => keyTable_1_2_port, Y => n921);
   U721 : INVX2 port map( A => keyTable_0_2_port, Y => n868);
   U722 : OAI22X1 port map( A => n554, B => n921, C => n553, D => n868, Y => 
                           n539);
   U723 : NOR2X1 port map( A => n540, B => n539, Y => n541);
   U724 : NAND3X1 port map( A => n543, B => n542, C => n541, Y => N477);
   U725 : AOI22X1 port map( A => keyTable_4_1_port, B => n550, C => 
                           keyTable_5_1_port, D => n549, Y => n548);
   U726 : AOI22X1 port map( A => keyTable_6_1_port, B => n164, C => 
                           keyTable_7_1_port, D => n170, Y => n547);
   U727 : INVX2 port map( A => keyTable_3_1_port, Y => n955);
   U728 : INVX2 port map( A => keyTable_2_1_port, Y => n939);
   U729 : OAI22X1 port map( A => n552, B => n955, C => n551, D => n939, Y => 
                           n545);
   U730 : INVX2 port map( A => keyTable_1_1_port, Y => n923);
   U731 : INVX2 port map( A => keyTable_0_1_port, Y => n866);
   U732 : OAI22X1 port map( A => n554, B => n923, C => n553, D => n866, Y => 
                           n544);
   U733 : NOR2X1 port map( A => n545, B => n544, Y => n546);
   U734 : NAND3X1 port map( A => n548, B => n547, C => n546, Y => N478);
   U735 : AOI22X1 port map( A => keyTable_4_0_port, B => n550, C => 
                           keyTable_5_0_port, D => n549, Y => n559);
   U736 : AOI22X1 port map( A => keyTable_6_0_port, B => n164, C => 
                           keyTable_7_0_port, D => n170, Y => n558);
   U737 : INVX2 port map( A => keyTable_3_0_port, Y => n957);
   U738 : INVX2 port map( A => keyTable_2_0_port, Y => n941);
   U739 : OAI22X1 port map( A => n552, B => n957, C => n551, D => n941, Y => 
                           n556);
   U740 : INVX2 port map( A => keyTable_1_0_port, Y => n925);
   U741 : INVX2 port map( A => keyTable_0_0_port, Y => n864);
   U742 : OAI22X1 port map( A => n554, B => n925, C => n553, D => n864, Y => 
                           n555);
   U743 : NOR2X1 port map( A => n556, B => n555, Y => n557);
   U744 : NAND3X1 port map( A => n559, B => n558, C => n557, Y => N479);
   U745 : NAND3X1 port map( A => n560, B => n7, C => n70, Y => n561);
   U746 : AND2X2 port map( A => n566, B => n22, Y => n590);
   U747 : NAND2X1 port map( A => n590, B => n54, Y => n582);
   U748 : INVX2 port map( A => n582, Y => n573);
   U749 : INVX2 port map( A => n48, Y => n568);
   U750 : INVX2 port map( A => n1090, Y => n587);
   U751 : NAND2X1 port map( A => N480, B => n587, Y => n567);
   U752 : OAI21X1 port map( A => n573, B => n568, C => n567, Y => n891);
   U753 : INVX2 port map( A => sj_1_port, Y => n570);
   U754 : NAND2X1 port map( A => N481, B => n587, Y => n569);
   U755 : OAI21X1 port map( A => n573, B => n570, C => n569, Y => n892);
   U756 : NAND2X1 port map( A => N482, B => n587, Y => n571);
   U757 : OAI21X1 port map( A => n573, B => n572, C => n571, Y => n893);
   U758 : NAND2X1 port map( A => sj_3_port, B => n582, Y => n575);
   U759 : NAND2X1 port map( A => N483, B => n587, Y => n574);
   U760 : NAND2X1 port map( A => n575, B => n574, Y => n894);
   U761 : NAND2X1 port map( A => sj_4_port, B => n582, Y => n577);
   U762 : NAND2X1 port map( A => N484, B => n587, Y => n576);
   U763 : NAND2X1 port map( A => n577, B => n576, Y => n895);
   U764 : NAND2X1 port map( A => sj_5_port, B => n582, Y => n579);
   U765 : NAND2X1 port map( A => N485, B => n587, Y => n578);
   U766 : NAND2X1 port map( A => n579, B => n578, Y => n896);
   U767 : NAND2X1 port map( A => sj_6_port, B => n582, Y => n581);
   U768 : NAND2X1 port map( A => N486, B => n587, Y => n580);
   U769 : NAND2X1 port map( A => n581, B => n580, Y => n897);
   U770 : NAND2X1 port map( A => sj_7_port, B => n582, Y => n584);
   U771 : INVX2 port map( A => N487, Y => n583);
   U772 : AOI22X1 port map( A => n584, B => n1090, C => n584, D => n583, Y => 
                           n1099);
   U773 : NAND2X1 port map( A => n106, B => n205, Y => n586);
   U774 : NOR2X1 port map( A => n587, B => n586, Y => n591);
   U775 : INVX2 port map( A => N518, Y => n593);
   U776 : NAND2X1 port map( A => intj_6_port, B => n55, Y => n592);
   U777 : OAI21X1 port map( A => n608, B => n593, C => n592, Y => n876);
   U778 : INVX2 port map( A => N517, Y => n595);
   U779 : NAND2X1 port map( A => intj_5_port, B => n55, Y => n594);
   U780 : OAI21X1 port map( A => n608, B => n595, C => n594, Y => n877);
   U781 : INVX2 port map( A => N516, Y => n597);
   U782 : NAND2X1 port map( A => intj_4_port, B => n55, Y => n596);
   U783 : OAI21X1 port map( A => n608, B => n597, C => n596, Y => n878);
   U784 : INVX2 port map( A => N515, Y => n599);
   U785 : NAND2X1 port map( A => intj_3_port, B => n55, Y => n598);
   U786 : OAI21X1 port map( A => n608, B => n599, C => n598, Y => n879);
   U787 : INVX2 port map( A => N514, Y => n601);
   U788 : NAND2X1 port map( A => intj_2_port, B => n55, Y => n600);
   U789 : OAI21X1 port map( A => n608, B => n601, C => n600, Y => n880);
   U790 : INVX2 port map( A => N513, Y => n603);
   U791 : NAND2X1 port map( A => intj_1_port, B => n55, Y => n602);
   U792 : OAI21X1 port map( A => n608, B => n603, C => n602, Y => n881);
   U793 : INVX2 port map( A => N512, Y => n605);
   U794 : NAND2X1 port map( A => intj_0_port, B => n55, Y => n604);
   U795 : OAI21X1 port map( A => n608, B => n605, C => n604, Y => n882);
   U796 : INVX2 port map( A => N519, Y => n607);
   U797 : NAND2X1 port map( A => intj_7_port, B => n55, Y => n606);
   U798 : OAI21X1 port map( A => n608, B => n607, C => n606, Y => n875);
   U799 : INVX2 port map( A => delaydata_6_port, Y => n610);
   U800 : INVX2 port map( A => BYTE(6), Y => n609);
   U801 : MUX2X1 port map( B => n610, A => n609, S => n191, Y => n1112);
   U802 : INVX2 port map( A => delaydata_5_port, Y => n612);
   U803 : INVX2 port map( A => BYTE(5), Y => n611);
   U804 : MUX2X1 port map( B => n612, A => n611, S => n192, Y => n1113);
   U805 : INVX2 port map( A => delaydata_4_port, Y => n614);
   U806 : INVX2 port map( A => BYTE(4), Y => n613);
   U807 : MUX2X1 port map( B => n614, A => n613, S => n191, Y => n1114);
   U808 : INVX2 port map( A => delaydata_3_port, Y => n616);
   U809 : INVX2 port map( A => BYTE(3), Y => n615);
   U810 : MUX2X1 port map( B => n616, A => n615, S => n192, Y => n1115);
   U811 : INVX2 port map( A => delaydata_2_port, Y => n618);
   U812 : INVX2 port map( A => BYTE(2), Y => n617);
   U813 : MUX2X1 port map( B => n618, A => n617, S => n191, Y => n1116);
   U814 : INVX2 port map( A => delaydata_1_port, Y => n620);
   U815 : INVX2 port map( A => BYTE(1), Y => n619);
   U816 : MUX2X1 port map( B => n620, A => n619, S => n192, Y => n1117);
   U817 : INVX2 port map( A => delaydata_0_port, Y => n622);
   U818 : INVX2 port map( A => BYTE(0), Y => n621);
   U819 : MUX2X1 port map( B => n622, A => n621, S => n191, Y => n1118);
   U820 : INVX2 port map( A => delaydata_7_port, Y => n624);
   U821 : INVX2 port map( A => BYTE(7), Y => n623);
   U822 : MUX2X1 port map( B => n624, A => n623, S => n192, Y => n1111);
   U823 : NAND3X1 port map( A => si_3_port, B => si_2_port, C => si_6_port, Y 
                           => n626);
   U824 : NAND2X1 port map( A => n588, B => si_7_port, Y => n625);
   U825 : NOR2X1 port map( A => n626, B => n625, Y => n627);
   U826 : NAND2X1 port map( A => n627, B => n589, Y => n1055);
   U827 : NAND2X1 port map( A => N431, B => n166, Y => n631);
   U828 : NAND2X1 port map( A => n629, B => n628, Y => n634);
   U829 : NAND2X1 port map( A => si_7_port, B => n634, Y => n630);
   U830 : NAND2X1 port map( A => n631, B => n630, Y => n900);
   U831 : NAND2X1 port map( A => N430, B => n166, Y => n633);
   U832 : NAND2X1 port map( A => si_6_port, B => n634, Y => n632);
   U833 : NAND2X1 port map( A => n633, B => n632, Y => n901);
   U834 : INVX2 port map( A => n634, Y => n643);
   U835 : NAND2X1 port map( A => N429, B => n166, Y => n635);
   U836 : OAI21X1 port map( A => n1105, B => n643, C => n635, Y => n902);
   U837 : NAND2X1 port map( A => N428, B => n166, Y => n636);
   U838 : OAI21X1 port map( A => n1104, B => n643, C => n636, Y => n903);
   U839 : NAND2X1 port map( A => N427, B => n166, Y => n637);
   U840 : OAI21X1 port map( A => n643, B => n638, C => n637, Y => n904);
   U841 : NAND2X1 port map( A => N426, B => n166, Y => n639);
   U842 : OAI21X1 port map( A => n643, B => n640, C => n639, Y => n905);
   U843 : NAND2X1 port map( A => N425, B => n166, Y => n641);
   U844 : OAI21X1 port map( A => n1103, B => n643, C => n641, Y => n906);
   U845 : NAND2X1 port map( A => N424, B => n166, Y => n642);
   U846 : OAI21X1 port map( A => n1102, B => n643, C => n642, Y => n907);
   U847 : NOR2X1 port map( A => n645, B => n644, Y => n651);
   U848 : NAND2X1 port map( A => n91, B => n203, Y => n648);
   U849 : NAND3X1 port map( A => n651, B => n71, C => n649, Y => n674);
   U850 : NAND2X1 port map( A => temp_6_port, B => n196, Y => n654);
   U851 : NAND3X1 port map( A => DATA_IN(6), B => n3, C => n675, Y => n653);
   U852 : NAND3X1 port map( A => N526, B => n676, C => n675, Y => n652);
   U853 : NAND3X1 port map( A => n654, B => n652, C => n653, Y => n857);
   U854 : NAND2X1 port map( A => temp_5_port, B => n196, Y => n657);
   U855 : NAND3X1 port map( A => DATA_IN(5), B => n3, C => n675, Y => n656);
   U856 : NAND3X1 port map( A => N525, B => n676, C => n675, Y => n655);
   U857 : NAND3X1 port map( A => n657, B => n655, C => n656, Y => n858);
   U858 : NAND2X1 port map( A => temp_4_port, B => n196, Y => n660);
   U859 : NAND3X1 port map( A => DATA_IN(4), B => n3, C => n675, Y => n659);
   U860 : NAND3X1 port map( A => N524, B => n676, C => n675, Y => n658);
   U861 : NAND3X1 port map( A => n660, B => n658, C => n659, Y => n859);
   U862 : NAND2X1 port map( A => temp_3_port, B => n196, Y => n663);
   U863 : NAND3X1 port map( A => DATA_IN(3), B => n3, C => n675, Y => n662);
   U864 : NAND3X1 port map( A => N523, B => n676, C => n151, Y => n661);
   U865 : NAND3X1 port map( A => n663, B => n661, C => n662, Y => n860);
   U866 : NAND2X1 port map( A => temp_2_port, B => n196, Y => n666);
   U867 : NAND3X1 port map( A => DATA_IN(2), B => n3, C => n675, Y => n665);
   U868 : NAND3X1 port map( A => N522, B => n676, C => n151, Y => n664);
   U869 : NAND3X1 port map( A => n666, B => n664, C => n665, Y => n861);
   U870 : NAND2X1 port map( A => temp_1_port, B => n196, Y => n669);
   U871 : NAND3X1 port map( A => DATA_IN(1), B => n3, C => n675, Y => n668);
   U872 : NAND3X1 port map( A => N521, B => n676, C => n675, Y => n667);
   U873 : NAND3X1 port map( A => n669, B => n667, C => n668, Y => n862);
   U874 : NAND2X1 port map( A => temp_0_port, B => n196, Y => n673);
   U875 : NAND3X1 port map( A => DATA_IN(0), B => n3, C => n151, Y => n672);
   U876 : NAND3X1 port map( A => N520, B => n676, C => n675, Y => n671);
   U877 : NAND3X1 port map( A => n673, B => n672, C => n671, Y => n863);
   U878 : NAND2X1 port map( A => temp_7_port, B => n196, Y => n679);
   U879 : NAND3X1 port map( A => DATA_IN(7), B => n3, C => n675, Y => n678);
   U880 : NAND3X1 port map( A => N527, B => n676, C => n151, Y => n677);
   U881 : NAND3X1 port map( A => n679, B => n677, C => n678, Y => n856);
   U882 : NAND3X1 port map( A => n682, B => n60, C => n57, Y => n785);
   U883 : NAND2X1 port map( A => n684, B => n141, Y => n1098);
   U884 : INVX2 port map( A => N413, Y => n686);
   U885 : NAND2X1 port map( A => prefillCounter_6_port, B => n149, Y => n685);
   U886 : OAI21X1 port map( A => n68, B => n686, C => n685, Y => n908);
   U887 : INVX2 port map( A => N412, Y => n688);
   U888 : NAND2X1 port map( A => n149, B => prefillCounter_5_port, Y => n687);
   U889 : OAI21X1 port map( A => n68, B => n688, C => n687, Y => n909);
   U890 : INVX2 port map( A => N411, Y => n690);
   U891 : NAND2X1 port map( A => prefillCounter_4_port, B => n149, Y => n689);
   U892 : OAI21X1 port map( A => n68, B => n690, C => n689, Y => n910);
   U893 : INVX2 port map( A => N410, Y => n701);
   U894 : NAND2X1 port map( A => prefillCounter_3_port, B => n149, Y => n692);
   U895 : OAI21X1 port map( A => n68, B => n701, C => n692, Y => n911);
   U896 : INVX2 port map( A => N409, Y => n766);
   U897 : NAND2X1 port map( A => prefillCounter_2_port, B => n149, Y => n765);
   U898 : OAI21X1 port map( A => n1098, B => n766, C => n765, Y => n912);
   U899 : INVX2 port map( A => N408, Y => n770);
   U900 : NAND2X1 port map( A => prefillCounter_1_port, B => n149, Y => n769);
   U901 : OAI21X1 port map( A => n1098, B => n770, C => n769, Y => n913);
   U914 : INVX2 port map( A => N414, Y => n784);
   U915 : NAND2X1 port map( A => prefillCounter_7_port, B => n149, Y => n783);
   U918 : OAI21X1 port map( A => n1098, B => n784, C => n783, Y => n914);
   U919 : INVX2 port map( A => KEY(7), Y => n787);
   U932 : NOR2X1 port map( A => n47, B => n785, Y => n786);
   U933 : MUX2X1 port map( B => n788, A => n787, S => n137, Y => n855);
   U934 : INVX2 port map( A => KEY(15), Y => n789);
   U935 : MUX2X1 port map( B => n790, A => n789, S => n78, Y => n854);
   U936 : INVX2 port map( A => KEY(0), Y => n791);
   U937 : MUX2X1 port map( B => n864, A => n791, S => n137, Y => n853);
   U938 : INVX2 port map( A => KEY(1), Y => n865);
   U939 : MUX2X1 port map( B => n866, A => n865, S => n82, Y => n852);
   U940 : INVX2 port map( A => KEY(2), Y => n867);
   U941 : MUX2X1 port map( B => n868, A => n867, S => n80, Y => n851);
   U942 : INVX2 port map( A => KEY(3), Y => n869);
   U943 : MUX2X1 port map( B => n870, A => n869, S => n137, Y => n850);
   U944 : INVX2 port map( A => KEY(4), Y => n871);
   U945 : MUX2X1 port map( B => n883, A => n871, S => n137, Y => n849);
   U946 : INVX2 port map( A => KEY(5), Y => n884);
   U947 : MUX2X1 port map( B => n885, A => n884, S => n137, Y => n848);
   U948 : INVX2 port map( A => KEY(6), Y => n886);
   U949 : MUX2X1 port map( B => n887, A => n886, S => n137, Y => n847);
   U950 : INVX2 port map( A => KEY(14), Y => n888);
   U951 : MUX2X1 port map( B => n889, A => n888, S => n78, Y => n846);
   U952 : INVX2 port map( A => KEY(13), Y => n890);
   U953 : MUX2X1 port map( B => n898, A => n890, S => n137, Y => n845);
   U954 : INVX2 port map( A => KEY(12), Y => n916);
   U955 : MUX2X1 port map( B => n917, A => n916, S => n77, Y => n844);
   U956 : INVX2 port map( A => KEY(11), Y => n918);
   U957 : MUX2X1 port map( B => n919, A => n918, S => n77, Y => n843);
   U958 : INVX2 port map( A => KEY(10), Y => n920);
   U959 : MUX2X1 port map( B => n921, A => n920, S => n77, Y => n842);
   U960 : INVX2 port map( A => KEY(9), Y => n922);
   U961 : MUX2X1 port map( B => n923, A => n922, S => n78, Y => n841);
   U962 : INVX2 port map( A => KEY(8), Y => n924);
   U963 : MUX2X1 port map( B => n925, A => n924, S => n78, Y => n840);
   U964 : INVX2 port map( A => KEY(23), Y => n926);
   U965 : MUX2X1 port map( B => n927, A => n926, S => n80, Y => n839);
   U966 : INVX2 port map( A => KEY(22), Y => n928);
   U967 : MUX2X1 port map( B => n929, A => n928, S => n143, Y => n838);
   U968 : INVX2 port map( A => KEY(21), Y => n930);
   U969 : MUX2X1 port map( B => n931, A => n930, S => n137, Y => n837);
   U970 : INVX2 port map( A => KEY(20), Y => n932);
   U971 : MUX2X1 port map( B => n933, A => n932, S => n137, Y => n836);
   U972 : INVX2 port map( A => KEY(19), Y => n934);
   U973 : MUX2X1 port map( B => n935, A => n934, S => n137, Y => n835);
   U974 : INVX2 port map( A => KEY(18), Y => n936);
   U975 : MUX2X1 port map( B => n937, A => n936, S => n143, Y => n834);
   U976 : INVX2 port map( A => KEY(17), Y => n938);
   U977 : MUX2X1 port map( B => n939, A => n938, S => n82, Y => n833);
   U978 : INVX2 port map( A => KEY(16), Y => n940);
   U979 : MUX2X1 port map( B => n941, A => n940, S => n137, Y => n832);
   U980 : INVX2 port map( A => KEY(31), Y => n942);
   U981 : MUX2X1 port map( B => n943, A => n942, S => n80, Y => n831);
   U982 : INVX2 port map( A => KEY(30), Y => n944);
   U983 : MUX2X1 port map( B => n945, A => n944, S => n82, Y => n830);
   U984 : INVX2 port map( A => KEY(29), Y => n946);
   U985 : MUX2X1 port map( B => n947, A => n946, S => n82, Y => n829);
   U986 : INVX2 port map( A => KEY(28), Y => n948);
   U987 : MUX2X1 port map( B => n949, A => n948, S => n80, Y => n828);
   U988 : INVX2 port map( A => KEY(27), Y => n950);
   U989 : MUX2X1 port map( B => n951, A => n950, S => n137, Y => n827);
   U990 : INVX2 port map( A => KEY(26), Y => n952);
   U991 : MUX2X1 port map( B => n953, A => n952, S => n143, Y => n826);
   U992 : INVX2 port map( A => KEY(25), Y => n954);
   U993 : MUX2X1 port map( B => n955, A => n954, S => n137, Y => n825);
   U994 : INVX2 port map( A => KEY(24), Y => n956);
   U995 : MUX2X1 port map( B => n957, A => n956, S => n143, Y => n824);
   U996 : INVX2 port map( A => keyTable_4_7_port, Y => n959);
   U997 : INVX2 port map( A => KEY(39), Y => n958);
   U998 : MUX2X1 port map( B => n959, A => n958, S => n137, Y => n823);
   U999 : INVX2 port map( A => keyTable_4_6_port, Y => n961);
   U1000 : INVX2 port map( A => KEY(38), Y => n960);
   U1001 : MUX2X1 port map( B => n961, A => n960, S => n77, Y => n822);
   U1002 : INVX2 port map( A => keyTable_4_5_port, Y => n963);
   U1003 : INVX2 port map( A => KEY(37), Y => n962);
   U1004 : MUX2X1 port map( B => n963, A => n962, S => n78, Y => n821);
   U1005 : INVX2 port map( A => keyTable_4_4_port, Y => n965);
   U1006 : INVX2 port map( A => KEY(36), Y => n964);
   U1007 : MUX2X1 port map( B => n965, A => n964, S => n78, Y => n820);
   U1008 : INVX2 port map( A => keyTable_4_3_port, Y => n967);
   U1009 : INVX2 port map( A => KEY(35), Y => n966);
   U1010 : MUX2X1 port map( B => n967, A => n966, S => n78, Y => n819);
   U1011 : INVX2 port map( A => keyTable_4_2_port, Y => n969);
   U1012 : INVX2 port map( A => KEY(34), Y => n968);
   U1013 : MUX2X1 port map( B => n969, A => n968, S => n80, Y => n818);
   U1014 : INVX2 port map( A => keyTable_4_1_port, Y => n971);
   U1015 : INVX2 port map( A => KEY(33), Y => n970);
   U1016 : MUX2X1 port map( B => n971, A => n970, S => n78, Y => n817);
   U1017 : INVX2 port map( A => keyTable_4_0_port, Y => n973);
   U1018 : INVX2 port map( A => KEY(32), Y => n972);
   U1019 : MUX2X1 port map( B => n973, A => n972, S => n77, Y => n816);
   U1020 : INVX2 port map( A => keyTable_5_7_port, Y => n975);
   U1021 : INVX2 port map( A => KEY(47), Y => n974);
   U1022 : MUX2X1 port map( B => n975, A => n974, S => n143, Y => n815);
   U1023 : INVX2 port map( A => keyTable_5_6_port, Y => n977);
   U1024 : INVX2 port map( A => KEY(46), Y => n976);
   U1025 : MUX2X1 port map( B => n977, A => n976, S => n143, Y => n814);
   U1026 : INVX2 port map( A => keyTable_5_5_port, Y => n979);
   U1027 : INVX2 port map( A => KEY(45), Y => n978);
   U1028 : MUX2X1 port map( B => n979, A => n978, S => n77, Y => n813);
   U1029 : INVX2 port map( A => keyTable_5_4_port, Y => n981);
   U1030 : INVX2 port map( A => KEY(44), Y => n980);
   U1031 : MUX2X1 port map( B => n981, A => n980, S => n80, Y => n812);
   U1032 : INVX2 port map( A => keyTable_5_3_port, Y => n983);
   U1033 : INVX2 port map( A => KEY(43), Y => n982);
   U1034 : MUX2X1 port map( B => n983, A => n982, S => n78, Y => n811);
   U1035 : INVX2 port map( A => keyTable_5_2_port, Y => n985);
   U1036 : INVX2 port map( A => KEY(42), Y => n984);
   U1037 : MUX2X1 port map( B => n985, A => n984, S => n143, Y => n810);
   U1038 : INVX2 port map( A => keyTable_5_1_port, Y => n987);
   U1039 : INVX2 port map( A => KEY(41), Y => n986);
   U1040 : MUX2X1 port map( B => n987, A => n986, S => n78, Y => n809);
   U1041 : INVX2 port map( A => keyTable_5_0_port, Y => n989);
   U1042 : INVX2 port map( A => KEY(40), Y => n988);
   U1043 : MUX2X1 port map( B => n989, A => n988, S => n77, Y => n808);
   U1044 : INVX2 port map( A => keyTable_6_7_port, Y => n991);
   U1045 : INVX2 port map( A => KEY(55), Y => n990);
   U1046 : MUX2X1 port map( B => n991, A => n990, S => n77, Y => n807);
   U1047 : INVX2 port map( A => keyTable_6_6_port, Y => n993);
   U1048 : INVX2 port map( A => KEY(54), Y => n992);
   U1049 : MUX2X1 port map( B => n993, A => n992, S => n78, Y => n806);
   U1050 : INVX2 port map( A => keyTable_6_5_port, Y => n995);
   U1051 : INVX2 port map( A => KEY(53), Y => n994);
   U1052 : MUX2X1 port map( B => n995, A => n994, S => n80, Y => n805);
   U1053 : INVX2 port map( A => keyTable_6_4_port, Y => n997);
   U1054 : INVX2 port map( A => KEY(52), Y => n996);
   U1055 : MUX2X1 port map( B => n997, A => n996, S => n82, Y => n804);
   U1056 : INVX2 port map( A => keyTable_6_3_port, Y => n999);
   U1057 : INVX2 port map( A => KEY(51), Y => n998);
   U1058 : MUX2X1 port map( B => n999, A => n998, S => n77, Y => n803);
   U1059 : INVX2 port map( A => keyTable_6_2_port, Y => n1001);
   U1060 : INVX2 port map( A => KEY(50), Y => n1000);
   U1061 : MUX2X1 port map( B => n1001, A => n1000, S => n82, Y => n802);
   U1062 : INVX2 port map( A => keyTable_6_1_port, Y => n1003);
   U1063 : INVX2 port map( A => KEY(49), Y => n1002);
   U1064 : MUX2X1 port map( B => n1003, A => n1002, S => n77, Y => n801);
   U1065 : INVX2 port map( A => keyTable_6_0_port, Y => n1005);
   U1066 : INVX2 port map( A => KEY(48), Y => n1004);
   U1067 : MUX2X1 port map( B => n1005, A => n1004, S => n82, Y => n800);
   U1068 : INVX2 port map( A => keyTable_7_7_port, Y => n1007);
   U1069 : INVX2 port map( A => KEY(63), Y => n1006);
   U1070 : MUX2X1 port map( B => n1007, A => n1006, S => n82, Y => n799);
   U1071 : INVX2 port map( A => keyTable_7_6_port, Y => n1009);
   U1072 : INVX2 port map( A => KEY(62), Y => n1008);
   U1073 : MUX2X1 port map( B => n1009, A => n1008, S => n80, Y => n798);
   U1074 : INVX2 port map( A => keyTable_7_5_port, Y => n1011);
   U1075 : INVX2 port map( A => KEY(61), Y => n1010);
   U1076 : MUX2X1 port map( B => n1011, A => n1010, S => n77, Y => n797);
   U1077 : INVX2 port map( A => keyTable_7_4_port, Y => n1013);
   U1078 : INVX2 port map( A => KEY(60), Y => n1012);
   U1079 : MUX2X1 port map( B => n1013, A => n1012, S => n143, Y => n796);
   U1080 : INVX2 port map( A => keyTable_7_3_port, Y => n1015);
   U1081 : INVX2 port map( A => KEY(59), Y => n1014);
   U1082 : MUX2X1 port map( B => n1015, A => n1014, S => n78, Y => n795);
   U1083 : INVX2 port map( A => keyTable_7_2_port, Y => n1017);
   U1084 : INVX2 port map( A => KEY(58), Y => n1016);
   U1085 : MUX2X1 port map( B => n1017, A => n1016, S => n77, Y => n794);
   U1086 : INVX2 port map( A => keyTable_7_1_port, Y => n1019);
   U1087 : INVX2 port map( A => KEY(57), Y => n1018);
   U1088 : MUX2X1 port map( B => n1019, A => n1018, S => n77, Y => n793);
   U1089 : INVX2 port map( A => keyTable_7_0_port, Y => n1021);
   U1090 : INVX2 port map( A => KEY(56), Y => n1020);
   U1091 : MUX2X1 port map( B => n1021, A => n1020, S => n78, Y => n792);
   U1092 : INVX2 port map( A => extratemp_0_port, Y => n1029);
   U1093 : INVX2 port map( A => DATA_IN(0), Y => n1028);
   U1094 : NAND2X1 port map( A => n28, B => n134, Y => n1023);
   U1095 : NAND2X1 port map( A => n1023, B => n1022, Y => n1024);
   U1096 : MUX2X1 port map( B => n1029, A => n1028, S => n1042, Y => n1127);
   U1097 : INVX2 port map( A => extratemp_1_port, Y => n1031);
   U1098 : INVX2 port map( A => DATA_IN(1), Y => n1030);
   U1099 : MUX2X1 port map( B => n1031, A => n1030, S => n1042, Y => n1128);
   U1100 : INVX2 port map( A => extratemp_2_port, Y => n1033);
   U1101 : INVX2 port map( A => DATA_IN(2), Y => n1032);
   U1102 : MUX2X1 port map( B => n1033, A => n1032, S => n1042, Y => n1129);
   U1103 : INVX2 port map( A => extratemp_3_port, Y => n1035);
   U1104 : INVX2 port map( A => DATA_IN(3), Y => n1034);
   U1105 : MUX2X1 port map( B => n1035, A => n1034, S => n1042, Y => n1130);
   U1106 : INVX2 port map( A => extratemp_4_port, Y => n1037);
   U1107 : INVX2 port map( A => DATA_IN(4), Y => n1036);
   U1108 : MUX2X1 port map( B => n1037, A => n1036, S => n1042, Y => n1131);
   U1109 : INVX2 port map( A => extratemp_5_port, Y => n1039);
   U1110 : INVX2 port map( A => DATA_IN(5), Y => n1038);
   U1111 : MUX2X1 port map( B => n1039, A => n1038, S => n1042, Y => n1132);
   U1112 : INVX2 port map( A => extratemp_6_port, Y => n1041);
   U1113 : INVX2 port map( A => DATA_IN(6), Y => n1040);
   U1114 : MUX2X1 port map( B => n1041, A => n1040, S => n1042, Y => n1133);
   U1115 : INVX2 port map( A => extratemp_7_port, Y => n1044);
   U1116 : INVX2 port map( A => DATA_IN(7), Y => n1043);
   U1117 : MUX2X1 port map( B => n1044, A => n1043, S => n1042, Y => n1134);
   U1118 : AOI21X1 port map( A => n12, B => n177, C => n1135, Y => n1053);
   U1119 : NAND2X1 port map( A => permuteComplete, B => n1046, Y => n1047);
   U1120 : NAND3X1 port map( A => n147, B => n70, C => n1047, Y => n1091);
   U1121 : INVX2 port map( A => n1091, Y => n1052);
   U1122 : OAI21X1 port map( A => n105, B => n107, C => n119, Y => n1049);
   U1123 : AOI22X1 port map( A => n1106, B => n1050, C => n134, D => n1049, Y 
                           => n1051);
   U1124 : NAND3X1 port map( A => n1053, B => n1052, C => n1051, Y => 
                           nextState_3_port);
   U1125 : OAI21X1 port map( A => n1055, B => n1057, C => n1054, Y => n1056);
   U1126 : NAND2X1 port map( A => n88, B => n1056, Y => n1059);
   U1127 : NAND2X1 port map( A => n1057, B => permuteComplete, Y => n1058);
   U1128 : NAND2X1 port map( A => n1059, B => n1058, Y => n899);
   U1129 : NAND3X1 port map( A => n1108, B => BYTE_READY, C => n1085, Y => 
                           n1063);
   U1130 : NAND2X1 port map( A => n128, B => n1084, Y => n1062);
   U1131 : NAND2X1 port map( A => n178, B => n1071, Y => n1061);
   U1132 : NAND3X1 port map( A => n1063, B => n1062, C => n1061, Y => n1064);
   U1133 : AOI21X1 port map( A => n1064, B => n1106, C => n645, Y => n1069);
   U1134 : NAND2X1 port map( A => n187, B => n30, Y => n1066);
   U1135 : NOR3X1 port map( A => n1067, B => n1066, C => n1135, Y => n1068);
   U1136 : NAND3X1 port map( A => n65, B => n1069, C => n1068, Y => 
                           nextState_0_port);
   U1137 : NAND2X1 port map( A => n105, B => n1071, Y => n1080);
   U1138 : INVX2 port map( A => n124, Y => n1072);
   U1139 : NAND2X1 port map( A => n1073, B => n1072, Y => n1079);
   U1140 : NAND2X1 port map( A => n1075, B => n133, Y => n1076);
   U1141 : AOI21X1 port map( A => n126, B => n1077, C => n1076, Y => n1078);
   U1142 : NAND3X1 port map( A => n1080, B => n1079, C => n1078, Y => 
                           nextState_4_port);
   U1143 : AND2X2 port map( A => n1082, B => n100, Y => n1083);
   U1144 : MUX2X1 port map( B => n177, A => n1083, S => n107, Y => n1095);
   U1145 : NAND2X1 port map( A => n155, B => n1084, Y => n1087);
   U1146 : NAND2X1 port map( A => n158, B => n1085, Y => n1086);
   U1147 : NAND2X1 port map( A => n1087, B => n1086, Y => n1088);
   U1148 : NAND2X1 port map( A => n1088, B => n1106, Y => n1094);
   U1149 : NAND2X1 port map( A => n1090, B => n93, Y => n1092);
   U1150 : NOR2X1 port map( A => n1092, B => n1091, Y => n1093);
   U1151 : NAND3X1 port map( A => n1095, B => n1094, C => n1093, Y => 
                           nextState_2_port);
   U1152 : INVX2 port map( A => N407, Y => n1097);
   U1153 : NAND2X1 port map( A => prefillCounter_0_port, B => n149, Y => n1096)
                           ;
   U1154 : OAI21X1 port map( A => n1098, B => n1097, C => n1096, Y => n915);
   U1155 : INVX2 port map( A => KEY_ERROR, Y => n1106);
   U1156 : INVX2 port map( A => BYTE_READY, Y => n1107);
   U1157 : INVX2 port map( A => n130, Y => n1108);
   U1158 : INVX2 port map( A => OPCODE(1), Y => n1109);
   U1159 : INVX2 port map( A => OPCODE(0), Y => n1110);
   n1137 <= '0';
   n1138 <= '0';

end SYN_bksa;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity transmitter_block_1 is

   port( PRGA_OUT : in std_logic_vector (7 downto 0);  clk, p_ready : in 
         std_logic;  prga_opcode : in std_logic_vector (1 downto 0);  rst : in 
         std_logic;  SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE : out std_logic);

end transmitter_block_1;

architecture SYN_struct of transmitter_block_1 is

   component tx_timer_1
      port( CLK, RST, SENDING : in std_logic;  SHIFT_ENABLE_R, SHIFT_ENABLE_E :
            out std_logic);
   end component;
   
   component tx_tcu_1
      port( clk, rst, p_ready, t_bitstuff : in std_logic;  PRGA_OUT : in 
            std_logic_vector (7 downto 0);  prga_opcode : in std_logic_vector 
            (1 downto 0);  t_crc : in std_logic_vector (15 downto 0);  sending,
            EOP, next_byte : out std_logic;  send_data : out std_logic_vector 
            (7 downto 0);  t_strobe : out std_logic);
   end component;
   
   component tx_shiftreg_1
      port( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe : in std_logic;  
            send_data : in std_logic_vector (7 downto 0);  d_encode : out 
            std_logic);
   end component;
   
   component tx_encode_1
      port( clk, rst, SHIFT_ENABLE_E, d_encode, EOP : in std_logic;  t_bitstuff
            , dp_tx_out, dm_tx_out : out std_logic);
   end component;
   
   component tx_CRC_CALC_1
      port( CLK, RST, EOP, T_STROBE : in std_logic;  PRGA_OPCODE : in 
            std_logic_vector (1 downto 0);  PRGA_OUT : in std_logic_vector (7 
            downto 0);  TX_CRC : out std_logic_vector (15 downto 0));
   end component;
   
   signal SENDING_port, t_strobe, EOP, TX_CRC_15_port, TX_CRC_14_port, 
      TX_CRC_13_port, TX_CRC_12_port, TX_CRC_11_port, TX_CRC_10_port, 
      TX_CRC_9_port, TX_CRC_8_port, TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port
      , TX_CRC_4_port, TX_CRC_3_port, TX_CRC_2_port, TX_CRC_1_port, 
      TX_CRC_0_port, SHIFT_ENABLE_E, d_encode, t_bitstuff, SHIFT_ENABLE_R, 
      send_data_7_port, send_data_6_port, send_data_5_port, send_data_4_port, 
      send_data_3_port, send_data_2_port, send_data_1_port, send_data_0_port : 
      std_logic;

begin
   SENDING <= SENDING_port;
   
   U_1 : tx_CRC_CALC_1 port map( CLK => clk, RST => rst, EOP => EOP, T_STROBE 
                           => t_strobe, PRGA_OPCODE(1) => prga_opcode(1), 
                           PRGA_OPCODE(0) => prga_opcode(0), PRGA_OUT(7) => 
                           PRGA_OUT(7), PRGA_OUT(6) => PRGA_OUT(6), PRGA_OUT(5)
                           => PRGA_OUT(5), PRGA_OUT(4) => PRGA_OUT(4), 
                           PRGA_OUT(3) => PRGA_OUT(3), PRGA_OUT(2) => 
                           PRGA_OUT(2), PRGA_OUT(1) => PRGA_OUT(1), PRGA_OUT(0)
                           => PRGA_OUT(0), TX_CRC(15) => TX_CRC_15_port, 
                           TX_CRC(14) => TX_CRC_14_port, TX_CRC(13) => 
                           TX_CRC_13_port, TX_CRC(12) => TX_CRC_12_port, 
                           TX_CRC(11) => TX_CRC_11_port, TX_CRC(10) => 
                           TX_CRC_10_port, TX_CRC(9) => TX_CRC_9_port, 
                           TX_CRC(8) => TX_CRC_8_port, TX_CRC(7) => 
                           TX_CRC_7_port, TX_CRC(6) => TX_CRC_6_port, TX_CRC(5)
                           => TX_CRC_5_port, TX_CRC(4) => TX_CRC_4_port, 
                           TX_CRC(3) => TX_CRC_3_port, TX_CRC(2) => 
                           TX_CRC_2_port, TX_CRC(1) => TX_CRC_1_port, TX_CRC(0)
                           => TX_CRC_0_port);
   U_0 : tx_encode_1 port map( clk => clk, rst => rst, SHIFT_ENABLE_E => 
                           SHIFT_ENABLE_E, d_encode => d_encode, EOP => EOP, 
                           t_bitstuff => t_bitstuff, dp_tx_out => dp_tx_out, 
                           dm_tx_out => dm_tx_out);
   U_2 : tx_shiftreg_1 port map( clk => clk, rst => rst, SHIFT_ENABLE_R => 
                           SHIFT_ENABLE_R, t_bitstuff => t_bitstuff, t_strobe 
                           => t_strobe, send_data(7) => send_data_7_port, 
                           send_data(6) => send_data_6_port, send_data(5) => 
                           send_data_5_port, send_data(4) => send_data_4_port, 
                           send_data(3) => send_data_3_port, send_data(2) => 
                           send_data_2_port, send_data(1) => send_data_1_port, 
                           send_data(0) => send_data_0_port, d_encode => 
                           d_encode);
   U_3 : tx_tcu_1 port map( clk => clk, rst => rst, p_ready => p_ready, 
                           t_bitstuff => t_bitstuff, PRGA_OUT(7) => PRGA_OUT(7)
                           , PRGA_OUT(6) => PRGA_OUT(6), PRGA_OUT(5) => 
                           PRGA_OUT(5), PRGA_OUT(4) => PRGA_OUT(4), PRGA_OUT(3)
                           => PRGA_OUT(3), PRGA_OUT(2) => PRGA_OUT(2), 
                           PRGA_OUT(1) => PRGA_OUT(1), PRGA_OUT(0) => 
                           PRGA_OUT(0), prga_opcode(1) => prga_opcode(1), 
                           prga_opcode(0) => prga_opcode(0), t_crc(15) => 
                           TX_CRC_15_port, t_crc(14) => TX_CRC_14_port, 
                           t_crc(13) => TX_CRC_13_port, t_crc(12) => 
                           TX_CRC_12_port, t_crc(11) => TX_CRC_11_port, 
                           t_crc(10) => TX_CRC_10_port, t_crc(9) => 
                           TX_CRC_9_port, t_crc(8) => TX_CRC_8_port, t_crc(7) 
                           => TX_CRC_7_port, t_crc(6) => TX_CRC_6_port, 
                           t_crc(5) => TX_CRC_5_port, t_crc(4) => TX_CRC_4_port
                           , t_crc(3) => TX_CRC_3_port, t_crc(2) => 
                           TX_CRC_2_port, t_crc(1) => TX_CRC_1_port, t_crc(0) 
                           => TX_CRC_0_port, sending => SENDING_port, EOP => 
                           EOP, next_byte => NEXT_BYTE, send_data(7) => 
                           send_data_7_port, send_data(6) => send_data_6_port, 
                           send_data(5) => send_data_5_port, send_data(4) => 
                           send_data_4_port, send_data(3) => send_data_3_port, 
                           send_data(2) => send_data_2_port, send_data(1) => 
                           send_data_1_port, send_data(0) => send_data_0_port, 
                           t_strobe => t_strobe);
   U_4 : tx_timer_1 port map( CLK => clk, RST => rst, SENDING => SENDING_port, 
                           SHIFT_ENABLE_R => SHIFT_ENABLE_R, SHIFT_ENABLE_E => 
                           SHIFT_ENABLE_E);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity receiver_block_rewire_1 is

   port( CLK, DM1_RX, DP1_RX, RST : in std_logic;  BS_ERROR, CRC_ERROR, 
         EOP_external : out std_logic;  OPCODE : out std_logic_vector (1 downto
         0);  RCV_DATA : out std_logic_vector (7 downto 0);  R_ERROR, W_ENABLE 
         : out std_logic);

end receiver_block_rewire_1;

architecture SYN_struct of receiver_block_rewire_1 is

   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component rx_timer_1
      port( CLK, RST, D_EDGE, RCVING : in std_logic;  SHIFT_ENABLE : out 
            std_logic);
   end component;
   
   component rx_shift_reg_1
      port( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF : in std_logic;  RCV_DATA 
            : out std_logic_vector (7 downto 0));
   end component;
   
   component rx_rcu_1
      port( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR : in 
            std_logic;  RX_CRC, RX_CHECK_CRC : in std_logic_vector (15 downto 
            0);  RCV_DATA : in std_logic_vector (7 downto 0);  RCVING, W_ENABLE
            , R_ERROR, CRC_ERROR : out std_logic;  OPCODE : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component rx_eopdetect_1
      port( DP1_RX, DM1_RX : in std_logic;  EOP : out std_logic);
   end component;
   
   component rx_edgedetect_1
      port( CLK, RST, DP1_RX : in std_logic;  D_EDGE : out std_logic);
   end component;
   
   component rx_decode_1
      port( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP : in std_logic;  D_ORIG, 
            BITSTUFF, BS_ERROR : out std_logic);
   end component;
   
   component rx_accumulator_1
      port( CLK, RST : in std_logic;  RCV_DATA : in std_logic_vector (7 downto 
            0);  W_ENABLE : in std_logic;  rx_CHECK_CRC : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component rx_CRC_CALC_1
      port( CLK, RST, W_ENABLE : in std_logic;  OPCODE : in std_logic_vector (1
            downto 0);  RCV_DATA : in std_logic_vector (7 downto 0);  RX_CRC : 
            out std_logic_vector (15 downto 0));
   end component;
   
   signal BS_ERROR_port, EOP_external_port, OPCODE_1_port, OPCODE_0_port, 
      RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, n8, RCV_DATA_1_port, RCV_DATA_0_port, W_ENABLE_port, 
      RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port, rx_CHECK_CRC_15_port, 
      rx_CHECK_CRC_14_port, rx_CHECK_CRC_13_port, rx_CHECK_CRC_12_port, 
      rx_CHECK_CRC_11_port, rx_CHECK_CRC_10_port, rx_CHECK_CRC_9_port, 
      rx_CHECK_CRC_8_port, rx_CHECK_CRC_7_port, rx_CHECK_CRC_6_port, 
      rx_CHECK_CRC_5_port, rx_CHECK_CRC_4_port, rx_CHECK_CRC_3_port, 
      rx_CHECK_CRC_2_port, rx_CHECK_CRC_1_port, rx_CHECK_CRC_0_port, 
      SHIFT_ENABLE, BITSTUFF, D_ORIG, D_EDGE, RCVING, n1, RCV_DATA_2_port, n3, 
      n4, n5, n6, n7 : std_logic;

begin
   BS_ERROR <= BS_ERROR_port;
   EOP_external <= EOP_external_port;
   OPCODE <= ( OPCODE_1_port, OPCODE_0_port );
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   W_ENABLE <= W_ENABLE_port;
   
   U_2 : rx_CRC_CALC_1 port map( CLK => CLK, RST => RST, W_ENABLE => n4, 
                           OPCODE(1) => n5, OPCODE(0) => n7, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           RX_CRC(15) => RX_CRC_15_port, RX_CRC(14) => 
                           RX_CRC_14_port, RX_CRC(13) => RX_CRC_13_port, 
                           RX_CRC(12) => RX_CRC_12_port, RX_CRC(11) => 
                           RX_CRC_11_port, RX_CRC(10) => RX_CRC_10_port, 
                           RX_CRC(9) => RX_CRC_9_port, RX_CRC(8) => 
                           RX_CRC_8_port, RX_CRC(7) => RX_CRC_7_port, RX_CRC(6)
                           => RX_CRC_6_port, RX_CRC(5) => RX_CRC_5_port, 
                           RX_CRC(4) => RX_CRC_4_port, RX_CRC(3) => 
                           RX_CRC_3_port, RX_CRC(2) => RX_CRC_2_port, RX_CRC(1)
                           => RX_CRC_1_port, RX_CRC(0) => RX_CRC_0_port);
   U_3 : rx_accumulator_1 port map( CLK => CLK, RST => RST, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           W_ENABLE => n4, rx_CHECK_CRC(15) => 
                           rx_CHECK_CRC_15_port, rx_CHECK_CRC(14) => 
                           rx_CHECK_CRC_14_port, rx_CHECK_CRC(13) => 
                           rx_CHECK_CRC_13_port, rx_CHECK_CRC(12) => 
                           rx_CHECK_CRC_12_port, rx_CHECK_CRC(11) => 
                           rx_CHECK_CRC_11_port, rx_CHECK_CRC(10) => 
                           rx_CHECK_CRC_10_port, rx_CHECK_CRC(9) => 
                           rx_CHECK_CRC_9_port, rx_CHECK_CRC(8) => 
                           rx_CHECK_CRC_8_port, rx_CHECK_CRC(7) => 
                           rx_CHECK_CRC_7_port, rx_CHECK_CRC(6) => 
                           rx_CHECK_CRC_6_port, rx_CHECK_CRC(5) => 
                           rx_CHECK_CRC_5_port, rx_CHECK_CRC(4) => 
                           rx_CHECK_CRC_4_port, rx_CHECK_CRC(3) => 
                           rx_CHECK_CRC_3_port, rx_CHECK_CRC(2) => 
                           rx_CHECK_CRC_2_port, rx_CHECK_CRC(1) => 
                           rx_CHECK_CRC_1_port, rx_CHECK_CRC(0) => 
                           rx_CHECK_CRC_0_port);
   U_1 : rx_decode_1 port map( CLK => CLK, RST => RST, DP1_RX => DP1_RX, 
                           SHIFT_ENABLE => n6, EOP => EOP_external_port, D_ORIG
                           => D_ORIG, BITSTUFF => BITSTUFF, BS_ERROR => 
                           BS_ERROR_port);
   U_0 : rx_edgedetect_1 port map( CLK => CLK, RST => RST, DP1_RX => DP1_RX, 
                           D_EDGE => D_EDGE);
   U_4 : rx_eopdetect_1 port map( DP1_RX => DP1_RX, DM1_RX => DM1_RX, EOP => 
                           EOP_external_port);
   U_5 : rx_rcu_1 port map( CLK => CLK, RST => RST, D_EDGE => n1, EOP => 
                           EOP_external_port, SHIFT_ENABLE => SHIFT_ENABLE, 
                           BITSTUFF => BITSTUFF, BS_ERROR => BS_ERROR_port, 
                           RX_CRC(15) => RX_CRC_15_port, RX_CRC(14) => 
                           RX_CRC_14_port, RX_CRC(13) => RX_CRC_13_port, 
                           RX_CRC(12) => RX_CRC_12_port, RX_CRC(11) => 
                           RX_CRC_11_port, RX_CRC(10) => RX_CRC_10_port, 
                           RX_CRC(9) => RX_CRC_9_port, RX_CRC(8) => 
                           RX_CRC_8_port, RX_CRC(7) => RX_CRC_7_port, RX_CRC(6)
                           => RX_CRC_6_port, RX_CRC(5) => RX_CRC_5_port, 
                           RX_CRC(4) => RX_CRC_4_port, RX_CRC(3) => 
                           RX_CRC_3_port, RX_CRC(2) => RX_CRC_2_port, RX_CRC(1)
                           => RX_CRC_1_port, RX_CRC(0) => RX_CRC_0_port, 
                           RX_CHECK_CRC(15) => rx_CHECK_CRC_15_port, 
                           RX_CHECK_CRC(14) => rx_CHECK_CRC_14_port, 
                           RX_CHECK_CRC(13) => rx_CHECK_CRC_13_port, 
                           RX_CHECK_CRC(12) => rx_CHECK_CRC_12_port, 
                           RX_CHECK_CRC(11) => rx_CHECK_CRC_11_port, 
                           RX_CHECK_CRC(10) => rx_CHECK_CRC_10_port, 
                           RX_CHECK_CRC(9) => rx_CHECK_CRC_9_port, 
                           RX_CHECK_CRC(8) => rx_CHECK_CRC_8_port, 
                           RX_CHECK_CRC(7) => rx_CHECK_CRC_7_port, 
                           RX_CHECK_CRC(6) => rx_CHECK_CRC_6_port, 
                           RX_CHECK_CRC(5) => rx_CHECK_CRC_5_port, 
                           RX_CHECK_CRC(4) => rx_CHECK_CRC_4_port, 
                           RX_CHECK_CRC(3) => rx_CHECK_CRC_3_port, 
                           RX_CHECK_CRC(2) => rx_CHECK_CRC_2_port, 
                           RX_CHECK_CRC(1) => rx_CHECK_CRC_1_port, 
                           RX_CHECK_CRC(0) => rx_CHECK_CRC_0_port, RCV_DATA(7) 
                           => RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => n8, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, RCVING => RCVING, 
                           W_ENABLE => W_ENABLE_port, R_ERROR => R_ERROR, 
                           CRC_ERROR => CRC_ERROR, OPCODE(1) => OPCODE_1_port, 
                           OPCODE(0) => OPCODE_0_port);
   U_6 : rx_shift_reg_1 port map( CLK => CLK, RST => RST, SHIFT_ENABLE => 
                           SHIFT_ENABLE, D_ORIG => D_ORIG, BITSTUFF => BITSTUFF
                           , RCV_DATA(7) => RCV_DATA_7_port, RCV_DATA(6) => 
                           RCV_DATA_6_port, RCV_DATA(5) => RCV_DATA_5_port, 
                           RCV_DATA(4) => RCV_DATA_4_port, RCV_DATA(3) => 
                           RCV_DATA_3_port, RCV_DATA(2) => n8, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port);
   U_7 : rx_timer_1 port map( CLK => CLK, RST => RST, D_EDGE => D_EDGE, RCVING 
                           => RCVING, SHIFT_ENABLE => SHIFT_ENABLE);
   U1 : BUFX2 port map( A => D_EDGE, Y => n1);
   U2 : BUFX2 port map( A => n8, Y => RCV_DATA_2_port);
   U3 : BUFX4 port map( A => SHIFT_ENABLE, Y => n6);
   U4 : INVX1 port map( A => W_ENABLE_port, Y => n3);
   U5 : INVX2 port map( A => n3, Y => n4);
   U6 : BUFX2 port map( A => OPCODE_1_port, Y => n5);
   U7 : BUFX2 port map( A => OPCODE_0_port, Y => n7);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity memoryblock_1 is

   port( CLK, NEXT_BYTE : in std_logic;  RCV_DATA : in std_logic_vector (7 
         downto 0);  RCV_OPCODE : in std_logic_vector (1 downto 0);  RST, 
         W_ENABLE, EOP : in std_logic;  EMPTY, FULL, B_READY : out std_logic;  
         PRGA_IN : out std_logic_vector (7 downto 0);  PRGA_OPCODE : out 
         std_logic_vector (1 downto 0));

end memoryblock_1;

architecture SYN_struct of memoryblock_1 is

   component RFIFO_1
      port( CLK, RST, W_ENABLE, R_ENABLE : in std_logic;  RCV_DATA : in 
            std_logic_vector (7 downto 0);  RCV_OPCODE : in std_logic_vector (1
            downto 0);  DATA : out std_logic_vector (7 downto 0);  OUT_OPCODE :
            out std_logic_vector (1 downto 0);  BYTE_COUNT : out 
            std_logic_vector (4 downto 0);  EMPTY, FULL : out std_logic);
   end component;
   
   component RBUFFER_1
      port( CLK, RST, NEXT_BYTE : in std_logic;  DATA : in std_logic_vector (7 
            downto 0);  OPCODE : in std_logic_vector (1 downto 0);  BYTE_COUNT 
            : in std_logic_vector (4 downto 0);  EOP : in std_logic;  B_READY, 
            R_ENABLE : out std_logic;  PRGA_IN : out std_logic_vector (7 downto
            0);  PRGA_OPCODE : out std_logic_vector (1 downto 0));
   end component;
   
   signal BYTE_COUNT_4_port, BYTE_COUNT_3_port, BYTE_COUNT_2_port, 
      BYTE_COUNT_1_port, BYTE_COUNT_0_port, DATA_7_port, DATA_6_port, 
      DATA_5_port, DATA_4_port, DATA_3_port, DATA_2_port, DATA_1_port, 
      DATA_0_port, OUT_OPCODE_1_port, OUT_OPCODE_0_port, R_ENABLE : std_logic;

begin
   
   U_0 : RBUFFER_1 port map( CLK => CLK, RST => RST, NEXT_BYTE => NEXT_BYTE, 
                           DATA(7) => DATA_7_port, DATA(6) => DATA_6_port, 
                           DATA(5) => DATA_5_port, DATA(4) => DATA_4_port, 
                           DATA(3) => DATA_3_port, DATA(2) => DATA_2_port, 
                           DATA(1) => DATA_1_port, DATA(0) => DATA_0_port, 
                           OPCODE(1) => OUT_OPCODE_1_port, OPCODE(0) => 
                           OUT_OPCODE_0_port, BYTE_COUNT(4) => 
                           BYTE_COUNT_4_port, BYTE_COUNT(3) => 
                           BYTE_COUNT_3_port, BYTE_COUNT(2) => 
                           BYTE_COUNT_2_port, BYTE_COUNT(1) => 
                           BYTE_COUNT_1_port, BYTE_COUNT(0) => 
                           BYTE_COUNT_0_port, EOP => EOP, B_READY => B_READY, 
                           R_ENABLE => R_ENABLE, PRGA_IN(7) => PRGA_IN(7), 
                           PRGA_IN(6) => PRGA_IN(6), PRGA_IN(5) => PRGA_IN(5), 
                           PRGA_IN(4) => PRGA_IN(4), PRGA_IN(3) => PRGA_IN(3), 
                           PRGA_IN(2) => PRGA_IN(2), PRGA_IN(1) => PRGA_IN(1), 
                           PRGA_IN(0) => PRGA_IN(0), PRGA_OPCODE(1) => 
                           PRGA_OPCODE(1), PRGA_OPCODE(0) => PRGA_OPCODE(0));
   U_1 : RFIFO_1 port map( CLK => CLK, RST => RST, W_ENABLE => W_ENABLE, 
                           R_ENABLE => R_ENABLE, RCV_DATA(7) => RCV_DATA(7), 
                           RCV_DATA(6) => RCV_DATA(6), RCV_DATA(5) => 
                           RCV_DATA(5), RCV_DATA(4) => RCV_DATA(4), RCV_DATA(3)
                           => RCV_DATA(3), RCV_DATA(2) => RCV_DATA(2), 
                           RCV_DATA(1) => RCV_DATA(1), RCV_DATA(0) => 
                           RCV_DATA(0), RCV_OPCODE(1) => RCV_OPCODE(1), 
                           RCV_OPCODE(0) => RCV_OPCODE(0), DATA(7) => 
                           DATA_7_port, DATA(6) => DATA_6_port, DATA(5) => 
                           DATA_5_port, DATA(4) => DATA_4_port, DATA(3) => 
                           DATA_3_port, DATA(2) => DATA_2_port, DATA(1) => 
                           DATA_1_port, DATA(0) => DATA_0_port, OUT_OPCODE(1) 
                           => OUT_OPCODE_1_port, OUT_OPCODE(0) => 
                           OUT_OPCODE_0_port, BYTE_COUNT(4) => 
                           BYTE_COUNT_4_port, BYTE_COUNT(3) => 
                           BYTE_COUNT_3_port, BYTE_COUNT(2) => 
                           BYTE_COUNT_2_port, BYTE_COUNT(1) => 
                           BYTE_COUNT_1_port, BYTE_COUNT(0) => 
                           BYTE_COUNT_0_port, EMPTY => EMPTY, FULL => FULL);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity EDBlock_1 is

   port( BYTE : in std_logic_vector (7 downto 0);  BYTE_READY, CLK : in 
         std_logic;  OPCODE : in std_logic_vector (1 downto 0);  RST, SERIAL_IN
         : in std_logic;  DATA_IN : in std_logic_vector (7 downto 0);  
         KEY_ERROR, PARITY_ERROR, PDATA_READY : out std_logic;  PROCESSED_DATA 
         : out std_logic_vector (7 downto 0);  PROG_ERROR, RBUF_FULL, W_ENABLE,
         R_ENABLE : out std_logic;  DATA, ADDR : out std_logic_vector (7 downto
         0));

end EDBlock_1;

architecture SYN_struct of EDBlock_1 is

   component uart_rcv_block_1
      port( CLK, RST, SERIAL_IN : in std_logic;  KEY_ERROR, PROG_ERROR : out 
            std_logic;  PLAINKEY : out std_logic_vector (63 downto 0);  
            RBUF_FULL, PARITY_ERROR : out std_logic);
   end component;
   
   component KSA_1
      port( KEY : in std_logic_vector (63 downto 0);  CLK, RST, KEY_ERROR, 
            BYTE_READY : in std_logic;  BYTE : in std_logic_vector (7 downto 0)
            ;  OPCODE : in std_logic_vector (1 downto 0);  DATA_IN : in 
            std_logic_vector (7 downto 0);  PROCESSED_DATA : out 
            std_logic_vector (7 downto 0);  PDATA_READY, W_ENABLE, R_ENABLE : 
            out std_logic;  ADDR, DATA : out std_logic_vector (7 downto 0));
   end component;
   
   signal KEY_ERROR_port, PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port,
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port : std_logic;

begin
   KEY_ERROR <= KEY_ERROR_port;
   
   U_0 : KSA_1 port map( KEY(63) => PLAINKEY_63_port, KEY(62) => 
                           PLAINKEY_62_port, KEY(61) => PLAINKEY_61_port, 
                           KEY(60) => PLAINKEY_60_port, KEY(59) => 
                           PLAINKEY_59_port, KEY(58) => PLAINKEY_58_port, 
                           KEY(57) => PLAINKEY_57_port, KEY(56) => 
                           PLAINKEY_56_port, KEY(55) => PLAINKEY_55_port, 
                           KEY(54) => PLAINKEY_54_port, KEY(53) => 
                           PLAINKEY_53_port, KEY(52) => PLAINKEY_52_port, 
                           KEY(51) => PLAINKEY_51_port, KEY(50) => 
                           PLAINKEY_50_port, KEY(49) => PLAINKEY_49_port, 
                           KEY(48) => PLAINKEY_48_port, KEY(47) => 
                           PLAINKEY_47_port, KEY(46) => PLAINKEY_46_port, 
                           KEY(45) => PLAINKEY_45_port, KEY(44) => 
                           PLAINKEY_44_port, KEY(43) => PLAINKEY_43_port, 
                           KEY(42) => PLAINKEY_42_port, KEY(41) => 
                           PLAINKEY_41_port, KEY(40) => PLAINKEY_40_port, 
                           KEY(39) => PLAINKEY_39_port, KEY(38) => 
                           PLAINKEY_38_port, KEY(37) => PLAINKEY_37_port, 
                           KEY(36) => PLAINKEY_36_port, KEY(35) => 
                           PLAINKEY_35_port, KEY(34) => PLAINKEY_34_port, 
                           KEY(33) => PLAINKEY_33_port, KEY(32) => 
                           PLAINKEY_32_port, KEY(31) => PLAINKEY_31_port, 
                           KEY(30) => PLAINKEY_30_port, KEY(29) => 
                           PLAINKEY_29_port, KEY(28) => PLAINKEY_28_port, 
                           KEY(27) => PLAINKEY_27_port, KEY(26) => 
                           PLAINKEY_26_port, KEY(25) => PLAINKEY_25_port, 
                           KEY(24) => PLAINKEY_24_port, KEY(23) => 
                           PLAINKEY_23_port, KEY(22) => PLAINKEY_22_port, 
                           KEY(21) => PLAINKEY_21_port, KEY(20) => 
                           PLAINKEY_20_port, KEY(19) => PLAINKEY_19_port, 
                           KEY(18) => PLAINKEY_18_port, KEY(17) => 
                           PLAINKEY_17_port, KEY(16) => PLAINKEY_16_port, 
                           KEY(15) => PLAINKEY_15_port, KEY(14) => 
                           PLAINKEY_14_port, KEY(13) => PLAINKEY_13_port, 
                           KEY(12) => PLAINKEY_12_port, KEY(11) => 
                           PLAINKEY_11_port, KEY(10) => PLAINKEY_10_port, 
                           KEY(9) => PLAINKEY_9_port, KEY(8) => PLAINKEY_8_port
                           , KEY(7) => PLAINKEY_7_port, KEY(6) => 
                           PLAINKEY_6_port, KEY(5) => PLAINKEY_5_port, KEY(4) 
                           => PLAINKEY_4_port, KEY(3) => PLAINKEY_3_port, 
                           KEY(2) => PLAINKEY_2_port, KEY(1) => PLAINKEY_1_port
                           , KEY(0) => PLAINKEY_0_port, CLK => CLK, RST => RST,
                           KEY_ERROR => KEY_ERROR_port, BYTE_READY => 
                           BYTE_READY, BYTE(7) => BYTE(7), BYTE(6) => BYTE(6), 
                           BYTE(5) => BYTE(5), BYTE(4) => BYTE(4), BYTE(3) => 
                           BYTE(3), BYTE(2) => BYTE(2), BYTE(1) => BYTE(1), 
                           BYTE(0) => BYTE(0), OPCODE(1) => OPCODE(1), 
                           OPCODE(0) => OPCODE(0), DATA_IN(7) => DATA_IN(7), 
                           DATA_IN(6) => DATA_IN(6), DATA_IN(5) => DATA_IN(5), 
                           DATA_IN(4) => DATA_IN(4), DATA_IN(3) => DATA_IN(3), 
                           DATA_IN(2) => DATA_IN(2), DATA_IN(1) => DATA_IN(1), 
                           DATA_IN(0) => DATA_IN(0), PROCESSED_DATA(7) => 
                           PROCESSED_DATA(7), PROCESSED_DATA(6) => 
                           PROCESSED_DATA(6), PROCESSED_DATA(5) => 
                           PROCESSED_DATA(5), PROCESSED_DATA(4) => 
                           PROCESSED_DATA(4), PROCESSED_DATA(3) => 
                           PROCESSED_DATA(3), PROCESSED_DATA(2) => 
                           PROCESSED_DATA(2), PROCESSED_DATA(1) => 
                           PROCESSED_DATA(1), PROCESSED_DATA(0) => 
                           PROCESSED_DATA(0), PDATA_READY => PDATA_READY, 
                           W_ENABLE => W_ENABLE, R_ENABLE => R_ENABLE, ADDR(7) 
                           => ADDR(7), ADDR(6) => ADDR(6), ADDR(5) => ADDR(5), 
                           ADDR(4) => ADDR(4), ADDR(3) => ADDR(3), ADDR(2) => 
                           ADDR(2), ADDR(1) => ADDR(1), ADDR(0) => ADDR(0), 
                           DATA(7) => DATA(7), DATA(6) => DATA(6), DATA(5) => 
                           DATA(5), DATA(4) => DATA(4), DATA(3) => DATA(3), 
                           DATA(2) => DATA(2), DATA(1) => DATA(1), DATA(0) => 
                           DATA(0));
   U_1 : uart_rcv_block_1 port map( CLK => CLK, RST => RST, SERIAL_IN => 
                           SERIAL_IN, KEY_ERROR => KEY_ERROR_port, PROG_ERROR 
                           => PROG_ERROR, PLAINKEY(63) => PLAINKEY_63_port, 
                           PLAINKEY(62) => PLAINKEY_62_port, PLAINKEY(61) => 
                           PLAINKEY_61_port, PLAINKEY(60) => PLAINKEY_60_port, 
                           PLAINKEY(59) => PLAINKEY_59_port, PLAINKEY(58) => 
                           PLAINKEY_58_port, PLAINKEY(57) => PLAINKEY_57_port, 
                           PLAINKEY(56) => PLAINKEY_56_port, PLAINKEY(55) => 
                           PLAINKEY_55_port, PLAINKEY(54) => PLAINKEY_54_port, 
                           PLAINKEY(53) => PLAINKEY_53_port, PLAINKEY(52) => 
                           PLAINKEY_52_port, PLAINKEY(51) => PLAINKEY_51_port, 
                           PLAINKEY(50) => PLAINKEY_50_port, PLAINKEY(49) => 
                           PLAINKEY_49_port, PLAINKEY(48) => PLAINKEY_48_port, 
                           PLAINKEY(47) => PLAINKEY_47_port, PLAINKEY(46) => 
                           PLAINKEY_46_port, PLAINKEY(45) => PLAINKEY_45_port, 
                           PLAINKEY(44) => PLAINKEY_44_port, PLAINKEY(43) => 
                           PLAINKEY_43_port, PLAINKEY(42) => PLAINKEY_42_port, 
                           PLAINKEY(41) => PLAINKEY_41_port, PLAINKEY(40) => 
                           PLAINKEY_40_port, PLAINKEY(39) => PLAINKEY_39_port, 
                           PLAINKEY(38) => PLAINKEY_38_port, PLAINKEY(37) => 
                           PLAINKEY_37_port, PLAINKEY(36) => PLAINKEY_36_port, 
                           PLAINKEY(35) => PLAINKEY_35_port, PLAINKEY(34) => 
                           PLAINKEY_34_port, PLAINKEY(33) => PLAINKEY_33_port, 
                           PLAINKEY(32) => PLAINKEY_32_port, PLAINKEY(31) => 
                           PLAINKEY_31_port, PLAINKEY(30) => PLAINKEY_30_port, 
                           PLAINKEY(29) => PLAINKEY_29_port, PLAINKEY(28) => 
                           PLAINKEY_28_port, PLAINKEY(27) => PLAINKEY_27_port, 
                           PLAINKEY(26) => PLAINKEY_26_port, PLAINKEY(25) => 
                           PLAINKEY_25_port, PLAINKEY(24) => PLAINKEY_24_port, 
                           PLAINKEY(23) => PLAINKEY_23_port, PLAINKEY(22) => 
                           PLAINKEY_22_port, PLAINKEY(21) => PLAINKEY_21_port, 
                           PLAINKEY(20) => PLAINKEY_20_port, PLAINKEY(19) => 
                           PLAINKEY_19_port, PLAINKEY(18) => PLAINKEY_18_port, 
                           PLAINKEY(17) => PLAINKEY_17_port, PLAINKEY(16) => 
                           PLAINKEY_16_port, PLAINKEY(15) => PLAINKEY_15_port, 
                           PLAINKEY(14) => PLAINKEY_14_port, PLAINKEY(13) => 
                           PLAINKEY_13_port, PLAINKEY(12) => PLAINKEY_12_port, 
                           PLAINKEY(11) => PLAINKEY_11_port, PLAINKEY(10) => 
                           PLAINKEY_10_port, PLAINKEY(9) => PLAINKEY_9_port, 
                           PLAINKEY(8) => PLAINKEY_8_port, PLAINKEY(7) => 
                           PLAINKEY_7_port, PLAINKEY(6) => PLAINKEY_6_port, 
                           PLAINKEY(5) => PLAINKEY_5_port, PLAINKEY(4) => 
                           PLAINKEY_4_port, PLAINKEY(3) => PLAINKEY_3_port, 
                           PLAINKEY(2) => PLAINKEY_2_port, PLAINKEY(1) => 
                           PLAINKEY_1_port, PLAINKEY(0) => PLAINKEY_0_port, 
                           RBUF_FULL => RBUF_FULL, PARITY_ERROR => PARITY_ERROR
                           );

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RMEDT_REWIRE_1 is

   port( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN : in std_logic;  DATA_IN : in 
         std_logic_vector (7 downto 0);  BS_ERROR, CRC_ERROR, EMPTY, FULL, 
         KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, R_ERROR, SENDING, 
         dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE : out std_logic;  DATA, 
         ADDR : out std_logic_vector (7 downto 0));

end RMEDT_REWIRE_1;

architecture SYN_struct of RMEDT_REWIRE_1 is

   component transmitter_block_1
      port( PRGA_OUT : in std_logic_vector (7 downto 0);  clk, p_ready : in 
            std_logic;  prga_opcode : in std_logic_vector (1 downto 0);  rst : 
            in std_logic;  SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE : out 
            std_logic);
   end component;
   
   component receiver_block_rewire_1
      port( CLK, DM1_RX, DP1_RX, RST : in std_logic;  BS_ERROR, CRC_ERROR, 
            EOP_external : out std_logic;  OPCODE : out std_logic_vector (1 
            downto 0);  RCV_DATA : out std_logic_vector (7 downto 0);  R_ERROR,
            W_ENABLE : out std_logic);
   end component;
   
   component memoryblock_1
      port( CLK, NEXT_BYTE : in std_logic;  RCV_DATA : in std_logic_vector (7 
            downto 0);  RCV_OPCODE : in std_logic_vector (1 downto 0);  RST, 
            W_ENABLE, EOP : in std_logic;  EMPTY, FULL, B_READY : out std_logic
            ;  PRGA_IN : out std_logic_vector (7 downto 0);  PRGA_OPCODE : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component EDBlock_1
      port( BYTE : in std_logic_vector (7 downto 0);  BYTE_READY, CLK : in 
            std_logic;  OPCODE : in std_logic_vector (1 downto 0);  RST, 
            SERIAL_IN : in std_logic;  DATA_IN : in std_logic_vector (7 downto 
            0);  KEY_ERROR, PARITY_ERROR, PDATA_READY : out std_logic;  
            PROCESSED_DATA : out std_logic_vector (7 downto 0);  PROG_ERROR, 
            RBUF_FULL, W_ENABLE, R_ENABLE : out std_logic;  DATA, ADDR : out 
            std_logic_vector (7 downto 0));
   end component;
   
   signal PRGA_IN_7_port, PRGA_IN_6_port, PRGA_IN_5_port, PRGA_IN_4_port, 
      PRGA_IN_3_port, PRGA_IN_2_port, PRGA_IN_1_port, PRGA_IN_0_port, B_READY, 
      PRGA_OPCODE_1_port, PRGA_OPCODE_0_port, PDATA_READY, 
      PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, PROCESSED_DATA_5_port, 
      PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, PROCESSED_DATA_2_port, 
      PROCESSED_DATA_1_port, PROCESSED_DATA_0_port, EOP_external, NEXT_BYTE, 
      RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      OPCODE_1_port, OPCODE_0_port, W_ENABLE : std_logic;

begin
   
   U_0 : EDBlock_1 port map( BYTE(7) => PRGA_IN_7_port, BYTE(6) => 
                           PRGA_IN_6_port, BYTE(5) => PRGA_IN_5_port, BYTE(4) 
                           => PRGA_IN_4_port, BYTE(3) => PRGA_IN_3_port, 
                           BYTE(2) => PRGA_IN_2_port, BYTE(1) => PRGA_IN_1_port
                           , BYTE(0) => PRGA_IN_0_port, BYTE_READY => B_READY, 
                           CLK => CLK, OPCODE(1) => PRGA_OPCODE_1_port, 
                           OPCODE(0) => PRGA_OPCODE_0_port, RST => RST, 
                           SERIAL_IN => SERIAL_IN, DATA_IN(7) => DATA_IN(7), 
                           DATA_IN(6) => DATA_IN(6), DATA_IN(5) => DATA_IN(5), 
                           DATA_IN(4) => DATA_IN(4), DATA_IN(3) => DATA_IN(3), 
                           DATA_IN(2) => DATA_IN(2), DATA_IN(1) => DATA_IN(1), 
                           DATA_IN(0) => DATA_IN(0), KEY_ERROR => KEY_ERROR, 
                           PARITY_ERROR => PARITY_ERROR, PDATA_READY => 
                           PDATA_READY, PROCESSED_DATA(7) => 
                           PROCESSED_DATA_7_port, PROCESSED_DATA(6) => 
                           PROCESSED_DATA_6_port, PROCESSED_DATA(5) => 
                           PROCESSED_DATA_5_port, PROCESSED_DATA(4) => 
                           PROCESSED_DATA_4_port, PROCESSED_DATA(3) => 
                           PROCESSED_DATA_3_port, PROCESSED_DATA(2) => 
                           PROCESSED_DATA_2_port, PROCESSED_DATA(1) => 
                           PROCESSED_DATA_1_port, PROCESSED_DATA(0) => 
                           PROCESSED_DATA_0_port, PROG_ERROR => PROG_ERROR, 
                           RBUF_FULL => RBUF_FULL, W_ENABLE => W_ENABLE_R, 
                           R_ENABLE => R_ENABLE, DATA(7) => DATA(7), DATA(6) =>
                           DATA(6), DATA(5) => DATA(5), DATA(4) => DATA(4), 
                           DATA(3) => DATA(3), DATA(2) => DATA(2), DATA(1) => 
                           DATA(1), DATA(0) => DATA(0), ADDR(7) => ADDR(7), 
                           ADDR(6) => ADDR(6), ADDR(5) => ADDR(5), ADDR(4) => 
                           ADDR(4), ADDR(3) => ADDR(3), ADDR(2) => ADDR(2), 
                           ADDR(1) => ADDR(1), ADDR(0) => ADDR(0));
   U_1 : memoryblock_1 port map( CLK => CLK, NEXT_BYTE => NEXT_BYTE, 
                           RCV_DATA(7) => RCV_DATA_7_port, RCV_DATA(6) => 
                           RCV_DATA_6_port, RCV_DATA(5) => RCV_DATA_5_port, 
                           RCV_DATA(4) => RCV_DATA_4_port, RCV_DATA(3) => 
                           RCV_DATA_3_port, RCV_DATA(2) => RCV_DATA_2_port, 
                           RCV_DATA(1) => RCV_DATA_1_port, RCV_DATA(0) => 
                           RCV_DATA_0_port, RCV_OPCODE(1) => OPCODE_1_port, 
                           RCV_OPCODE(0) => OPCODE_0_port, RST => RST, W_ENABLE
                           => W_ENABLE, EOP => EOP_external, EMPTY => EMPTY, 
                           FULL => FULL, B_READY => B_READY, PRGA_IN(7) => 
                           PRGA_IN_7_port, PRGA_IN(6) => PRGA_IN_6_port, 
                           PRGA_IN(5) => PRGA_IN_5_port, PRGA_IN(4) => 
                           PRGA_IN_4_port, PRGA_IN(3) => PRGA_IN_3_port, 
                           PRGA_IN(2) => PRGA_IN_2_port, PRGA_IN(1) => 
                           PRGA_IN_1_port, PRGA_IN(0) => PRGA_IN_0_port, 
                           PRGA_OPCODE(1) => PRGA_OPCODE_1_port, PRGA_OPCODE(0)
                           => PRGA_OPCODE_0_port);
   U_2 : receiver_block_rewire_1 port map( CLK => CLK, DM1_RX => DM1_RX, DP1_RX
                           => DP1_RX, RST => RST, BS_ERROR => BS_ERROR, 
                           CRC_ERROR => CRC_ERROR, EOP_external => EOP_external
                           , OPCODE(1) => OPCODE_1_port, OPCODE(0) => 
                           OPCODE_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, R_ERROR => R_ERROR, 
                           W_ENABLE => W_ENABLE);
   U_3 : transmitter_block_1 port map( PRGA_OUT(7) => PROCESSED_DATA_7_port, 
                           PRGA_OUT(6) => PROCESSED_DATA_6_port, PRGA_OUT(5) =>
                           PROCESSED_DATA_5_port, PRGA_OUT(4) => 
                           PROCESSED_DATA_4_port, PRGA_OUT(3) => 
                           PROCESSED_DATA_3_port, PRGA_OUT(2) => 
                           PROCESSED_DATA_2_port, PRGA_OUT(1) => 
                           PROCESSED_DATA_1_port, PRGA_OUT(0) => 
                           PROCESSED_DATA_0_port, clk => CLK, p_ready => 
                           PDATA_READY, prga_opcode(1) => PRGA_OPCODE_1_port, 
                           prga_opcode(0) => PRGA_OPCODE_0_port, rst => RST, 
                           SENDING => SENDING, dm_tx_out => dm_tx_out, 
                           dp_tx_out => dp_tx_out, NEXT_BYTE => NEXT_BYTE);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rmedt_square is

   port( CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN : in std_logic;  DATA_IN_H
         , DATA_IN_S : in std_logic_vector (7 downto 0);  BSE_H, BSE_S, CRCE_H,
         CRCE_S, DMTH, DMTS, DPTH, DPTS, EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H
         , RE_S, c_key_error, c_parity_error, c_prog_error, host_is_sending, 
         slave_is_sending, W_ENABLE_H, W_ENABLE_S, R_ENABLE_H, R_ENABLE_S : out
         std_logic;  DATA_H, DATA_S, ADDR_H, ADDR_S : out std_logic_vector (7 
         downto 0));

end rmedt_square;

architecture SYN_struct of rmedt_square is

   component RMEDT_REWIRE_0
      port( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN : in std_logic;  DATA_IN : in 
            std_logic_vector (7 downto 0);  BS_ERROR, CRC_ERROR, EMPTY, FULL, 
            KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, R_ERROR, SENDING, 
            dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE : out std_logic;  DATA, 
            ADDR : out std_logic_vector (7 downto 0));
   end component;
   
   component RMEDT_REWIRE_1
      port( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN : in std_logic;  DATA_IN : in 
            std_logic_vector (7 downto 0);  BS_ERROR, CRC_ERROR, EMPTY, FULL, 
            KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, R_ERROR, SENDING, 
            dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE : out std_logic;  DATA, 
            ADDR : out std_logic_vector (7 downto 0));
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal KEY_ERROR, KEY_ERROR1, PARITY_ERROR, PARITY_ERROR1, PROG_ERROR, 
      PROG_ERROR1, n_1036, n_1037 : std_logic;

begin
   
   U1 : OR2X2 port map( A => PROG_ERROR, B => PROG_ERROR1, Y => c_prog_error);
   U2 : OR2X2 port map( A => PARITY_ERROR, B => PARITY_ERROR1, Y => 
                           c_parity_error);
   U3 : OR2X2 port map( A => KEY_ERROR, B => KEY_ERROR1, Y => c_key_error);
   U_0 : RMEDT_REWIRE_1 port map( CLK => CLK, DM1_RX => DMRH, DP1_RX => DPRH, 
                           RST => RST, SERIAL_IN => SERIAL_IN, DATA_IN(7) => 
                           DATA_IN_H(7), DATA_IN(6) => DATA_IN_H(6), DATA_IN(5)
                           => DATA_IN_H(5), DATA_IN(4) => DATA_IN_H(4), 
                           DATA_IN(3) => DATA_IN_H(3), DATA_IN(2) => 
                           DATA_IN_H(2), DATA_IN(1) => DATA_IN_H(1), DATA_IN(0)
                           => DATA_IN_H(0), BS_ERROR => BSE_H, CRC_ERROR => 
                           CRCE_H, EMPTY => EMPTY_H, FULL => FULL_H, KEY_ERROR 
                           => KEY_ERROR, PROG_ERROR => PROG_ERROR, PARITY_ERROR
                           => PARITY_ERROR, RBUF_FULL => n_1036, R_ERROR => 
                           RE_H, SENDING => host_is_sending, dm_tx_out => DMTS,
                           dp_tx_out => DPTS, W_ENABLE_R => W_ENABLE_H, 
                           R_ENABLE => R_ENABLE_H, DATA(7) => DATA_H(7), 
                           DATA(6) => DATA_H(6), DATA(5) => DATA_H(5), DATA(4) 
                           => DATA_H(4), DATA(3) => DATA_H(3), DATA(2) => 
                           DATA_H(2), DATA(1) => DATA_H(1), DATA(0) => 
                           DATA_H(0), ADDR(7) => ADDR_H(7), ADDR(6) => 
                           ADDR_H(6), ADDR(5) => ADDR_H(5), ADDR(4) => 
                           ADDR_H(4), ADDR(3) => ADDR_H(3), ADDR(2) => 
                           ADDR_H(2), ADDR(1) => ADDR_H(1), ADDR(0) => 
                           ADDR_H(0));
   U_1 : RMEDT_REWIRE_0 port map( CLK => CLK, DM1_RX => DMRS, DP1_RX => DPRS, 
                           RST => RST, SERIAL_IN => SERIAL_IN, DATA_IN(7) => 
                           DATA_IN_S(7), DATA_IN(6) => DATA_IN_S(6), DATA_IN(5)
                           => DATA_IN_S(5), DATA_IN(4) => DATA_IN_S(4), 
                           DATA_IN(3) => DATA_IN_S(3), DATA_IN(2) => 
                           DATA_IN_S(2), DATA_IN(1) => DATA_IN_S(1), DATA_IN(0)
                           => DATA_IN_S(0), BS_ERROR => BSE_S, CRC_ERROR => 
                           CRCE_S, EMPTY => EMPTY_S, FULL => FULL_S, KEY_ERROR 
                           => KEY_ERROR1, PROG_ERROR => PROG_ERROR1, 
                           PARITY_ERROR => PARITY_ERROR1, RBUF_FULL => n_1037, 
                           R_ERROR => RE_S, SENDING => slave_is_sending, 
                           dm_tx_out => DMTH, dp_tx_out => DPTH, W_ENABLE_R => 
                           W_ENABLE_S, R_ENABLE => R_ENABLE_S, DATA(7) => 
                           DATA_S(7), DATA(6) => DATA_S(6), DATA(5) => 
                           DATA_S(5), DATA(4) => DATA_S(4), DATA(3) => 
                           DATA_S(3), DATA(2) => DATA_S(2), DATA(1) => 
                           DATA_S(1), DATA(0) => DATA_S(0), ADDR(7) => 
                           ADDR_S(7), ADDR(6) => ADDR_S(6), ADDR(5) => 
                           ADDR_S(5), ADDR(4) => ADDR_S(4), ADDR(3) => 
                           ADDR_S(3), ADDR(2) => ADDR_S(2), ADDR(1) => 
                           ADDR_S(1), ADDR(0) => ADDR_S(0));

end SYN_struct;
