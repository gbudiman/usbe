
library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

package CONV_PACK_rmedt_square is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_rmedt_square;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_add_3 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_1_DW01_add_3;

architecture SYN_rpl of KSA_1_DW01_add_3 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n6, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : XOR2X1 port map( A => B(3), B => A(3), Y => n1);
   U2 : XOR2X1 port map( A => carry_3_port, B => n1, Y => SUM(3));
   U3 : NAND2X1 port map( A => carry_3_port, B => B(3), Y => n2);
   U4 : NAND2X1 port map( A => carry_3_port, B => A(3), Y => n3);
   U5 : NAND2X1 port map( A => B(3), B => A(3), Y => n4);
   U6 : NAND3X1 port map( A => n3, B => n2, C => n4, Y => carry_4_port);
   U7 : XOR2X1 port map( A => B(7), B => A(7), Y => n5);
   U8 : XOR2X1 port map( A => carry_7_port, B => n5, Y => SUM(7));
   U9 : AND2X2 port map( A => B(0), B => A(0), Y => n6);
   U10 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_add_2 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_1_DW01_add_2;

architecture SYN_rpl of KSA_1_DW01_add_2 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22 : std_logic;

begin
   
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => n22, YS
                           => SUM(7));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : XOR2X1 port map( A => A(5), B => B(5), Y => n2);
   U3 : XOR2X1 port map( A => n2, B => carry_5_port, Y => SUM(5));
   U4 : NAND2X1 port map( A => A(5), B => B(5), Y => n3);
   U5 : NAND2X1 port map( A => A(5), B => carry_5_port, Y => n4);
   U6 : NAND2X1 port map( A => B(5), B => carry_5_port, Y => n5);
   U7 : NAND3X1 port map( A => n3, B => n4, C => n5, Y => carry_6_port);
   U8 : XOR2X1 port map( A => A(6), B => B(6), Y => n6);
   U9 : XOR2X1 port map( A => n6, B => carry_6_port, Y => SUM(6));
   U10 : NAND2X1 port map( A => A(6), B => B(6), Y => n7);
   U11 : NAND2X1 port map( A => A(6), B => carry_6_port, Y => n8);
   U12 : NAND2X1 port map( A => B(6), B => carry_6_port, Y => n9);
   U13 : NAND3X1 port map( A => n7, B => n8, C => n9, Y => carry_7_port);
   U14 : XOR2X1 port map( A => B(1), B => A(1), Y => n10);
   U15 : XOR2X1 port map( A => n1, B => n10, Y => SUM(1));
   U16 : NAND2X1 port map( A => n1, B => B(1), Y => n11);
   U17 : NAND2X1 port map( A => n1, B => A(1), Y => n12);
   U18 : NAND2X1 port map( A => B(1), B => A(1), Y => n13);
   U19 : NAND3X1 port map( A => n12, B => n11, C => n13, Y => carry_2_port);
   U20 : XOR2X1 port map( A => A(2), B => B(2), Y => n14);
   U21 : XOR2X1 port map( A => n14, B => carry_2_port, Y => SUM(2));
   U22 : NAND2X1 port map( A => A(2), B => B(2), Y => n15);
   U23 : NAND2X1 port map( A => A(2), B => carry_2_port, Y => n16);
   U24 : NAND2X1 port map( A => B(2), B => carry_2_port, Y => n17);
   U25 : NAND3X1 port map( A => n15, B => n16, C => n17, Y => carry_3_port);
   U26 : XOR2X1 port map( A => A(3), B => B(3), Y => n18);
   U27 : XOR2X1 port map( A => n18, B => carry_3_port, Y => SUM(3));
   U28 : NAND2X1 port map( A => A(3), B => B(3), Y => n19);
   U29 : NAND2X1 port map( A => A(3), B => carry_3_port, Y => n20);
   U30 : NAND2X1 port map( A => B(3), B => carry_3_port, Y => n21);
   U31 : NAND3X1 port map( A => n19, B => n20, C => n21, Y => carry_4_port);
   U32 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_add_3 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_0_DW01_add_3;

architecture SYN_rpl of KSA_0_DW01_add_3 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n6, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : XOR2X1 port map( A => B(4), B => A(4), Y => n1);
   U2 : XOR2X1 port map( A => carry_4_port, B => n1, Y => SUM(4));
   U3 : NAND2X1 port map( A => carry_4_port, B => B(4), Y => n2);
   U4 : NAND2X1 port map( A => carry_4_port, B => A(4), Y => n3);
   U5 : NAND2X1 port map( A => B(4), B => A(4), Y => n4);
   U6 : NAND3X1 port map( A => n3, B => n2, C => n4, Y => carry_5_port);
   U7 : XOR2X1 port map( A => B(7), B => A(7), Y => n5);
   U8 : XOR2X1 port map( A => carry_7_port, B => n5, Y => SUM(7));
   U9 : AND2X2 port map( A => B(0), B => A(0), Y => n6);
   U10 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_add_2 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_0_DW01_add_2;

architecture SYN_rpl of KSA_0_DW01_add_2 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : 
      std_logic;

begin
   
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => n12, YS
                           => SUM(7));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n1, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : XOR2X1 port map( A => A(5), B => n10, Y => n2);
   U3 : XOR2X1 port map( A => n2, B => carry_5_port, Y => SUM(5));
   U4 : NAND2X1 port map( A => A(5), B => n10, Y => n3);
   U5 : NAND2X1 port map( A => A(5), B => carry_5_port, Y => n4);
   U6 : NAND2X1 port map( A => n10, B => carry_5_port, Y => n5);
   U7 : NAND3X1 port map( A => n3, B => n4, C => n5, Y => carry_6_port);
   U8 : XOR2X1 port map( A => A(6), B => n11, Y => n6);
   U9 : XOR2X1 port map( A => n6, B => carry_6_port, Y => SUM(6));
   U10 : NAND2X1 port map( A => A(6), B => n11, Y => n7);
   U11 : NAND2X1 port map( A => A(6), B => carry_6_port, Y => n8);
   U12 : NAND2X1 port map( A => n11, B => carry_6_port, Y => n9);
   U13 : NAND3X1 port map( A => n7, B => n8, C => n9, Y => carry_7_port);
   U14 : BUFX2 port map( A => B(5), Y => n10);
   U15 : BUFX2 port map( A => B(6), Y => n11);
   U16 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_inc_2 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_1_DW01_inc_2;

architecture SYN_rpl of KSA_1_DW01_inc_2 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_inc_1 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_1_DW01_inc_1;

architecture SYN_rpl of KSA_1_DW01_inc_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_1_DW01_inc_0;

architecture SYN_rpl of KSA_1_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_add_1 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_1_DW01_add_1;

architecture SYN_rpl of KSA_1_DW01_add_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2 : std_logic;

begin
   
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => n2, YS 
                           => SUM(7));
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n1, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1_DW01_add_0 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_1_DW01_add_0;

architecture SYN_rpl of KSA_1_DW01_add_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2 : std_logic;

begin
   
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => n2, YS 
                           => SUM(7));
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n1, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity keyreg_1_DW01_add_0 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end keyreg_1_DW01_add_0;

architecture SYN_rpl of keyreg_1_DW01_add_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => n10, YS
                           => SUM(7));
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n9, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : XOR2X1 port map( A => A(3), B => B(3), Y => n1);
   U2 : XOR2X1 port map( A => n1, B => carry_3_port, Y => SUM(3));
   U3 : NAND2X1 port map( A => A(3), B => B(3), Y => n2);
   U4 : NAND2X1 port map( A => A(3), B => carry_3_port, Y => n3);
   U5 : NAND2X1 port map( A => B(3), B => carry_3_port, Y => n4);
   U6 : NAND3X1 port map( A => n2, B => n3, C => n4, Y => carry_4_port);
   U7 : XOR2X1 port map( A => A(4), B => B(4), Y => n5);
   U8 : XOR2X1 port map( A => n5, B => carry_4_port, Y => SUM(4));
   U9 : NAND2X1 port map( A => A(4), B => B(4), Y => n6);
   U10 : NAND2X1 port map( A => A(4), B => carry_4_port, Y => n7);
   U11 : NAND2X1 port map( A => B(4), B => carry_4_port, Y => n8);
   U12 : NAND3X1 port map( A => n6, B => n7, C => n8, Y => carry_5_port);
   U13 : AND2X2 port map( A => B(0), B => A(0), Y => n9);
   U14 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_timer_1_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end uart_timer_1_DW01_inc_0;

architecture SYN_rpl of uart_timer_1_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_tcu_1_DW01_inc_0 is

   port( A : in std_logic_vector (6 downto 0);  SUM : out std_logic_vector (6 
         downto 0));

end tx_tcu_1_DW01_inc_0;

architecture SYN_rpl of tx_tcu_1_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port 
      : std_logic;

begin
   
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_6_port, B => A(6), Y => SUM(6));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_inc_2 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_0_DW01_inc_2;

architecture SYN_rpl of KSA_0_DW01_inc_2 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_inc_1 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_0_DW01_inc_1;

architecture SYN_rpl of KSA_0_DW01_inc_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end KSA_0_DW01_inc_0;

architecture SYN_rpl of KSA_0_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_add_1 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_0_DW01_add_1;

architecture SYN_rpl of KSA_0_DW01_add_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2 : std_logic;

begin
   
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => n2, YS 
                           => SUM(7));
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n1, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0_DW01_add_0 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end KSA_0_DW01_add_0;

architecture SYN_rpl of KSA_0_DW01_add_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2 : std_logic;

begin
   
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => n2, YS 
                           => SUM(7));
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n1, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity keyreg_0_DW01_add_0 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end keyreg_0_DW01_add_0;

architecture SYN_rpl of keyreg_0_DW01_add_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, n1, n2 : std_logic;

begin
   
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => n2, YS 
                           => SUM(7));
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n1, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_timer_0_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end uart_timer_0_DW01_inc_0;

architecture SYN_rpl of uart_timer_0_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_tcu_0_DW01_inc_0 is

   port( A : in std_logic_vector (6 downto 0);  SUM : out std_logic_vector (6 
         downto 0));

end tx_tcu_0_DW01_inc_0;

architecture SYN_rpl of tx_tcu_0_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port 
      : std_logic;

begin
   
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_6_port, B => A(6), Y => SUM(6));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_timer_0 is

   port( CLK, RST, TIMER_TRIG : in std_logic;  STOP_RCVING, SHIFT_STROBE : out 
         std_logic);

end uart_timer_0;

architecture SYN_timerB of uart_timer_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component uart_timer_0_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal state_7_port, state_6_port, state_5_port, state_4_port, state_3_port,
      state_2_port, state_1_port, state_0_port, nextState_7_port, 
      nextState_6_port, nextState_5_port, nextState_4_port, nextState_3_port, 
      nextState_2_port, nextState_1_port, nextState_0_port, N26, N27, N28, N29,
      N30, N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26_port
      , n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110 : std_logic;

begin
   
   U21 : OR2X2 port map( A => state_7_port, B => n95, Y => n96);
   U38 : OAI21X1 port map( A => n20, B => n27_port, C => n110, Y => n81);
   U39 : NAND2X1 port map( A => N33, B => n109, Y => n110);
   U40 : OAI21X1 port map( A => n26_port, B => n20, C => n108, Y => n80);
   U41 : NAND2X1 port map( A => N32, B => n109, Y => n108);
   U42 : OAI21X1 port map( A => n25, B => n20, C => n107, Y => n79);
   U43 : NAND2X1 port map( A => N31, B => n109, Y => n107);
   U44 : OAI21X1 port map( A => n20, B => n24, C => n106, Y => n78);
   U45 : NAND2X1 port map( A => N30, B => n109, Y => n106);
   U46 : OAI21X1 port map( A => n23, B => n20, C => n105, Y => n77);
   U47 : NAND2X1 port map( A => N29, B => n109, Y => n105);
   U48 : OAI21X1 port map( A => n22, B => n20, C => n104, Y => n76);
   U49 : NAND2X1 port map( A => N28, B => n109, Y => n104);
   U50 : OAI21X1 port map( A => n20, B => n21, C => n103, Y => n75);
   U51 : NAND2X1 port map( A => N27, B => n109, Y => n103);
   U52 : OAI21X1 port map( A => n19, B => n20, C => n102, Y => n74);
   U53 : NAND2X1 port map( A => N26, B => n109, Y => n102);
   U54 : NOR2X1 port map( A => n101, B => n73, Y => n109);
   U55 : NOR2X1 port map( A => n73, B => TIMER_TRIG, Y => n101);
   U56 : NOR2X1 port map( A => n100, B => n99, Y => n73);
   U57 : NAND3X1 port map( A => nextState_6_port, B => nextState_5_port, C => 
                           n98, Y => n99);
   U58 : NOR2X1 port map( A => n22, B => n23, Y => n98);
   U59 : NAND3X1 port map( A => nextState_0_port, B => n21, C => n97, Y => n100
                           );
   U60 : NOR2X1 port map( A => nextState_7_port, B => nextState_4_port, Y => 
                           n97);
   U61 : NOR2X1 port map( A => state_0_port, B => n96, Y => SHIFT_STROBE);
   U62 : AOI21X1 port map( A => n94, B => n32_port, C => n93, Y => n95);
   U63 : OAI21X1 port map( A => n33_port, B => n92, C => n91, Y => n93);
   U64 : NAND3X1 port map( A => state_6_port, B => state_1_port, C => n90, Y =>
                           n91);
   U65 : AOI21X1 port map( A => n89, B => n88, C => state_3_port, Y => n90);
   U66 : NAND3X1 port map( A => n33_port, B => n31_port, C => state_4_port, Y 
                           => n88);
   U67 : NAND3X1 port map( A => state_2_port, B => n32_port, C => state_5_port,
                           Y => n89);
   U68 : NAND2X1 port map( A => state_4_port, B => n87, Y => n92);
   U69 : OAI21X1 port map( A => state_2_port, B => n28_port, C => n86, Y => n94
                           );
   U70 : NAND3X1 port map( A => state_2_port, B => n29_port, C => n30_port, Y 
                           => n86);
   U71 : OAI22X1 port map( A => state_6_port, B => n84, C => n29_port, D => n85
                           , Y => n87);
   U72 : NAND3X1 port map( A => n34, B => n31_port, C => state_3_port, Y => n85
                           );
   U73 : AOI22X1 port map( A => n83, B => state_1_port, C => n82, D => 
                           state_5_port, Y => n84);
   U74 : XOR2X1 port map( A => n34, B => state_3_port, Y => n82);
   U75 : NOR2X1 port map( A => state_5_port, B => state_3_port, Y => n83);
   add_39 : uart_timer_0_DW01_inc_0 port map( A(7) => nextState_7_port, A(6) =>
                           nextState_6_port, A(5) => nextState_5_port, A(4) => 
                           nextState_4_port, A(3) => nextState_3_port, A(2) => 
                           nextState_2_port, A(1) => nextState_1_port, A(0) => 
                           nextState_0_port, SUM(7) => N33, SUM(6) => N32, 
                           SUM(5) => N31, SUM(4) => N30, SUM(3) => N29, SUM(2) 
                           => N28, SUM(1) => N27, SUM(0) => N26);
   state_reg_3_inst : DFFSR port map( D => nextState_3_port, CLK => CLK, R => 
                           n18, S => n17, Q => state_3_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n18, S => n16, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n18, S => n15, Q => state_1_port);
   state_reg_5_inst : DFFSR port map( D => nextState_5_port, CLK => CLK, R => 
                           n18, S => n14, Q => state_5_port);
   state_reg_6_inst : DFFSR port map( D => nextState_6_port, CLK => CLK, R => 
                           n18, S => n13, Q => state_6_port);
   state_reg_4_inst : DFFSR port map( D => nextState_4_port, CLK => CLK, R => 
                           n18, S => n12, Q => state_4_port);
   state_reg_7_inst : DFFSR port map( D => nextState_7_port, CLK => CLK, R => 
                           n18, S => n11, Q => state_7_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n18, S => n10, Q => state_0_port);
   STOP_RCVING_reg : DFFSR port map( D => n73, CLK => CLK, R => n18, S => n9, Q
                           => STOP_RCVING);
   nextState_reg_3_inst : DFFSR port map( D => n77, CLK => CLK, R => n18, S => 
                           n8, Q => nextState_3_port);
   nextState_reg_2_inst : DFFSR port map( D => n76, CLK => CLK, R => n18, S => 
                           n7, Q => nextState_2_port);
   nextState_reg_0_inst : DFFSR port map( D => n74, CLK => CLK, R => n18, S => 
                           n6, Q => nextState_0_port);
   nextState_reg_4_inst : DFFSR port map( D => n78, CLK => CLK, R => n18, S => 
                           n5, Q => nextState_4_port);
   nextState_reg_1_inst : DFFSR port map( D => n75, CLK => CLK, R => n18, S => 
                           n4, Q => nextState_1_port);
   nextState_reg_5_inst : DFFSR port map( D => n79, CLK => CLK, R => n18, S => 
                           n3, Q => nextState_5_port);
   nextState_reg_6_inst : DFFSR port map( D => n80, CLK => CLK, R => n18, S => 
                           n2, Q => nextState_6_port);
   nextState_reg_7_inst : DFFSR port map( D => n81, CLK => CLK, R => n18, S => 
                           n1, Q => nextState_7_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   U20 : INVX2 port map( A => RST, Y => n18);
   U22 : INVX2 port map( A => nextState_0_port, Y => n19);
   U23 : INVX2 port map( A => n101, Y => n20);
   U24 : INVX2 port map( A => nextState_1_port, Y => n21);
   U25 : INVX2 port map( A => nextState_2_port, Y => n22);
   U26 : INVX2 port map( A => nextState_3_port, Y => n23);
   U27 : INVX2 port map( A => nextState_4_port, Y => n24);
   U28 : INVX2 port map( A => nextState_5_port, Y => n25);
   U29 : INVX2 port map( A => nextState_6_port, Y => n26_port);
   U30 : INVX2 port map( A => nextState_7_port, Y => n27_port);
   U31 : INVX2 port map( A => n87, Y => n28_port);
   U32 : INVX2 port map( A => state_6_port, Y => n29_port);
   U33 : INVX2 port map( A => n85, Y => n30_port);
   U34 : INVX2 port map( A => state_5_port, Y => n31_port);
   U35 : INVX2 port map( A => state_4_port, Y => n32_port);
   U36 : INVX2 port map( A => state_2_port, Y => n33_port);
   U37 : INVX2 port map( A => state_1_port, Y => n34);

end SYN_timerB;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity keyreg_0 is

   port( CLK, RST, SBE, OE, RBUF_FULL : in std_logic;  RCV_DATA : in 
         std_logic_vector (7 downto 0);  PLAINKEY : out std_logic_vector (63 
         downto 0);  KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR : out 
         std_logic);

end keyreg_0;

architecture SYN_keyb of keyreg_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component keyreg_0_DW01_add_0
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port, 
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port, CLR_RBUFF_port, state_3_port, state_2_port, state_1_port
      , state_0_port, parityError, keyCount_3_port, keyCount_2_port, 
      keyCount_1_port, keyCount_0_port, address_7_port, address_6_port, 
      address_5_port, address_4_port, address_3_port, address_2_port, 
      address_1_port, address_0_port, currentPlainKey_63_port, 
      currentPlainKey_62_port, currentPlainKey_61_port, currentPlainKey_60_port
      , currentPlainKey_59_port, currentPlainKey_58_port, 
      currentPlainKey_57_port, currentPlainKey_56_port, currentPlainKey_55_port
      , currentPlainKey_54_port, currentPlainKey_53_port, 
      currentPlainKey_52_port, currentPlainKey_51_port, currentPlainKey_50_port
      , currentPlainKey_49_port, currentPlainKey_48_port, 
      currentPlainKey_47_port, currentPlainKey_46_port, currentPlainKey_45_port
      , currentPlainKey_44_port, currentPlainKey_43_port, 
      currentPlainKey_42_port, currentPlainKey_41_port, currentPlainKey_40_port
      , currentPlainKey_39_port, currentPlainKey_38_port, 
      currentPlainKey_37_port, currentPlainKey_36_port, currentPlainKey_35_port
      , currentPlainKey_34_port, currentPlainKey_33_port, 
      currentPlainKey_32_port, currentPlainKey_31_port, currentPlainKey_30_port
      , currentPlainKey_29_port, currentPlainKey_28_port, 
      currentPlainKey_27_port, currentPlainKey_26_port, currentPlainKey_25_port
      , currentPlainKey_24_port, currentPlainKey_23_port, 
      currentPlainKey_22_port, currentPlainKey_21_port, currentPlainKey_20_port
      , currentPlainKey_19_port, currentPlainKey_18_port, 
      currentPlainKey_17_port, currentPlainKey_16_port, currentPlainKey_15_port
      , currentPlainKey_14_port, currentPlainKey_13_port, 
      currentPlainKey_12_port, currentPlainKey_11_port, currentPlainKey_10_port
      , currentPlainKey_9_port, currentPlainKey_8_port, currentPlainKey_7_port,
      currentPlainKey_6_port, currentPlainKey_5_port, currentPlainKey_4_port, 
      currentPlainKey_3_port, currentPlainKey_2_port, currentPlainKey_1_port, 
      currentPlainKey_0_port, parityAccumulator_7_port, 
      parityAccumulator_6_port, parityAccumulator_5_port, 
      parityAccumulator_4_port, parityAccumulator_3_port, 
      parityAccumulator_2_port, parityAccumulator_1_port, 
      parityAccumulator_0_port, nextParityError, N694, N1792, N1793, N1794, 
      N1795, N1796, N1797, N1798, N1799, n1, n2, n4, n5, n6, n7, n8, n9, n10, 
      n11, n14, n16, n17, n19, n20, n21, n23, n25, n27, n29, n31, n33, n35, n37
      , n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63, n65, 
      n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95
      , n97, n99, n101, n103, n105, n107, n109, n111, n113, n115, n117, n119, 
      n121, n123, n125, n127, n129, n131, n133, n135, n137, n139, n141, n143, 
      n145, n147, n149, n150, n151, n153, n154, n156, n158, n160, n161, n165, 
      n166, n168, n172, n173, n175, n177, n178, n180, n181, n183, n184, n185, 
      n186, n187, n188, n189, n192, n193, n195, n197, n203, n205, n206, n207, 
      n208, n209, n210, n217, n219, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n240, n241, n242, n243, n244, 
      n245, n247, n248, n249, n250, n255, n257, n258, n259, n260, n261, n262, 
      n263, n264, n265, n266, n267, n268, n269, n270, n271, n275, n277, n278, 
      n279, n280, n281, n282, n284, n285, n286, n287, n289, n291, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n311, n312, n313, 
      n314, n315, n316, n317, n319, n320, n321, n322, n324, n326, n327, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n343, n344, 
      n345, n346, n347, n348, n350, n351, n352, n353, n355, n357, n360, n361, 
      n362, n363, n364, n365, n366, n367, n368, n369, n370, n373, n374, n375, 
      n376, n377, n378, n380, n381, n382, n383, n385, n387, n390, n391, n392, 
      n393, n394, n395, n396, n397, n398, n399, n400, n404, n405, n406, n407, 
      n408, n409, n411, n412, n413, n414, n416, n418, n419, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n435, n436, n437, n438, 
      n439, n440, n441, n443, n444, n445, n446, n448, n450, n452, n453, n454, 
      n455, n456, n457, n458, n459, n460, n461, n462, n465, n466, n467, n468, 
      n469, n471, n472, n473, n474, n476, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n492, n493, n494, n495, n496, n498, n499, 
      n500, n501, n503, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n519, n520, n521, n522, n523, n525, n526, n527, n528, n530, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n547, 
      n548, n549, n550, n551, n552, n554, n555, n556, n557, n559, n561, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n576, n577, 
      n578, n579, n580, n582, n583, n584, n585, n587, n590, n591, n592, n593, 
      n594, n595, n596, n597, n598, n599, n600, n603, n604, n605, n606, n607, 
      n609, n610, n611, n612, n614, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n630, n631, n632, n633, n634, n636, n637, n638, 
      n639, n641, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, 
      n654, n657, n658, n659, n660, n661, n662, n663, n665, n666, n667, n668, 
      n670, n672, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n687, n688, n689, n690, n691, n693, n694_port, n695, n696, n698, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n714, 
      n715, n716, n717, n718, n720, n721, n722, n723, n725, n728, n729, n730, 
      n731, n732, n733, n734, n735, n736, n737, n738, n741, n742, n743, n744, 
      n745, n747, n748, n749, n750, n752, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n769, n770, n771, n772, n773, n774, n776, 
      n777, n778, n779, n781, n783, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n798, n799, n800, n801, n802, n804, n805, n806, 
      n807, n809, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, 
      n822, n825, n826, n827, n828, n829, n831, n832, n833, n834, n836, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n852, n853, 
      n854, n855, n856, n858, n859, n860, n861, n863, n866, n867, n868, n869, 
      n870, n871, n872, n873, n874, n875, n876, n879, n880, n881, n882, n883, 
      n884, n885, n887, n888, n889, n890, n892, n894, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n909, n910, n911, n912, n913, 
      n915, n916, n917, n918, n920, n923, n924, n925, n926, n927, n928, n929, 
      n930, n931, n932, n933, n936, n937, n938, n939, n940, n942, n943, n944, 
      n945, n947, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n963, n964, n965, n966, n967, n969, n970, n971, n972, n974, n977, 
      n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1003, n1005, 
      n1007, n1008, n1009, n1010, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1032, n1035, n1036, n1037, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, 
      n1056, n1057, n1058, n1059, n1060, n1061, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1091, 
      n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1102, 
      n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, 
      n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, 
      n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, 
      n1139, n1140, n1141, n1142, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1161, 
      n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, 
      n1172, n1173, n1174, n1175, n1176, n1177, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
      n1268, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, PROG_ERROR_port, n1482, n1483, n1484, 
      n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
      n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, 
      n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, 
      n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
      n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, 
      n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, 
      n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, 
      n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, 
      n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, 
      n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, 
      n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, 
      n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, 
      n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, 
      n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, 
      n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, 
      n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, 
      n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, 
      n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, 
      n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, 
      n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, 
      n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
      n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
      n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 
      n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, 
      n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, 
      n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, 
      n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
      n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, 
      n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
      n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, 
      n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792_port, n1793_port, 
      n1794_port, n1795_port, n1796_port, n1797_port, n1798_port, n1799_port, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, 
      n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
      n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
      n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, 
      n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
      n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
      n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, 
      n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
      n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n_1020 : 
      std_logic;

begin
   PLAINKEY <= ( PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port, 
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port );
   PROG_ERROR <= PROG_ERROR_port;
   CLR_RBUFF <= CLR_RBUFF_port;
   
   n2038 <= '0';
   keyCount_reg_0_inst : DFFPOSX1 port map( D => n1577, CLK => CLK, Q => 
                           keyCount_0_port);
   keyCount_reg_2_inst : DFFPOSX1 port map( D => n1584, CLK => CLK, Q => 
                           keyCount_2_port);
   keyCount_reg_3_inst : DFFPOSX1 port map( D => n1578, CLK => CLK, Q => 
                           keyCount_3_port);
   parityAccumulator_reg_0_inst : DFFPOSX1 port map( D => n1585, CLK => CLK, Q 
                           => parityAccumulator_0_port);
   parityAccumulator_reg_1_inst : DFFPOSX1 port map( D => n1586, CLK => CLK, Q 
                           => parityAccumulator_1_port);
   parityAccumulator_reg_2_inst : DFFPOSX1 port map( D => n1587, CLK => CLK, Q 
                           => parityAccumulator_2_port);
   parityAccumulator_reg_3_inst : DFFPOSX1 port map( D => n1588, CLK => CLK, Q 
                           => parityAccumulator_3_port);
   parityAccumulator_reg_4_inst : DFFPOSX1 port map( D => n1589, CLK => CLK, Q 
                           => parityAccumulator_4_port);
   parityAccumulator_reg_5_inst : DFFPOSX1 port map( D => n1590, CLK => CLK, Q 
                           => parityAccumulator_5_port);
   parityAccumulator_reg_6_inst : DFFPOSX1 port map( D => n1591, CLK => CLK, Q 
                           => parityAccumulator_6_port);
   parityAccumulator_reg_7_inst : DFFPOSX1 port map( D => n1592, CLK => CLK, Q 
                           => parityAccumulator_7_port);
   keyCount_reg_1_inst : DFFPOSX1 port map( D => n1583, CLK => CLK, Q => 
                           keyCount_1_port);
   address_reg_7_inst : DFFPOSX1 port map( D => n1593, CLK => CLK, Q => 
                           address_7_port);
   address_reg_6_inst : DFFPOSX1 port map( D => n1594, CLK => CLK, Q => 
                           address_6_port);
   address_reg_5_inst : DFFPOSX1 port map( D => n1595, CLK => CLK, Q => 
                           address_5_port);
   address_reg_4_inst : DFFPOSX1 port map( D => n1596, CLK => CLK, Q => 
                           address_4_port);
   address_reg_3_inst : DFFPOSX1 port map( D => n1597, CLK => CLK, Q => 
                           address_3_port);
   address_reg_2_inst : DFFPOSX1 port map( D => n1598, CLK => CLK, Q => 
                           address_2_port);
   address_reg_1_inst : DFFPOSX1 port map( D => n1599, CLK => CLK, Q => 
                           address_1_port);
   address_reg_0_inst : DFFPOSX1 port map( D => n1600, CLK => CLK, Q => 
                           address_0_port);
   currentPlainKey_reg_63_inst : DFFPOSX1 port map( D => n1664, CLK => CLK, Q 
                           => currentPlainKey_63_port);
   currentPlainKey_reg_62_inst : DFFPOSX1 port map( D => n1663, CLK => CLK, Q 
                           => currentPlainKey_62_port);
   currentPlainKey_reg_61_inst : DFFPOSX1 port map( D => n1662, CLK => CLK, Q 
                           => currentPlainKey_61_port);
   currentPlainKey_reg_60_inst : DFFPOSX1 port map( D => n1661, CLK => CLK, Q 
                           => currentPlainKey_60_port);
   currentPlainKey_reg_59_inst : DFFPOSX1 port map( D => n1660, CLK => CLK, Q 
                           => currentPlainKey_59_port);
   currentPlainKey_reg_58_inst : DFFPOSX1 port map( D => n1659, CLK => CLK, Q 
                           => currentPlainKey_58_port);
   currentPlainKey_reg_57_inst : DFFPOSX1 port map( D => n1658, CLK => CLK, Q 
                           => currentPlainKey_57_port);
   currentPlainKey_reg_56_inst : DFFPOSX1 port map( D => n1657, CLK => CLK, Q 
                           => currentPlainKey_56_port);
   currentPlainKey_reg_55_inst : DFFPOSX1 port map( D => n1656, CLK => CLK, Q 
                           => currentPlainKey_55_port);
   currentPlainKey_reg_54_inst : DFFPOSX1 port map( D => n1655, CLK => CLK, Q 
                           => currentPlainKey_54_port);
   currentPlainKey_reg_53_inst : DFFPOSX1 port map( D => n1654, CLK => CLK, Q 
                           => currentPlainKey_53_port);
   currentPlainKey_reg_52_inst : DFFPOSX1 port map( D => n1653, CLK => CLK, Q 
                           => currentPlainKey_52_port);
   currentPlainKey_reg_51_inst : DFFPOSX1 port map( D => n1652, CLK => CLK, Q 
                           => currentPlainKey_51_port);
   currentPlainKey_reg_50_inst : DFFPOSX1 port map( D => n1651, CLK => CLK, Q 
                           => currentPlainKey_50_port);
   currentPlainKey_reg_49_inst : DFFPOSX1 port map( D => n1650, CLK => CLK, Q 
                           => currentPlainKey_49_port);
   currentPlainKey_reg_48_inst : DFFPOSX1 port map( D => n1649, CLK => CLK, Q 
                           => currentPlainKey_48_port);
   currentPlainKey_reg_47_inst : DFFPOSX1 port map( D => n1648, CLK => CLK, Q 
                           => currentPlainKey_47_port);
   currentPlainKey_reg_46_inst : DFFPOSX1 port map( D => n1647, CLK => CLK, Q 
                           => currentPlainKey_46_port);
   currentPlainKey_reg_45_inst : DFFPOSX1 port map( D => n1646, CLK => CLK, Q 
                           => currentPlainKey_45_port);
   currentPlainKey_reg_44_inst : DFFPOSX1 port map( D => n1645, CLK => CLK, Q 
                           => currentPlainKey_44_port);
   currentPlainKey_reg_43_inst : DFFPOSX1 port map( D => n1644, CLK => CLK, Q 
                           => currentPlainKey_43_port);
   currentPlainKey_reg_42_inst : DFFPOSX1 port map( D => n1643, CLK => CLK, Q 
                           => currentPlainKey_42_port);
   currentPlainKey_reg_41_inst : DFFPOSX1 port map( D => n1642, CLK => CLK, Q 
                           => currentPlainKey_41_port);
   currentPlainKey_reg_40_inst : DFFPOSX1 port map( D => n1641, CLK => CLK, Q 
                           => currentPlainKey_40_port);
   currentPlainKey_reg_39_inst : DFFPOSX1 port map( D => n1640, CLK => CLK, Q 
                           => currentPlainKey_39_port);
   currentPlainKey_reg_38_inst : DFFPOSX1 port map( D => n1639, CLK => CLK, Q 
                           => currentPlainKey_38_port);
   currentPlainKey_reg_37_inst : DFFPOSX1 port map( D => n1638, CLK => CLK, Q 
                           => currentPlainKey_37_port);
   currentPlainKey_reg_36_inst : DFFPOSX1 port map( D => n1637, CLK => CLK, Q 
                           => currentPlainKey_36_port);
   currentPlainKey_reg_35_inst : DFFPOSX1 port map( D => n1636, CLK => CLK, Q 
                           => currentPlainKey_35_port);
   currentPlainKey_reg_34_inst : DFFPOSX1 port map( D => n1635, CLK => CLK, Q 
                           => currentPlainKey_34_port);
   currentPlainKey_reg_33_inst : DFFPOSX1 port map( D => n1634, CLK => CLK, Q 
                           => currentPlainKey_33_port);
   currentPlainKey_reg_32_inst : DFFPOSX1 port map( D => n1633, CLK => CLK, Q 
                           => currentPlainKey_32_port);
   currentPlainKey_reg_31_inst : DFFPOSX1 port map( D => n1632, CLK => CLK, Q 
                           => currentPlainKey_31_port);
   currentPlainKey_reg_30_inst : DFFPOSX1 port map( D => n1631, CLK => CLK, Q 
                           => currentPlainKey_30_port);
   currentPlainKey_reg_29_inst : DFFPOSX1 port map( D => n1630, CLK => CLK, Q 
                           => currentPlainKey_29_port);
   currentPlainKey_reg_28_inst : DFFPOSX1 port map( D => n1629, CLK => CLK, Q 
                           => currentPlainKey_28_port);
   currentPlainKey_reg_27_inst : DFFPOSX1 port map( D => n1628, CLK => CLK, Q 
                           => currentPlainKey_27_port);
   currentPlainKey_reg_26_inst : DFFPOSX1 port map( D => n1627, CLK => CLK, Q 
                           => currentPlainKey_26_port);
   currentPlainKey_reg_25_inst : DFFPOSX1 port map( D => n1626, CLK => CLK, Q 
                           => currentPlainKey_25_port);
   currentPlainKey_reg_24_inst : DFFPOSX1 port map( D => n1625, CLK => CLK, Q 
                           => currentPlainKey_24_port);
   currentPlainKey_reg_23_inst : DFFPOSX1 port map( D => n1624, CLK => CLK, Q 
                           => currentPlainKey_23_port);
   currentPlainKey_reg_22_inst : DFFPOSX1 port map( D => n1623, CLK => CLK, Q 
                           => currentPlainKey_22_port);
   currentPlainKey_reg_21_inst : DFFPOSX1 port map( D => n1622, CLK => CLK, Q 
                           => currentPlainKey_21_port);
   currentPlainKey_reg_20_inst : DFFPOSX1 port map( D => n1621, CLK => CLK, Q 
                           => currentPlainKey_20_port);
   currentPlainKey_reg_19_inst : DFFPOSX1 port map( D => n1620, CLK => CLK, Q 
                           => currentPlainKey_19_port);
   currentPlainKey_reg_18_inst : DFFPOSX1 port map( D => n1619, CLK => CLK, Q 
                           => currentPlainKey_18_port);
   currentPlainKey_reg_17_inst : DFFPOSX1 port map( D => n1618, CLK => CLK, Q 
                           => currentPlainKey_17_port);
   currentPlainKey_reg_16_inst : DFFPOSX1 port map( D => n1617, CLK => CLK, Q 
                           => currentPlainKey_16_port);
   currentPlainKey_reg_15_inst : DFFPOSX1 port map( D => n1616, CLK => CLK, Q 
                           => currentPlainKey_15_port);
   currentPlainKey_reg_14_inst : DFFPOSX1 port map( D => n1615, CLK => CLK, Q 
                           => currentPlainKey_14_port);
   currentPlainKey_reg_13_inst : DFFPOSX1 port map( D => n1614, CLK => CLK, Q 
                           => currentPlainKey_13_port);
   currentPlainKey_reg_12_inst : DFFPOSX1 port map( D => n1613, CLK => CLK, Q 
                           => currentPlainKey_12_port);
   currentPlainKey_reg_11_inst : DFFPOSX1 port map( D => n1612, CLK => CLK, Q 
                           => currentPlainKey_11_port);
   currentPlainKey_reg_10_inst : DFFPOSX1 port map( D => n1611, CLK => CLK, Q 
                           => currentPlainKey_10_port);
   currentPlainKey_reg_9_inst : DFFPOSX1 port map( D => n1610, CLK => CLK, Q =>
                           currentPlainKey_9_port);
   currentPlainKey_reg_8_inst : DFFPOSX1 port map( D => n1609, CLK => CLK, Q =>
                           currentPlainKey_8_port);
   currentPlainKey_reg_7_inst : DFFPOSX1 port map( D => n1608, CLK => CLK, Q =>
                           currentPlainKey_7_port);
   currentPlainKey_reg_6_inst : DFFPOSX1 port map( D => n1607, CLK => CLK, Q =>
                           currentPlainKey_6_port);
   currentPlainKey_reg_5_inst : DFFPOSX1 port map( D => n1606, CLK => CLK, Q =>
                           currentPlainKey_5_port);
   currentPlainKey_reg_4_inst : DFFPOSX1 port map( D => n1605, CLK => CLK, Q =>
                           currentPlainKey_4_port);
   currentPlainKey_reg_3_inst : DFFPOSX1 port map( D => n1604, CLK => CLK, Q =>
                           currentPlainKey_3_port);
   currentPlainKey_reg_2_inst : DFFPOSX1 port map( D => n1603, CLK => CLK, Q =>
                           currentPlainKey_2_port);
   currentPlainKey_reg_1_inst : DFFPOSX1 port map( D => n1602, CLK => CLK, Q =>
                           currentPlainKey_1_port);
   currentPlainKey_reg_0_inst : DFFPOSX1 port map( D => n1601, CLK => CLK, Q =>
                           currentPlainKey_0_port);
   PLAINKEY_reg_63_inst : DFFPOSX1 port map( D => n1665, CLK => CLK, Q => 
                           PLAINKEY_63_port);
   PLAINKEY_reg_62_inst : DFFPOSX1 port map( D => n1666, CLK => CLK, Q => 
                           PLAINKEY_62_port);
   PLAINKEY_reg_61_inst : DFFPOSX1 port map( D => n1667, CLK => CLK, Q => 
                           PLAINKEY_61_port);
   PLAINKEY_reg_60_inst : DFFPOSX1 port map( D => n1668, CLK => CLK, Q => 
                           PLAINKEY_60_port);
   PLAINKEY_reg_59_inst : DFFPOSX1 port map( D => n1669, CLK => CLK, Q => 
                           PLAINKEY_59_port);
   PLAINKEY_reg_58_inst : DFFPOSX1 port map( D => n1670, CLK => CLK, Q => 
                           PLAINKEY_58_port);
   PLAINKEY_reg_57_inst : DFFPOSX1 port map( D => n1671, CLK => CLK, Q => 
                           PLAINKEY_57_port);
   PLAINKEY_reg_56_inst : DFFPOSX1 port map( D => n1672, CLK => CLK, Q => 
                           PLAINKEY_56_port);
   PLAINKEY_reg_55_inst : DFFPOSX1 port map( D => n1673, CLK => CLK, Q => 
                           PLAINKEY_55_port);
   PLAINKEY_reg_54_inst : DFFPOSX1 port map( D => n1674, CLK => CLK, Q => 
                           PLAINKEY_54_port);
   PLAINKEY_reg_53_inst : DFFPOSX1 port map( D => n1675, CLK => CLK, Q => 
                           PLAINKEY_53_port);
   PLAINKEY_reg_52_inst : DFFPOSX1 port map( D => n1676, CLK => CLK, Q => 
                           PLAINKEY_52_port);
   PLAINKEY_reg_51_inst : DFFPOSX1 port map( D => n1677, CLK => CLK, Q => 
                           PLAINKEY_51_port);
   PLAINKEY_reg_50_inst : DFFPOSX1 port map( D => n1678, CLK => CLK, Q => 
                           PLAINKEY_50_port);
   PLAINKEY_reg_49_inst : DFFPOSX1 port map( D => n1679, CLK => CLK, Q => 
                           PLAINKEY_49_port);
   PLAINKEY_reg_48_inst : DFFPOSX1 port map( D => n1680, CLK => CLK, Q => 
                           PLAINKEY_48_port);
   PLAINKEY_reg_47_inst : DFFPOSX1 port map( D => n1681, CLK => CLK, Q => 
                           PLAINKEY_47_port);
   PLAINKEY_reg_46_inst : DFFPOSX1 port map( D => n1682, CLK => CLK, Q => 
                           PLAINKEY_46_port);
   PLAINKEY_reg_45_inst : DFFPOSX1 port map( D => n1683, CLK => CLK, Q => 
                           PLAINKEY_45_port);
   PLAINKEY_reg_44_inst : DFFPOSX1 port map( D => n1684, CLK => CLK, Q => 
                           PLAINKEY_44_port);
   PLAINKEY_reg_43_inst : DFFPOSX1 port map( D => n1685, CLK => CLK, Q => 
                           PLAINKEY_43_port);
   PLAINKEY_reg_42_inst : DFFPOSX1 port map( D => n1686, CLK => CLK, Q => 
                           PLAINKEY_42_port);
   PLAINKEY_reg_41_inst : DFFPOSX1 port map( D => n1687, CLK => CLK, Q => 
                           PLAINKEY_41_port);
   PLAINKEY_reg_40_inst : DFFPOSX1 port map( D => n1688, CLK => CLK, Q => 
                           PLAINKEY_40_port);
   PLAINKEY_reg_39_inst : DFFPOSX1 port map( D => n1689, CLK => CLK, Q => 
                           PLAINKEY_39_port);
   PLAINKEY_reg_38_inst : DFFPOSX1 port map( D => n1690, CLK => CLK, Q => 
                           PLAINKEY_38_port);
   PLAINKEY_reg_37_inst : DFFPOSX1 port map( D => n1691, CLK => CLK, Q => 
                           PLAINKEY_37_port);
   PLAINKEY_reg_36_inst : DFFPOSX1 port map( D => n1692, CLK => CLK, Q => 
                           PLAINKEY_36_port);
   PLAINKEY_reg_35_inst : DFFPOSX1 port map( D => n1693, CLK => CLK, Q => 
                           PLAINKEY_35_port);
   PLAINKEY_reg_34_inst : DFFPOSX1 port map( D => n1694, CLK => CLK, Q => 
                           PLAINKEY_34_port);
   PLAINKEY_reg_33_inst : DFFPOSX1 port map( D => n1695, CLK => CLK, Q => 
                           PLAINKEY_33_port);
   PLAINKEY_reg_32_inst : DFFPOSX1 port map( D => n1696, CLK => CLK, Q => 
                           PLAINKEY_32_port);
   PLAINKEY_reg_31_inst : DFFPOSX1 port map( D => n1697, CLK => CLK, Q => 
                           PLAINKEY_31_port);
   PLAINKEY_reg_30_inst : DFFPOSX1 port map( D => n1698, CLK => CLK, Q => 
                           PLAINKEY_30_port);
   PLAINKEY_reg_29_inst : DFFPOSX1 port map( D => n1699, CLK => CLK, Q => 
                           PLAINKEY_29_port);
   PLAINKEY_reg_28_inst : DFFPOSX1 port map( D => n1700, CLK => CLK, Q => 
                           PLAINKEY_28_port);
   PLAINKEY_reg_27_inst : DFFPOSX1 port map( D => n1701, CLK => CLK, Q => 
                           PLAINKEY_27_port);
   PLAINKEY_reg_26_inst : DFFPOSX1 port map( D => n1702, CLK => CLK, Q => 
                           PLAINKEY_26_port);
   PLAINKEY_reg_25_inst : DFFPOSX1 port map( D => n1703, CLK => CLK, Q => 
                           PLAINKEY_25_port);
   PLAINKEY_reg_24_inst : DFFPOSX1 port map( D => n1704, CLK => CLK, Q => 
                           PLAINKEY_24_port);
   PLAINKEY_reg_23_inst : DFFPOSX1 port map( D => n1705, CLK => CLK, Q => 
                           PLAINKEY_23_port);
   PLAINKEY_reg_22_inst : DFFPOSX1 port map( D => n1706, CLK => CLK, Q => 
                           PLAINKEY_22_port);
   PLAINKEY_reg_21_inst : DFFPOSX1 port map( D => n1707, CLK => CLK, Q => 
                           PLAINKEY_21_port);
   PLAINKEY_reg_20_inst : DFFPOSX1 port map( D => n1708, CLK => CLK, Q => 
                           PLAINKEY_20_port);
   PLAINKEY_reg_19_inst : DFFPOSX1 port map( D => n1709, CLK => CLK, Q => 
                           PLAINKEY_19_port);
   PLAINKEY_reg_18_inst : DFFPOSX1 port map( D => n1710, CLK => CLK, Q => 
                           PLAINKEY_18_port);
   PLAINKEY_reg_17_inst : DFFPOSX1 port map( D => n1711, CLK => CLK, Q => 
                           PLAINKEY_17_port);
   PLAINKEY_reg_16_inst : DFFPOSX1 port map( D => n1712, CLK => CLK, Q => 
                           PLAINKEY_16_port);
   PLAINKEY_reg_15_inst : DFFPOSX1 port map( D => n1713, CLK => CLK, Q => 
                           PLAINKEY_15_port);
   PLAINKEY_reg_14_inst : DFFPOSX1 port map( D => n1714, CLK => CLK, Q => 
                           PLAINKEY_14_port);
   PLAINKEY_reg_13_inst : DFFPOSX1 port map( D => n1715, CLK => CLK, Q => 
                           PLAINKEY_13_port);
   PLAINKEY_reg_12_inst : DFFPOSX1 port map( D => n1716, CLK => CLK, Q => 
                           PLAINKEY_12_port);
   PLAINKEY_reg_11_inst : DFFPOSX1 port map( D => n1717, CLK => CLK, Q => 
                           PLAINKEY_11_port);
   PLAINKEY_reg_10_inst : DFFPOSX1 port map( D => n1718, CLK => CLK, Q => 
                           PLAINKEY_10_port);
   PLAINKEY_reg_9_inst : DFFPOSX1 port map( D => n1719, CLK => CLK, Q => 
                           PLAINKEY_9_port);
   PLAINKEY_reg_8_inst : DFFPOSX1 port map( D => n1720, CLK => CLK, Q => 
                           PLAINKEY_8_port);
   PLAINKEY_reg_7_inst : DFFPOSX1 port map( D => n1721, CLK => CLK, Q => 
                           PLAINKEY_7_port);
   PLAINKEY_reg_6_inst : DFFPOSX1 port map( D => n1722, CLK => CLK, Q => 
                           PLAINKEY_6_port);
   PLAINKEY_reg_5_inst : DFFPOSX1 port map( D => n1723, CLK => CLK, Q => 
                           PLAINKEY_5_port);
   PLAINKEY_reg_4_inst : DFFPOSX1 port map( D => n1724, CLK => CLK, Q => 
                           PLAINKEY_4_port);
   PLAINKEY_reg_3_inst : DFFPOSX1 port map( D => n1725, CLK => CLK, Q => 
                           PLAINKEY_3_port);
   PLAINKEY_reg_2_inst : DFFPOSX1 port map( D => n1726, CLK => CLK, Q => 
                           PLAINKEY_2_port);
   PLAINKEY_reg_1_inst : DFFPOSX1 port map( D => n1727, CLK => CLK, Q => 
                           PLAINKEY_1_port);
   PLAINKEY_reg_0_inst : DFFPOSX1 port map( D => n1728, CLK => CLK, Q => 
                           PLAINKEY_0_port);
   U9 : NAND3X1 port map( A => parityAccumulator_7_port, B => 
                           parityAccumulator_6_port, C => n2035, Y => n2036);
   U10 : NOR2X1 port map( A => n1486, B => n1487, Y => n2035);
   U11 : NAND3X1 port map( A => parityAccumulator_3_port, B => 
                           parityAccumulator_2_port, C => n2034, Y => n2037);
   U12 : NOR2X1 port map( A => n1482, B => n1483, Y => n2034);
   U13 : OAI21X1 port map( A => n223, B => n1569, C => n2033, Y => n1728);
   U14 : NAND2X1 port map( A => PLAINKEY_0_port, B => n227, Y => n2033);
   U15 : OAI21X1 port map( A => n223, B => n1568, C => n2032, Y => n1727);
   U16 : NAND2X1 port map( A => PLAINKEY_1_port, B => RST, Y => n2032);
   U17 : OAI21X1 port map( A => n223, B => n1567, C => n2031, Y => n1726);
   U18 : NAND2X1 port map( A => PLAINKEY_2_port, B => RST, Y => n2031);
   U19 : OAI21X1 port map( A => n223, B => n1566, C => n2030, Y => n1725);
   U20 : NAND2X1 port map( A => PLAINKEY_3_port, B => RST, Y => n2030);
   U21 : OAI21X1 port map( A => n223, B => n1565, C => n2029, Y => n1724);
   U22 : NAND2X1 port map( A => PLAINKEY_4_port, B => n227, Y => n2029);
   U24 : OAI21X1 port map( A => n223, B => n1564, C => n2028, Y => n1723);
   U25 : NAND2X1 port map( A => PLAINKEY_5_port, B => n228, Y => n2028);
   U27 : OAI21X1 port map( A => n223, B => n1563, C => n2027, Y => n1722);
   U28 : NAND2X1 port map( A => PLAINKEY_6_port, B => n229, Y => n2027);
   U30 : OAI21X1 port map( A => n223, B => n1562, C => n2026, Y => n1721);
   U31 : NAND2X1 port map( A => PLAINKEY_7_port, B => RST, Y => n2026);
   U33 : OAI21X1 port map( A => n223, B => n1561, C => n2025, Y => n1720);
   U34 : NAND2X1 port map( A => PLAINKEY_8_port, B => n227, Y => n2025);
   U36 : OAI21X1 port map( A => n224, B => n1560, C => n2024, Y => n1719);
   U37 : NAND2X1 port map( A => PLAINKEY_9_port, B => n228, Y => n2024);
   U39 : OAI21X1 port map( A => n224, B => n1559, C => n2023, Y => n1718);
   U40 : NAND2X1 port map( A => PLAINKEY_10_port, B => n229, Y => n2023);
   U42 : OAI21X1 port map( A => n224, B => n1558, C => n2022, Y => n1717);
   U43 : NAND2X1 port map( A => PLAINKEY_11_port, B => n229, Y => n2022);
   U45 : OAI21X1 port map( A => n224, B => n1557, C => n2021, Y => n1716);
   U46 : NAND2X1 port map( A => PLAINKEY_12_port, B => n229, Y => n2021);
   U48 : OAI21X1 port map( A => n224, B => n1556, C => n2020, Y => n1715);
   U49 : NAND2X1 port map( A => PLAINKEY_13_port, B => n229, Y => n2020);
   U51 : OAI21X1 port map( A => n224, B => n1555, C => n2019, Y => n1714);
   U52 : NAND2X1 port map( A => PLAINKEY_14_port, B => n229, Y => n2019);
   U54 : OAI21X1 port map( A => n224, B => n1554, C => n2018, Y => n1713);
   U55 : NAND2X1 port map( A => PLAINKEY_15_port, B => n229, Y => n2018);
   U57 : OAI21X1 port map( A => n225, B => n1553, C => n2017, Y => n1712);
   U58 : NAND2X1 port map( A => PLAINKEY_16_port, B => n229, Y => n2017);
   U60 : OAI21X1 port map( A => n225, B => n1552, C => n2016, Y => n1711);
   U61 : NAND2X1 port map( A => PLAINKEY_17_port, B => n229, Y => n2016);
   U63 : OAI21X1 port map( A => n225, B => n1551, C => n2015, Y => n1710);
   U64 : NAND2X1 port map( A => PLAINKEY_18_port, B => n229, Y => n2015);
   U66 : OAI21X1 port map( A => n225, B => n1550, C => n2014, Y => n1709);
   U67 : NAND2X1 port map( A => PLAINKEY_19_port, B => n229, Y => n2014);
   U69 : OAI21X1 port map( A => n225, B => n1549, C => n2013, Y => n1708);
   U70 : NAND2X1 port map( A => PLAINKEY_20_port, B => n229, Y => n2013);
   U72 : OAI21X1 port map( A => n225, B => n1548, C => n2012, Y => n1707);
   U73 : NAND2X1 port map( A => PLAINKEY_21_port, B => n229, Y => n2012);
   U75 : OAI21X1 port map( A => n225, B => n1547, C => n2011, Y => n1706);
   U76 : NAND2X1 port map( A => PLAINKEY_22_port, B => n229, Y => n2011);
   U78 : OAI21X1 port map( A => n226, B => n1546, C => n2010, Y => n1705);
   U79 : NAND2X1 port map( A => PLAINKEY_23_port, B => n229, Y => n2010);
   U81 : OAI21X1 port map( A => n225, B => n1545, C => n2009, Y => n1704);
   U82 : NAND2X1 port map( A => PLAINKEY_24_port, B => n229, Y => n2009);
   U84 : OAI21X1 port map( A => n224, B => n1544, C => n2008, Y => n1703);
   U85 : NAND2X1 port map( A => PLAINKEY_25_port, B => n229, Y => n2008);
   U87 : OAI21X1 port map( A => n226, B => n1543, C => n2007, Y => n1702);
   U88 : NAND2X1 port map( A => PLAINKEY_26_port, B => n229, Y => n2007);
   U90 : OAI21X1 port map( A => n226, B => n1542, C => n2006, Y => n1701);
   U91 : NAND2X1 port map( A => PLAINKEY_27_port, B => n229, Y => n2006);
   U93 : OAI21X1 port map( A => n225, B => n1541, C => n2005, Y => n1700);
   U94 : NAND2X1 port map( A => PLAINKEY_28_port, B => n229, Y => n2005);
   U96 : OAI21X1 port map( A => n226, B => n1540, C => n2004, Y => n1699);
   U97 : NAND2X1 port map( A => PLAINKEY_29_port, B => n228, Y => n2004);
   U99 : OAI21X1 port map( A => n226, B => n1539, C => n2003, Y => n1698);
   U100 : NAND2X1 port map( A => PLAINKEY_30_port, B => n228, Y => n2003);
   U102 : OAI21X1 port map( A => n225, B => n1538, C => n2002, Y => n1697);
   U103 : NAND2X1 port map( A => PLAINKEY_31_port, B => n228, Y => n2002);
   U105 : OAI21X1 port map( A => RST, B => n1537, C => n2001, Y => n1696);
   U106 : NAND2X1 port map( A => PLAINKEY_32_port, B => n228, Y => n2001);
   U108 : OAI21X1 port map( A => n226, B => n1536, C => n2000, Y => n1695);
   U109 : NAND2X1 port map( A => PLAINKEY_33_port, B => n228, Y => n2000);
   U111 : OAI21X1 port map( A => n229, B => n1535, C => n1999, Y => n1694);
   U112 : NAND2X1 port map( A => PLAINKEY_34_port, B => n228, Y => n1999);
   U114 : OAI21X1 port map( A => n226, B => n1534, C => n1998, Y => n1693);
   U115 : NAND2X1 port map( A => PLAINKEY_35_port, B => n228, Y => n1998);
   U117 : OAI21X1 port map( A => n226, B => n1533, C => n1997, Y => n1692);
   U118 : NAND2X1 port map( A => PLAINKEY_36_port, B => n228, Y => n1997);
   U120 : OAI21X1 port map( A => n227, B => n1532, C => n1996, Y => n1691);
   U121 : NAND2X1 port map( A => PLAINKEY_37_port, B => n228, Y => n1996);
   U123 : OAI21X1 port map( A => n223, B => n1531, C => n1995, Y => n1690);
   U124 : NAND2X1 port map( A => PLAINKEY_38_port, B => n228, Y => n1995);
   U126 : OAI21X1 port map( A => n226, B => n1530, C => n1994, Y => n1689);
   U127 : NAND2X1 port map( A => PLAINKEY_39_port, B => n228, Y => n1994);
   U129 : OAI21X1 port map( A => n225, B => n1529, C => n1993, Y => n1688);
   U130 : NAND2X1 port map( A => PLAINKEY_40_port, B => n228, Y => n1993);
   U132 : OAI21X1 port map( A => n226, B => n1528, C => n1992, Y => n1687);
   U133 : NAND2X1 port map( A => PLAINKEY_41_port, B => n228, Y => n1992);
   U135 : OAI21X1 port map( A => n226, B => n1527, C => n1991, Y => n1686);
   U136 : NAND2X1 port map( A => PLAINKEY_42_port, B => n228, Y => n1991);
   U138 : OAI21X1 port map( A => RST, B => n1526, C => n1990, Y => n1685);
   U139 : NAND2X1 port map( A => PLAINKEY_43_port, B => n228, Y => n1990);
   U141 : OAI21X1 port map( A => n224, B => n1525, C => n1989, Y => n1684);
   U142 : NAND2X1 port map( A => PLAINKEY_44_port, B => n227, Y => n1989);
   U144 : OAI21X1 port map( A => n224, B => n1524, C => n1988, Y => n1683);
   U145 : NAND2X1 port map( A => PLAINKEY_45_port, B => n227, Y => n1988);
   U147 : OAI21X1 port map( A => n228, B => n1523, C => n1987, Y => n1682);
   U148 : NAND2X1 port map( A => PLAINKEY_46_port, B => n228, Y => n1987);
   U150 : OAI21X1 port map( A => n224, B => n1522, C => n1986, Y => n1681);
   U151 : NAND2X1 port map( A => PLAINKEY_47_port, B => n227, Y => n1986);
   U153 : OAI21X1 port map( A => n226, B => n1521, C => n1985, Y => n1680);
   U154 : NAND2X1 port map( A => PLAINKEY_48_port, B => n227, Y => n1985);
   U156 : OAI21X1 port map( A => n226, B => n1520, C => n1984, Y => n1679);
   U157 : NAND2X1 port map( A => PLAINKEY_49_port, B => n227, Y => n1984);
   U159 : OAI21X1 port map( A => n226, B => n1519, C => n1983, Y => n1678);
   U160 : NAND2X1 port map( A => PLAINKEY_50_port, B => n227, Y => n1983);
   U162 : OAI21X1 port map( A => n225, B => n1518, C => n1982, Y => n1677);
   U163 : NAND2X1 port map( A => PLAINKEY_51_port, B => n227, Y => n1982);
   U165 : OAI21X1 port map( A => n226, B => n1517, C => n1981, Y => n1676);
   U166 : NAND2X1 port map( A => PLAINKEY_52_port, B => n227, Y => n1981);
   U168 : OAI21X1 port map( A => n225, B => n1516, C => n1980, Y => n1675);
   U169 : NAND2X1 port map( A => PLAINKEY_53_port, B => n227, Y => n1980);
   U171 : OAI21X1 port map( A => n225, B => n1515, C => n1979, Y => n1674);
   U172 : NAND2X1 port map( A => PLAINKEY_54_port, B => n227, Y => n1979);
   U174 : OAI21X1 port map( A => n224, B => n1514, C => n1978, Y => n1673);
   U175 : NAND2X1 port map( A => PLAINKEY_55_port, B => n228, Y => n1978);
   U177 : OAI21X1 port map( A => n225, B => n1513, C => n1977, Y => n1672);
   U178 : NAND2X1 port map( A => PLAINKEY_56_port, B => n227, Y => n1977);
   U180 : OAI21X1 port map( A => n224, B => n1512, C => n1976, Y => n1671);
   U181 : NAND2X1 port map( A => PLAINKEY_57_port, B => n227, Y => n1976);
   U183 : OAI21X1 port map( A => n224, B => n1511, C => n1975, Y => n1670);
   U184 : NAND2X1 port map( A => PLAINKEY_58_port, B => n227, Y => n1975);
   U186 : OAI21X1 port map( A => n224, B => n1510, C => n1974, Y => n1669);
   U187 : NAND2X1 port map( A => PLAINKEY_59_port, B => n227, Y => n1974);
   U188 : OAI21X1 port map( A => n223, B => n1509, C => n1973, Y => n1668);
   U189 : NAND2X1 port map( A => PLAINKEY_60_port, B => n227, Y => n1973);
   U191 : OAI21X1 port map( A => n223, B => n1508, C => n1972, Y => n1667);
   U192 : NAND2X1 port map( A => PLAINKEY_61_port, B => n227, Y => n1972);
   U194 : OAI21X1 port map( A => n223, B => n1507, C => n1971, Y => n1666);
   U195 : NAND2X1 port map( A => PLAINKEY_62_port, B => n227, Y => n1971);
   U196 : OAI21X1 port map( A => n223, B => n1506, C => n1970, Y => n1665);
   U197 : NAND2X1 port map( A => PLAINKEY_63_port, B => n228, Y => n1970);
   U202 : OAI21X1 port map( A => n1445, B => n1965, C => n1967, Y => n1968);
   U203 : AOI22X1 port map( A => n1964, B => n1963, C => n1494, D => n1572, Y 
                           => n1965);
   U205 : OAI22X1 port map( A => RCV_DATA(3), B => n1962, C => n1495, D => 
                           n1961, Y => n1964);
   U206 : AOI22X1 port map( A => n1960, B => n1959, C => n1496, D => n1574, Y 
                           => n1961);
   U208 : OAI22X1 port map( A => n1958, B => n1497, C => n221, D => n1957, Y =>
                           n1960);
   U210 : NAND2X1 port map( A => n21, B => n6, Y => n1957);
   U211 : AOI22X1 port map( A => n1956, B => n1575, C => n1503, D => n1506, Y 
                           => n1958);
   U213 : NOR2X1 port map( A => n1955, B => n127, Y => n1956);
   U220 : OAI22X1 port map( A => n1967, B => n1571, C => n1966, D => n1572, Y 
                           => n1953);
   U221 : OAI21X1 port map( A => n1963, B => n1573, C => n1952, Y => n1954);
   U222 : AOI22X1 port map( A => RCV_DATA(2), B => n1495, C => n1492, D => 
                           n1951, Y => n1952);
   U223 : OAI21X1 port map( A => n1959, B => n222, C => n1950, Y => n1951);
   U224 : NAND2X1 port map( A => n1949, B => n1959, Y => n1950);
   U225 : OAI21X1 port map( A => n1955, B => n1948, C => n1947, Y => n1949);
   U226 : OAI21X1 port map( A => n1946, B => n1955, C => 
                           currentPlainKey_62_port, Y => n1947);
   U227 : NAND2X1 port map( A => n20, B => n6, Y => n1959);
   U233 : OAI21X1 port map( A => n1943, B => n1942, C => n1969, Y => n1944);
   U234 : OAI22X1 port map( A => n1967, B => n1572, C => n1963, D => n1574, Y 
                           => n1942);
   U235 : OAI21X1 port map( A => n1941, B => n1945, C => n1940, Y => n1943);
   U236 : AOI22X1 port map( A => n221, B => n1495, C => RCV_DATA(3), D => n1445
                           , Y => n1940);
   U238 : NAND2X1 port map( A => n1939, B => n1962, Y => n1945);
   U239 : NAND2X1 port map( A => n19, B => n6, Y => n1962);
   U240 : AOI22X1 port map( A => n1938, B => n139, C => currentPlainKey_61_port
                           , D => n1502, Y => n1941);
   U242 : NOR2X1 port map( A => n1955, B => n1937, Y => n1938);
   U252 : OAI21X1 port map( A => n1955, B => n1935, C => n1934, Y => n1936);
   U253 : OAI21X1 port map( A => n1933, B => n1955, C => 
                           currentPlainKey_60_port, Y => n1934);
   U264 : OAI21X1 port map( A => n1967, B => n1574, C => n1929, Y => n1930);
   U265 : AOI22X1 port map( A => n1932, B => n1928, C => n221, D => n1445, Y =>
                           n1929);
   U266 : OAI22X1 port map( A => n1927, B => n1510, C => n1575, D => n1501, Y 
                           => n1928);
   U270 : NOR2X1 port map( A => n1955, B => n1926, Y => n1927);
   U271 : NOR2X1 port map( A => n1445, B => n1493, Y => n1932);
   U284 : OAI22X1 port map( A => n1967, B => n222, C => n1493, D => n1924, Y =>
                           n1925);
   U285 : AOI22X1 port map( A => n1923, B => n139, C => currentPlainKey_58_port
                           , D => n1500, Y => n1924);
   U287 : NOR2X1 port map( A => n1955, B => n1922, Y => n1923);
   U300 : AOI22X1 port map( A => n1919, B => n1969, C => n221, D => n1446, Y =>
                           n1920);
   U303 : OAI21X1 port map( A => n1955, B => n1918, C => n1917, Y => n1919);
   U304 : OAI21X1 port map( A => n1916, B => n1955, C => 
                           currentPlainKey_57_port, Y => n1917);
   U314 : OAI21X1 port map( A => n1955, B => n1914, C => n1913, Y => n1915);
   U315 : OAI21X1 port map( A => n1912, B => n1955, C => 
                           currentPlainKey_56_port, Y => n1913);
   U316 : NAND2X1 port map( A => address_3_port, B => n1911, Y => n1955);
   U330 : AOI22X1 port map( A => n1908, B => n1931, C => n1447, D => n221, Y =>
                           n1909);
   U333 : OAI21X1 port map( A => n151, B => n1907, C => n1906, Y => n1908);
   U334 : OAI21X1 port map( A => n127, B => n151, C => currentPlainKey_55_port,
                           Y => n1906);
   U344 : OAI21X1 port map( A => n1948, B => n151, C => n1904, Y => n1905);
   U345 : OAI21X1 port map( A => n1946, B => n151, C => currentPlainKey_54_port
                           , Y => n1904);
   U359 : AOI22X1 port map( A => n1901, B => n1921, C => n1448, D => n221, Y =>
                           n1902);
   U362 : OAI21X1 port map( A => n151, B => n1900, C => n1899, Y => n1901);
   U363 : OAI21X1 port map( A => n1937, B => n151, C => currentPlainKey_53_port
                           , Y => n1899);
   U373 : OAI21X1 port map( A => n1935, B => n151, C => n1897, Y => n1898);
   U374 : OAI21X1 port map( A => n1933, B => n151, C => currentPlainKey_52_port
                           , Y => n1897);
   U388 : AOI22X1 port map( A => n1894, B => n1910, C => n1449, D => n221, Y =>
                           n1895);
   U391 : OAI21X1 port map( A => n151, B => n1893, C => n1892, Y => n1894);
   U392 : OAI21X1 port map( A => n1926, B => n151, C => currentPlainKey_51_port
                           , Y => n1892);
   U402 : OAI21X1 port map( A => n151, B => n1890, C => n1889, Y => n1891);
   U403 : OAI21X1 port map( A => n1922, B => n151, C => currentPlainKey_50_port
                           , Y => n1889);
   U417 : AOI22X1 port map( A => n1886, B => n1903, C => n1450, D => n221, Y =>
                           n1887);
   U422 : OAI21X1 port map( A => n1918, B => n151, C => n1884, Y => n1886);
   U423 : OAI21X1 port map( A => n1916, B => n151, C => currentPlainKey_49_port
                           , Y => n1884);
   U433 : OAI21X1 port map( A => n1914, B => n151, C => n1882, Y => n1883);
   U434 : OAI21X1 port map( A => n1912, B => n151, C => currentPlainKey_48_port
                           , Y => n1882);
   U449 : AOI22X1 port map( A => n1879, B => n1896, C => n1451, D => n221, Y =>
                           n1880);
   U452 : OAI21X1 port map( A => n1907, B => n150, C => n1878, Y => n1879);
   U453 : OAI21X1 port map( A => n127, B => n150, C => currentPlainKey_47_port,
                           Y => n1878);
   U463 : OAI21X1 port map( A => n1948, B => n150, C => n1876, Y => n1877);
   U464 : OAI21X1 port map( A => n1946, B => n150, C => currentPlainKey_46_port
                           , Y => n1876);
   U478 : AOI22X1 port map( A => n1873, B => n1888, C => n1452, D => n221, Y =>
                           n1874);
   U481 : OAI21X1 port map( A => n1900, B => n150, C => n1872, Y => n1873);
   U482 : OAI21X1 port map( A => n1937, B => n150, C => currentPlainKey_45_port
                           , Y => n1872);
   U492 : OAI21X1 port map( A => n1935, B => n150, C => n1870, Y => n1871);
   U493 : OAI21X1 port map( A => n1933, B => n150, C => currentPlainKey_44_port
                           , Y => n1870);
   U507 : AOI22X1 port map( A => n1867, B => n1881, C => n1453, D => n221, Y =>
                           n1868);
   U510 : OAI21X1 port map( A => n1893, B => n150, C => n1866, Y => n1867);
   U511 : OAI21X1 port map( A => n1926, B => n150, C => currentPlainKey_43_port
                           , Y => n1866);
   U521 : OAI21X1 port map( A => n1890, B => n150, C => n1864, Y => n1865);
   U522 : OAI21X1 port map( A => n1922, B => n150, C => currentPlainKey_42_port
                           , Y => n1864);
   U536 : AOI22X1 port map( A => n1861, B => n1875, C => n1454, D => n221, Y =>
                           n1862);
   U539 : OAI21X1 port map( A => n1918, B => n150, C => n1860, Y => n1861);
   U540 : OAI21X1 port map( A => n1916, B => n150, C => currentPlainKey_41_port
                           , Y => n1860);
   U550 : OAI21X1 port map( A => n1914, B => n150, C => n1858, Y => n1859);
   U551 : OAI21X1 port map( A => n1912, B => n150, C => currentPlainKey_40_port
                           , Y => n1858);
   U566 : AOI22X1 port map( A => n1854, B => n1869, C => n1455, D => n221, Y =>
                           n1855);
   U569 : OAI21X1 port map( A => n1907, B => n149, C => n1853, Y => n1854);
   U570 : OAI21X1 port map( A => n127, B => n149, C => currentPlainKey_39_port,
                           Y => n1853);
   U580 : OAI21X1 port map( A => n1948, B => n149, C => n1851, Y => n1852);
   U581 : OAI21X1 port map( A => n1946, B => n149, C => currentPlainKey_38_port
                           , Y => n1851);
   U595 : AOI22X1 port map( A => n1848, B => n1863, C => n1456, D => n221, Y =>
                           n1849);
   U598 : OAI21X1 port map( A => n1900, B => n149, C => n1847, Y => n1848);
   U599 : OAI21X1 port map( A => n1937, B => n149, C => currentPlainKey_37_port
                           , Y => n1847);
   U609 : OAI21X1 port map( A => n1935, B => n149, C => n1845, Y => n1846);
   U610 : OAI21X1 port map( A => n1933, B => n149, C => currentPlainKey_36_port
                           , Y => n1845);
   U624 : AOI22X1 port map( A => n1842, B => n1856, C => n1457, D => n221, Y =>
                           n1843);
   U627 : OAI21X1 port map( A => n1893, B => n149, C => n1841, Y => n1842);
   U628 : OAI21X1 port map( A => n1926, B => n149, C => currentPlainKey_35_port
                           , Y => n1841);
   U638 : OAI21X1 port map( A => n1890, B => n149, C => n1839, Y => n1840);
   U639 : OAI21X1 port map( A => n1922, B => n149, C => currentPlainKey_34_port
                           , Y => n1839);
   U653 : AOI22X1 port map( A => n1836, B => n1850, C => n1458, D => n221, Y =>
                           n1837);
   U658 : OAI21X1 port map( A => n1918, B => n149, C => n1835, Y => n1836);
   U659 : OAI21X1 port map( A => n1916, B => n149, C => currentPlainKey_33_port
                           , Y => n1835);
   U669 : OAI21X1 port map( A => n1914, B => n149, C => n1833, Y => n1834);
   U670 : OAI21X1 port map( A => n1912, B => n149, C => currentPlainKey_32_port
                           , Y => n1833);
   U672 : NOR2X1 port map( A => n1504, B => address_4_port, Y => n1857);
   U686 : AOI22X1 port map( A => n1830, B => n1844, C => n1459, D => n221, Y =>
                           n1831);
   U689 : OAI21X1 port map( A => n1907, B => n147, C => n1829, Y => n1830);
   U690 : OAI21X1 port map( A => n127, B => n147, C => currentPlainKey_31_port,
                           Y => n1829);
   U700 : OAI21X1 port map( A => n1948, B => n147, C => n1827, Y => n1828);
   U701 : OAI21X1 port map( A => n1946, B => n147, C => currentPlainKey_30_port
                           , Y => n1827);
   U715 : AOI22X1 port map( A => n1824, B => n1838, C => n1460, D => n221, Y =>
                           n1825);
   U718 : OAI21X1 port map( A => n1900, B => n147, C => n1823, Y => n1824);
   U719 : OAI21X1 port map( A => n1937, B => n147, C => currentPlainKey_29_port
                           , Y => n1823);
   U729 : OAI21X1 port map( A => n1935, B => n147, C => n1821, Y => n1822);
   U730 : OAI21X1 port map( A => n1933, B => n147, C => currentPlainKey_28_port
                           , Y => n1821);
   U744 : AOI22X1 port map( A => n1818, B => n1832, C => n1461, D => n221, Y =>
                           n1819);
   U747 : OAI21X1 port map( A => n1893, B => n147, C => n1817, Y => n1818);
   U748 : OAI21X1 port map( A => n1926, B => n147, C => currentPlainKey_27_port
                           , Y => n1817);
   U758 : OAI21X1 port map( A => n1890, B => n147, C => n1815, Y => n1816);
   U759 : OAI21X1 port map( A => n1922, B => n147, C => currentPlainKey_26_port
                           , Y => n1815);
   U773 : AOI22X1 port map( A => n1812, B => n1826, C => n1462, D => n221, Y =>
                           n1813);
   U776 : OAI21X1 port map( A => n1918, B => n147, C => n1811, Y => n1812);
   U777 : OAI21X1 port map( A => n1916, B => n147, C => currentPlainKey_25_port
                           , Y => n1811);
   U787 : OAI21X1 port map( A => n1914, B => n147, C => n1809, Y => n1810);
   U788 : OAI21X1 port map( A => n1912, B => n147, C => currentPlainKey_24_port
                           , Y => n1809);
   U803 : AOI22X1 port map( A => n1805, B => n1820, C => n1463, D => n221, Y =>
                           n1806);
   U806 : OAI21X1 port map( A => n1907, B => n145, C => n1804, Y => n1805);
   U807 : OAI21X1 port map( A => n127, B => n145, C => currentPlainKey_23_port,
                           Y => n1804);
   U817 : OAI21X1 port map( A => n1948, B => n145, C => n1802, Y => n1803);
   U818 : OAI21X1 port map( A => n1946, B => n145, C => currentPlainKey_22_port
                           , Y => n1802);
   U832 : AOI22X1 port map( A => n1799_port, B => n1814, C => n1464, D => n221,
                           Y => n1800);
   U835 : OAI21X1 port map( A => n1900, B => n145, C => n1798_port, Y => 
                           n1799_port);
   U836 : OAI21X1 port map( A => n1937, B => n145, C => currentPlainKey_21_port
                           , Y => n1798_port);
   U846 : OAI21X1 port map( A => n1935, B => n145, C => n1796_port, Y => 
                           n1797_port);
   U847 : OAI21X1 port map( A => n1933, B => n145, C => currentPlainKey_20_port
                           , Y => n1796_port);
   U861 : AOI22X1 port map( A => n1793_port, B => n1807, C => n1465, D => n221,
                           Y => n1794_port);
   U864 : OAI21X1 port map( A => n1893, B => n145, C => n1792_port, Y => 
                           n1793_port);
   U865 : OAI21X1 port map( A => n1926, B => n145, C => currentPlainKey_19_port
                           , Y => n1792_port);
   U875 : OAI21X1 port map( A => n1890, B => n145, C => n1790, Y => n1791);
   U876 : OAI21X1 port map( A => n1922, B => n145, C => currentPlainKey_18_port
                           , Y => n1790);
   U890 : AOI22X1 port map( A => n1787, B => n1801, C => n1466, D => n221, Y =>
                           n1788);
   U895 : OAI21X1 port map( A => n1918, B => n145, C => n1786, Y => n1787);
   U896 : OAI21X1 port map( A => n1916, B => n145, C => currentPlainKey_17_port
                           , Y => n1786);
   U906 : OAI21X1 port map( A => n1914, B => n145, C => n1784, Y => n1785);
   U907 : OAI21X1 port map( A => n1912, B => n145, C => currentPlainKey_16_port
                           , Y => n1784);
   U909 : NOR2X1 port map( A => n1505, B => address_5_port, Y => n1808);
   U923 : AOI22X1 port map( A => n1781, B => n1795_port, C => n1467, D => n221,
                           Y => n1782);
   U926 : OAI21X1 port map( A => n1907, B => n143, C => n1780, Y => n1781);
   U927 : OAI21X1 port map( A => n127, B => n143, C => currentPlainKey_15_port,
                           Y => n1780);
   U937 : OAI21X1 port map( A => n1948, B => n143, C => n1778, Y => n1779);
   U938 : OAI21X1 port map( A => n1946, B => n143, C => currentPlainKey_14_port
                           , Y => n1778);
   U952 : AOI22X1 port map( A => n1775, B => n1789, C => n1468, D => n221, Y =>
                           n1776);
   U955 : OAI21X1 port map( A => n1900, B => n143, C => n1774, Y => n1775);
   U956 : OAI21X1 port map( A => n1937, B => n143, C => currentPlainKey_13_port
                           , Y => n1774);
   U966 : OAI21X1 port map( A => n1935, B => n143, C => n1772, Y => n1773);
   U967 : OAI21X1 port map( A => n1933, B => n143, C => currentPlainKey_12_port
                           , Y => n1772);
   U981 : AOI22X1 port map( A => n1769, B => n1783, C => n1469, D => n221, Y =>
                           n1770);
   U984 : OAI21X1 port map( A => n1893, B => n143, C => n1768, Y => n1769);
   U985 : OAI21X1 port map( A => n1926, B => n143, C => currentPlainKey_11_port
                           , Y => n1768);
   U995 : OAI21X1 port map( A => n1890, B => n143, C => n1766, Y => n1767);
   U996 : OAI21X1 port map( A => n1922, B => n143, C => currentPlainKey_10_port
                           , Y => n1766);
   U1010 : AOI22X1 port map( A => n1763, B => n1777, C => n1470, D => n221, Y 
                           => n1764);
   U1014 : OAI21X1 port map( A => n1918, B => n143, C => n1762, Y => n1763);
   U1015 : OAI21X1 port map( A => n1916, B => n143, C => currentPlainKey_9_port
                           , Y => n1762);
   U1025 : OAI21X1 port map( A => n1914, B => n143, C => n1760, Y => n1761);
   U1026 : OAI21X1 port map( A => n1912, B => n143, C => currentPlainKey_8_port
                           , Y => n1760);
   U1041 : AOI22X1 port map( A => n1757, B => n1771, C => n1471, D => n221, Y 
                           => n1758);
   U1044 : OAI21X1 port map( A => n1907, B => n141, C => n1756, Y => n1757);
   U1045 : OAI21X1 port map( A => n127, B => n141, C => currentPlainKey_7_port,
                           Y => n1756);
   U1046 : NAND2X1 port map( A => n139, B => n7, Y => n1907);
   U1057 : OAI21X1 port map( A => n1948, B => n141, C => n1753, Y => n1754);
   U1058 : OAI21X1 port map( A => n1946, B => n141, C => currentPlainKey_6_port
                           , Y => n1753);
   U1059 : NAND2X1 port map( A => n139, B => n125, Y => n1948);
   U1074 : AOI22X1 port map( A => n1751, B => n1765, C => n1472, D => n221, Y 
                           => n1752);
   U1077 : OAI21X1 port map( A => n1900, B => n141, C => n1750, Y => n1751);
   U1078 : OAI21X1 port map( A => n1937, B => n141, C => currentPlainKey_5_port
                           , Y => n1750);
   U1079 : NAND2X1 port map( A => n139, B => n1474, Y => n1900);
   U1090 : OAI21X1 port map( A => n1935, B => n141, C => n1747, Y => n1748);
   U1091 : OAI21X1 port map( A => n1933, B => n141, C => currentPlainKey_4_port
                           , Y => n1747);
   U1092 : NAND2X1 port map( A => n139, B => n129, Y => n1935);
   U1111 : OAI21X1 port map( A => n1893, B => n141, C => n1745, Y => n1746);
   U1112 : OAI21X1 port map( A => n1926, B => n141, C => currentPlainKey_3_port
                           , Y => n1745);
   U1113 : NAND2X1 port map( A => n139, B => n1477, Y => n1893);
   U1126 : OAI21X1 port map( A => n1890, B => n141, C => n1743, Y => n1744);
   U1127 : OAI21X1 port map( A => n1922, B => n141, C => currentPlainKey_2_port
                           , Y => n1743);
   U1128 : NAND2X1 port map( A => n139, B => n131, Y => n1890);
   U1154 : NOR2X1 port map( A => address_6_port, B => address_7_port, Y => 
                           n1885);
   U1155 : OAI21X1 port map( A => n1918, B => n141, C => n1741, Y => n1742);
   U1156 : OAI21X1 port map( A => n1916, B => n141, C => currentPlainKey_1_port
                           , Y => n1741);
   U1157 : NAND2X1 port map( A => n139, B => n119, Y => n1918);
   U1182 : AOI22X1 port map( A => n9, B => n1572, C => n1739, D => n1738, Y => 
                           n1740);
   U1183 : AOI21X1 port map( A => n1737, B => n1749, C => n9, Y => n1738);
   U1184 : OAI21X1 port map( A => n222, B => n1755, C => n1736, Y => n1737);
   U1185 : NAND2X1 port map( A => n16, B => n1735, Y => n1736);
   U1186 : OAI21X1 port map( A => n1914, B => n141, C => n1734, Y => n1735);
   U1187 : OAI21X1 port map( A => n1912, B => n141, C => currentPlainKey_0_port
                           , Y => n1734);
   U1189 : NOR2X1 port map( A => address_4_port, B => address_5_port, Y => 
                           n1759);
   U1190 : NAND2X1 port map( A => n139, B => n1473, Y => n1914);
   U1199 : AOI22X1 port map( A => n1475, B => RCV_DATA(2), C => n1498, D => 
                           RCV_DATA(3), Y => n1739);
   U1220 : NOR2X1 port map( A => n1504, B => n1505, Y => n1911);
   U1273 : OAI21X1 port map( A => n1476, B => n1480, C => n1733, Y => n1584);
   U1274 : NAND3X1 port map( A => keyCount_0_port, B => n1480, C => n1732, Y =>
                           n1733);
   U1305 : NAND2X1 port map( A => n1576, B => n1570, Y => n1730);
   U1314 : NAND3X1 port map( A => keyCount_2_port, B => keyCount_1_port, C => 
                           n1729, Y => n1731);
   U1315 : NOR2X1 port map( A => keyCount_3_port, B => n1479, Y => n1729);
   U254 : AND2X2 port map( A => n1932, B => n1963, Y => n1939);
   r577 : keyreg_0_DW01_add_0 port map( A(7) => parityAccumulator_7_port, A(6) 
                           => parityAccumulator_6_port, A(5) => 
                           parityAccumulator_5_port, A(4) => 
                           parityAccumulator_4_port, A(3) => 
                           parityAccumulator_3_port, A(2) => 
                           parityAccumulator_2_port, A(1) => 
                           parityAccumulator_1_port, A(0) => 
                           parityAccumulator_0_port, B(7) => RCV_DATA(7), B(6) 
                           => RCV_DATA(6), B(5) => RCV_DATA(5), B(4) => 
                           RCV_DATA(4), B(3) => RCV_DATA(3), B(2) => 
                           RCV_DATA(2), B(1) => n221, B(0) => n139, CI => n2038
                           , SUM(7) => N1799, SUM(6) => N1798, SUM(5) => N1797,
                           SUM(4) => N1796, SUM(3) => N1795, SUM(2) => N1794, 
                           SUM(1) => N1793, SUM(0) => N1792, CO => n_1020);
   state_reg_0_inst : DFFSR port map( D => n1580, CLK => CLK, R => n234, S => 
                           n69, Q => state_0_port);
   state_reg_3_inst : DFFSR port map( D => n1579, CLK => CLK, R => n234, S => 
                           n67, Q => state_3_port);
   state_reg_2_inst : DFFSR port map( D => n1581, CLK => CLK, R => n234, S => 
                           n65, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => n1582, CLK => CLK, R => n234, S => 
                           n63, Q => state_1_port);
   parityError_reg : DFFSR port map( D => nextParityError, CLK => CLK, R => 
                           n234, S => n61, Q => parityError);
   PARITY_ERROR_reg : DFFSR port map( D => nextParityError, CLK => CLK, R => 
                           n234, S => n59, Q => PARITY_ERROR);
   U3 : INVX8 port map( A => n154, Y => n153);
   U4 : INVX2 port map( A => n101, Y => n103);
   U5 : BUFX2 port map( A => n1181, Y => n181);
   U7 : BUFX2 port map( A => n75, Y => n188);
   U8 : BUFX2 port map( A => n1364, Y => n203);
   U23 : INVX2 port map( A => n123, Y => n1391);
   U26 : BUFX2 port map( A => n1367, Y => n219);
   U29 : INVX1 port map( A => n139, Y => n1575);
   U32 : AND2X2 port map( A => n79, B => n1478, Y => n1);
   U35 : AND2X2 port map( A => n81, B => n1478, Y => n2);
   U38 : AND2X2 port map( A => n83, B => n1478, Y => n4);
   U41 : AND2X2 port map( A => n6, B => n1478, Y => n5);
   U44 : AND2X2 port map( A => n1911, B => n1885, Y => n6);
   U47 : AND2X2 port map( A => n53, B => address_0_port, Y => n7);
   U50 : INVX2 port map( A => n11, Y => n154);
   U53 : AND2X2 port map( A => n1477, B => address_3_port, Y => n8);
   U56 : AND2X2 port map( A => n266, B => n19, Y => n9);
   U59 : AND2X2 port map( A => n266, B => n8, Y => n10);
   U62 : INVX2 port map( A => n121, Y => n123);
   U65 : INVX2 port map( A => state_3_port, Y => n115);
   U68 : AND2X2 port map( A => n188, B => n1420, Y => n11);
   U71 : AND2X2 port map( A => n1432, B => n103, Y => n14);
   U74 : AND2X2 port map( A => n295, B => n1755, Y => n16);
   U77 : AND2X2 port map( A => n131, B => address_3_port, Y => n17);
   U80 : AND2X2 port map( A => n129, B => address_3_port, Y => n19);
   U83 : AND2X2 port map( A => n1474, B => address_3_port, Y => n20);
   U86 : AND2X2 port map( A => n125, B => address_3_port, Y => n21);
   U89 : AND2X2 port map( A => n7, B => address_3_port, Y => n23);
   U92 : AND2X2 port map( A => n1473, B => address_3_port, Y => n25);
   U95 : AND2X2 port map( A => n313, B => n340, Y => n27);
   U98 : AND2X2 port map( A => n1888, B => n1010, Y => n29);
   U101 : AND2X2 port map( A => n1875, B => n950, Y => n31);
   U104 : AND2X2 port map( A => n1777, B => n455, Y => n33);
   U107 : AND2X2 port map( A => n1789, B => n515, Y => n35);
   U110 : AND2X2 port map( A => n1826, B => n702, Y => n37);
   U113 : AND2X2 port map( A => n1838, B => n762, Y => n39);
   U116 : AND2X2 port map( A => n1765, B => n392, Y => n41);
   U119 : AND2X2 port map( A => n1801, B => n578, Y => n43);
   U122 : AND2X2 port map( A => n1814, B => n639, Y => n45);
   U125 : AND2X2 port map( A => n1850, B => n825, Y => n47);
   U128 : AND2X2 port map( A => n1863, B => n885, Y => n49);
   U131 : AND2X2 port map( A => n1903, B => n1069, Y => n51);
   U134 : AND2X2 port map( A => address_1_port, B => address_2_port, Y => n53);
   U137 : AND2X2 port map( A => n1939, B => n1936, Y => n55);
   U140 : AND2X2 port map( A => n266, B => n17, Y => n57);
   n59 <= '1';
   n61 <= '1';
   n63 <= '1';
   n65 <= '1';
   n67 <= '1';
   n69 <= '1';
   U161 : INVX1 port map( A => RCV_DATA(0), Y => n137);
   U164 : INVX4 port map( A => n133, Y => n1132);
   U167 : INVX1 port map( A => state_1_port, Y => n244);
   U170 : NAND2X1 port map( A => n111, B => n14, Y => n1425);
   U173 : AND2X1 port map( A => n249, B => n1425, Y => n113);
   U176 : INVX2 port map( A => n91, Y => n71);
   U179 : INVX4 port map( A => n166, Y => n156);
   U182 : AND2X1 port map( A => n1098, B => n221, Y => n73);
   U185 : INVX8 port map( A => n222, Y => n221);
   U190 : INVX2 port map( A => n137, Y => n139);
   U193 : INVX2 port map( A => n231, Y => n226);
   U198 : INVX2 port map( A => n231, Y => n225);
   U199 : INVX2 port map( A => n230, Y => n224);
   U200 : INVX2 port map( A => n230, Y => n223);
   U201 : INVX2 port map( A => n232, Y => n227);
   U204 : INVX2 port map( A => n232, Y => n228);
   U207 : INVX2 port map( A => n233, Y => n229);
   U209 : INVX2 port map( A => n188, Y => n187);
   U212 : BUFX2 port map( A => n234, Y => n232);
   U214 : BUFX2 port map( A => n232, Y => n231);
   U215 : BUFX2 port map( A => n233, Y => n230);
   U216 : BUFX2 port map( A => n234, Y => n233);
   U217 : INVX2 port map( A => n73, Y => n135);
   U218 : INVX2 port map( A => n73, Y => n133);
   U219 : INVX2 port map( A => n189, Y => n186);
   U228 : INVX2 port map( A => n189, Y => n185);
   U229 : INVX2 port map( A => RST, Y => n234);
   U230 : BUFX2 port map( A => n1360, Y => n192);
   U231 : BUFX2 port map( A => n1360, Y => n193);
   U232 : BUFX2 port map( A => n1360, Y => n195);
   U237 : BUFX2 port map( A => n1360, Y => n197);
   U241 : BUFX2 port map( A => n1364, Y => n206);
   U243 : INVX2 port map( A => n165, Y => n160);
   U244 : BUFX2 port map( A => n1364, Y => n205);
   U245 : BUFX2 port map( A => n1181, Y => n183);
   U246 : BUFX2 port map( A => n1181, Y => n180);
   U247 : BUFX2 port map( A => n1181, Y => n178);
   U248 : INVX2 port map( A => n165, Y => n161);
   U249 : INVX2 port map( A => n166, Y => n158);
   U250 : AND2X2 port map( A => n264, B => n1414, Y => n75);
   U251 : BUFX2 port map( A => n1181, Y => n184);
   U255 : BUFX2 port map( A => n1364, Y => n207);
   U256 : INVX2 port map( A => n77, Y => n141);
   U257 : INVX2 port map( A => n85, Y => n151);
   U258 : INVX2 port map( A => n87, Y => n145);
   U259 : INVX2 port map( A => n89, Y => n149);
   U260 : INVX2 port map( A => n177, Y => n173);
   U261 : INVX2 port map( A => n177, Y => n172);
   U262 : INVX2 port map( A => n175, Y => n168);
   U263 : INVX2 port map( A => n1158, Y => n165);
   U267 : INVX2 port map( A => n1158, Y => n166);
   U268 : AND2X2 port map( A => n1759, B => n1478, Y => n77);
   U269 : AND2X2 port map( A => n1857, B => n1885, Y => n79);
   U272 : AND2X2 port map( A => n1759, B => n1885, Y => n81);
   U273 : AND2X2 port map( A => n1808, B => n1885, Y => n83);
   U274 : INVX2 port map( A => n1946, Y => n125);
   U275 : AND2X2 port map( A => n1911, B => n1478, Y => n85);
   U276 : AND2X2 port map( A => n1808, B => n1478, Y => n87);
   U277 : AND2X2 port map( A => n1857, B => n1478, Y => n89);
   U278 : INVX2 port map( A => n93, Y => n143);
   U279 : INVX2 port map( A => n95, Y => n147);
   U280 : INVX2 port map( A => n97, Y => n150);
   U281 : INVX2 port map( A => RCV_DATA(1), Y => n222);
   U282 : AND2X2 port map( A => n11, B => RCV_DATA(2), Y => n91);
   U283 : INVX2 port map( A => n1916, Y => n119);
   U286 : INVX2 port map( A => n1933, Y => n129);
   U288 : INVX2 port map( A => n1922, Y => n131);
   U289 : INVX2 port map( A => n7, Y => n127);
   U290 : AND2X2 port map( A => n1759, B => address_3_port, Y => n93);
   U291 : AND2X2 port map( A => n1808, B => address_3_port, Y => n95);
   U292 : AND2X2 port map( A => n1857, B => address_3_port, Y => n97);
   U293 : NAND2X1 port map( A => n188, B => n1420, Y => n99);
   U294 : INVX2 port map( A => state_2_port, Y => n101);
   U295 : AND2X2 port map( A => n109, B => n1413, Y => n117);
   U296 : BUFX2 port map( A => state_0_port, Y => n105);
   U297 : INVX1 port map( A => n115, Y => n107);
   U298 : INVX2 port map( A => n1427, Y => n1406);
   U299 : INVX2 port map( A => state_0_port, Y => n1432);
   U301 : NOR2X1 port map( A => state_1_port, B => state_0_port, Y => n109);
   U302 : INVX1 port map( A => n109, Y => n1408);
   U305 : AND2X2 port map( A => state_1_port, B => n115, Y => n111);
   U306 : INVX1 port map( A => n123, Y => n1395);
   U307 : INVX1 port map( A => n123, Y => n1393);
   U308 : INVX1 port map( A => n123, Y => n1399);
   U309 : BUFX2 port map( A => n91, Y => n177);
   U310 : BUFX2 port map( A => n91, Y => n175);
   U311 : INVX1 port map( A => n117, Y => n1424);
   U312 : BUFX2 port map( A => n75, Y => n189);
   U313 : INVX1 port map( A => n1426, Y => n1384);
   U317 : INVX2 port map( A => n1403, Y => n121);
   U318 : INVX1 port map( A => n1361, Y => n1098);
   U319 : BUFX4 port map( A => n1367, Y => n208);
   U320 : BUFX4 port map( A => n1367, Y => n209);
   U321 : BUFX4 port map( A => n1367, Y => n210);
   U322 : BUFX4 port map( A => n1367, Y => n217);
   U323 : NAND2X1 port map( A => address_0_port, B => address_1_port, Y => n240
                           );
   U324 : OR2X2 port map( A => address_2_port, B => n240, Y => n1926);
   U325 : INVX2 port map( A => n1926, Y => n1477);
   U326 : NAND2X1 port map( A => n8, B => n6, Y => n1963);
   U327 : INVX2 port map( A => address_2_port, Y => n262);
   U328 : INVX2 port map( A => address_1_port, Y => n261);
   U329 : NAND3X1 port map( A => address_0_port, B => n262, C => n261, Y => 
                           n1916);
   U331 : NAND2X1 port map( A => n119, B => address_3_port, Y => n269);
   U332 : INVX2 port map( A => n269, Y => n917);
   U335 : NAND2X1 port map( A => n917, B => n6, Y => n1967);
   U336 : INVX2 port map( A => n103, Y => n1413);
   U337 : NAND3X1 port map( A => n111, B => n1432, C => n1413, Y => n1438);
   U338 : NAND3X1 port map( A => n103, B => n105, C => n111, Y => n1411);
   U339 : NAND2X1 port map( A => n1438, B => n1411, Y => CLR_RBUFF_port);
   U340 : NAND3X1 port map( A => n109, B => n103, C => n115, Y => n241);
   U341 : INVX2 port map( A => n241, Y => PROG_ERROR_port);
   U342 : NAND3X1 port map( A => n111, B => n105, C => n1413, Y => n1427);
   U343 : OAI21X1 port map( A => n107, B => n1424, C => n1427, Y => n243);
   U346 : NAND2X1 port map( A => n1425, B => n241, Y => n242);
   U347 : NOR3X1 port map( A => CLR_RBUFF_port, B => n243, C => n242, Y => 
                           n1371);
   U348 : NAND2X1 port map( A => n117, B => n107, Y => n1426);
   U349 : NAND3X1 port map( A => n105, B => n244, C => n115, Y => n245);
   U350 : INVX2 port map( A => n245, Y => n247);
   U351 : NAND2X1 port map( A => n247, B => n103, Y => n1414);
   U352 : INVX2 port map( A => n1414, Y => n1435);
   U353 : NAND2X1 port map( A => n247, B => n1413, Y => n249);
   U354 : INVX2 port map( A => n249, Y => n1383);
   U355 : AOI21X1 port map( A => n1435, B => parityError, C => n1383, Y => n248
                           );
   U356 : NAND3X1 port map( A => n1371, B => n1426, C => n248, Y => KEY_ERROR);
   U357 : NOR2X1 port map( A => PROG_ERROR_port, B => n223, Y => n255);
   U358 : NAND2X1 port map( A => n249, B => n1425, Y => n1419);
   U360 : NOR2X1 port map( A => n1406, B => n1419, Y => n250);
   U361 : NAND3X1 port map( A => n255, B => n1426, C => n250, Y => n1403);
   U364 : NAND2X1 port map( A => n1391, B => n1411, Y => n1442);
   U365 : INVX2 port map( A => n1442, Y => n264);
   U366 : INVX2 port map( A => n1438, Y => n1420);
   U367 : NAND2X1 port map( A => n264, B => n1420, Y => n1444);
   U368 : NOR2X1 port map( A => n1490, B => n1444, Y => n1732);
   U369 : NAND2X1 port map( A => keyCount_1_port, B => keyCount_0_port, Y => 
                           n257);
   U370 : NAND2X1 port map( A => n1420, B => n257, Y => n258);
   U371 : NAND2X1 port map( A => n264, B => n258, Y => n1439);
   U372 : INVX2 port map( A => n1439, Y => n1476);
   U375 : INVX2 port map( A => address_0_port, Y => n263);
   U376 : NAND2X1 port map( A => n53, B => n263, Y => n1946);
   U377 : NAND3X1 port map( A => address_6_port, B => address_7_port, C => 
                           n1911, Y => n268);
   U378 : INVX2 port map( A => n268, Y => n266);
   U379 : NAND2X1 port map( A => n266, B => n21, Y => n295);
   U380 : INVX2 port map( A => n295, Y => n1475);
   U381 : NAND2X1 port map( A => address_0_port, B => address_2_port, Y => n259
                           );
   U382 : OR2X2 port map( A => address_1_port, B => n259, Y => n1937);
   U383 : INVX2 port map( A => n1937, Y => n1474);
   U384 : NAND2X1 port map( A => n266, B => n20, Y => n1749);
   U385 : INVX2 port map( A => n1749, Y => n1498);
   U386 : NOR2X1 port map( A => address_2_port, B => address_0_port, Y => n260)
                           ;
   U387 : NAND2X1 port map( A => n260, B => n261, Y => n1912);
   U389 : INVX2 port map( A => n1912, Y => n1473);
   U390 : INVX2 port map( A => address_3_port, Y => n1478);
   U393 : NAND2X1 port map( A => n266, B => n23, Y => n1755);
   U394 : NAND3X1 port map( A => address_2_port, B => n263, C => n261, Y => 
                           n1933);
   U395 : INVX2 port map( A => RCV_DATA(4), Y => n1572);
   U396 : NAND3X1 port map( A => address_1_port, B => n263, C => n262, Y => 
                           n1922);
   U397 : NAND2X1 port map( A => n2, B => n129, Y => n1765);
   U398 : INVX2 port map( A => n1765, Y => n1472);
   U399 : NAND2X1 port map( A => n2, B => n125, Y => n1771);
   U400 : INVX2 port map( A => n1771, Y => n1471);
   U401 : NAND2X1 port map( A => n81, B => n25, Y => n1777);
   U404 : INVX2 port map( A => n1777, Y => n1470);
   U405 : NAND2X1 port map( A => n81, B => n17, Y => n1783);
   U406 : INVX2 port map( A => n1783, Y => n1469);
   U407 : NAND2X1 port map( A => n81, B => n19, Y => n1789);
   U408 : INVX2 port map( A => n1789, Y => n1468);
   U409 : NAND2X1 port map( A => n81, B => n21, Y => n1795_port);
   U410 : INVX2 port map( A => n1795_port, Y => n1467);
   U411 : NAND2X1 port map( A => n4, B => n1473, Y => n1801);
   U412 : INVX2 port map( A => n1801, Y => n1466);
   U413 : NAND2X1 port map( A => n4, B => n131, Y => n1807);
   U414 : INVX2 port map( A => n1807, Y => n1465);
   U415 : NAND2X1 port map( A => n4, B => n129, Y => n1814);
   U416 : INVX2 port map( A => n1814, Y => n1464);
   U418 : NAND2X1 port map( A => n4, B => n125, Y => n1820);
   U419 : INVX2 port map( A => n1820, Y => n1463);
   U420 : NAND2X1 port map( A => n83, B => n25, Y => n1826);
   U421 : INVX2 port map( A => n1826, Y => n1462);
   U424 : NAND2X1 port map( A => n83, B => n17, Y => n1832);
   U425 : INVX2 port map( A => n1832, Y => n1461);
   U426 : NAND2X1 port map( A => n83, B => n19, Y => n1838);
   U427 : INVX2 port map( A => n1838, Y => n1460);
   U428 : NAND2X1 port map( A => n83, B => n21, Y => n1844);
   U429 : INVX2 port map( A => n1844, Y => n1459);
   U430 : NAND2X1 port map( A => n1, B => n1473, Y => n1850);
   U431 : INVX2 port map( A => n1850, Y => n1458);
   U432 : NAND2X1 port map( A => n1, B => n131, Y => n1856);
   U435 : INVX2 port map( A => n1856, Y => n1457);
   U436 : NAND2X1 port map( A => n1, B => n129, Y => n1863);
   U437 : INVX2 port map( A => n1863, Y => n1456);
   U438 : NAND2X1 port map( A => n1, B => n125, Y => n1869);
   U439 : INVX2 port map( A => n1869, Y => n1455);
   U440 : NAND2X1 port map( A => n79, B => n25, Y => n1875);
   U441 : INVX2 port map( A => n1875, Y => n1454);
   U442 : NAND2X1 port map( A => n79, B => n17, Y => n1881);
   U443 : INVX2 port map( A => n1881, Y => n1453);
   U444 : NAND2X1 port map( A => n19, B => n79, Y => n1888);
   U445 : INVX2 port map( A => n1888, Y => n1452);
   U446 : NAND2X1 port map( A => n21, B => n79, Y => n1896);
   U447 : INVX2 port map( A => n1896, Y => n1451);
   U448 : NAND2X1 port map( A => n5, B => n1473, Y => n1903);
   U450 : INVX2 port map( A => n1903, Y => n1450);
   U451 : NAND2X1 port map( A => n5, B => n131, Y => n1910);
   U454 : INVX2 port map( A => n1910, Y => n1449);
   U455 : NAND2X1 port map( A => n5, B => n129, Y => n1921);
   U456 : INVX2 port map( A => n1921, Y => n1448);
   U457 : NAND2X1 port map( A => n5, B => n125, Y => n1931);
   U458 : INVX2 port map( A => n1931, Y => n1447);
   U459 : NAND2X1 port map( A => n25, B => n6, Y => n1969);
   U460 : INVX2 port map( A => n1969, Y => n1446);
   U461 : NAND2X1 port map( A => n6, B => n17, Y => n1966);
   U462 : INVX2 port map( A => n1966, Y => n1445);
   U465 : INVX2 port map( A => RCV_DATA(2), Y => n1574);
   U466 : INVX2 port map( A => RCV_DATA(3), Y => n1573);
   U467 : INVX2 port map( A => RCV_DATA(5), Y => n1571);
   U468 : INVX2 port map( A => currentPlainKey_3_port, Y => n1566);
   U469 : INVX2 port map( A => currentPlainKey_2_port, Y => n1567);
   U470 : INVX2 port map( A => currentPlainKey_1_port, Y => n1568);
   U471 : NAND2X1 port map( A => n187, B => currentPlainKey_0_port, Y => n277);
   U472 : NAND2X1 port map( A => n188, B => n1420, Y => n1361);
   U473 : NAND2X1 port map( A => n11, B => RCV_DATA(5), Y => n1171);
   U474 : OAI21X1 port map( A => n10, B => n99, C => n1171, Y => n265);
   U475 : OAI21X1 port map( A => n1740, B => n10, C => n265, Y => n267);
   U476 : NAND2X1 port map( A => RCV_DATA(6), B => n11, Y => n320);
   U477 : MUX2X1 port map( B => n267, A => n320, S => n57, Y => n271);
   U479 : NAND2X1 port map( A => RCV_DATA(7), B => n153, Y => n1267);
   U480 : INVX2 port map( A => n1267, Y => n1367);
   U483 : NOR2X1 port map( A => n269, B => n268, Y => n270);
   U484 : MUX2X1 port map( B => n271, A => n210, S => n270, Y => n275);
   U485 : NAND2X1 port map( A => n277, B => n275, Y => n1601);
   U486 : NAND2X1 port map( A => n185, B => currentPlainKey_1_port, Y => n291);
   U487 : NAND2X1 port map( A => n1098, B => RCV_DATA(3), Y => n1158);
   U488 : INVX2 port map( A => n1742, Y => n278);
   U489 : NAND2X1 port map( A => n2, B => n1473, Y => n313);
   U490 : INVX2 port map( A => n313, Y => n376);
   U491 : MUX2X1 port map( B => n278, A => n222, S => n376, Y => n280);
   U494 : NOR2X1 port map( A => n1574, B => n1755, Y => n279);
   U495 : AOI21X1 port map( A => n16, B => n280, C => n279, Y => n281);
   U496 : NOR2X1 port map( A => n281, B => n1361, Y => n282);
   U497 : AOI21X1 port map( A => n1475, B => n165, C => n282, Y => n284);
   U498 : NAND2X1 port map( A => n11, B => RCV_DATA(4), Y => n1169);
   U499 : MUX2X1 port map( B => n284, A => n1169, S => n1498, Y => n285);
   U500 : INVX2 port map( A => n1171, Y => n1364);
   U501 : MUX2X1 port map( B => n285, A => n203, S => n9, Y => n286);
   U502 : MUX2X1 port map( B => n286, A => n320, S => n10, Y => n287);
   U503 : MUX2X1 port map( B => n287, A => n219, S => n57, Y => n289);
   U504 : NAND2X1 port map( A => n291, B => n289, Y => n1602);
   U505 : NAND2X1 port map( A => n185, B => currentPlainKey_2_port, Y => n305);
   U506 : NOR2X1 port map( A => n1169, B => n295, Y => n301);
   U508 : NAND2X1 port map( A => n2, B => n119, Y => n340);
   U509 : NAND2X1 port map( A => n27, B => n1098, Y => n331);
   U512 : INVX2 port map( A => n1744, Y => n296);
   U513 : OAI22X1 port map( A => n133, B => n340, C => n331, D => n296, Y => 
                           n298);
   U514 : OAI22X1 port map( A => n1755, B => n156, C => n71, D => n313, Y => 
                           n297);
   U515 : AOI21X1 port map( A => n16, B => n298, C => n297, Y => n299);
   U516 : MUX2X1 port map( B => n299, A => n1171, S => n1498, Y => n300);
   U517 : NOR2X1 port map( A => n301, B => n300, Y => n302);
   U518 : MUX2X1 port map( B => n302, A => n320, S => n9, Y => n303);
   U519 : MUX2X1 port map( B => n303, A => n219, S => n10, Y => n304);
   U520 : NAND2X1 port map( A => n305, B => n304, Y => n1603);
   U523 : NAND2X1 port map( A => n186, B => currentPlainKey_3_port, Y => n327);
   U524 : NAND2X1 port map( A => n1475, B => n203, Y => n319);
   U525 : INVX2 port map( A => n331, Y => n311);
   U526 : NAND2X1 port map( A => n1746, B => n311, Y => n312);
   U527 : NAND2X1 port map( A => n2, B => n131, Y => n343);
   U528 : INVX2 port map( A => n343, Y => n422);
   U529 : MUX2X1 port map( B => n312, A => n135, S => n422, Y => n315);
   U530 : OAI22X1 port map( A => n156, B => n313, C => n71, D => n340, Y => 
                           n314);
   U531 : OAI21X1 port map( A => n315, B => n314, C => n16, Y => n317);
   U532 : INVX2 port map( A => n1169, Y => n1181);
   U533 : INVX2 port map( A => n1755, Y => n370);
   U534 : NAND2X1 port map( A => n181, B => n370, Y => n316);
   U535 : NAND3X1 port map( A => n319, B => n317, C => n316, Y => n321);
   U537 : INVX2 port map( A => n320, Y => n1360);
   U538 : MUX2X1 port map( B => n321, A => n195, S => n1498, Y => n322);
   U541 : MUX2X1 port map( B => n322, A => n1267, S => n9, Y => n324);
   U542 : INVX2 port map( A => n324, Y => n326);
   U543 : NAND2X1 port map( A => n327, B => n326, Y => n1604);
   U544 : AOI22X1 port map( A => currentPlainKey_4_port, B => n186, C => n1475,
                           D => n192, Y => n339);
   U545 : NAND2X1 port map( A => n376, B => n178, Y => n336);
   U546 : OAI22X1 port map( A => n160, B => n340, C => n71, D => n343, Y => 
                           n333);
   U547 : NAND2X1 port map( A => n2, B => n1477, Y => n380);
   U548 : NAND2X1 port map( A => n343, B => n380, Y => n362);
   U549 : INVX2 port map( A => n362, Y => n418);
   U552 : NAND2X1 port map( A => n1748, B => n418, Y => n330);
   U553 : OAI22X1 port map( A => n133, B => n380, C => n331, D => n330, Y => 
                           n332);
   U554 : OAI21X1 port map( A => n333, B => n332, C => n16, Y => n335);
   U555 : NAND2X1 port map( A => n207, B => n370, Y => n334);
   U556 : NAND3X1 port map( A => n336, B => n335, C => n334, Y => n337);
   U557 : MUX2X1 port map( B => n337, A => n219, S => n1498, Y => n338);
   U558 : NAND2X1 port map( A => n339, B => n338, Y => n1605);
   U559 : NAND2X1 port map( A => n1475, B => n219, Y => n360);
   U560 : INVX2 port map( A => n340, Y => n400);
   U561 : NAND2X1 port map( A => n400, B => n178, Y => n351);
   U562 : NOR2X1 port map( A => n160, B => n343, Y => n347);
   U563 : INVX2 port map( A => n1752, Y => n344);
   U564 : NAND3X1 port map( A => n418, B => n153, C => n344, Y => n345);
   U565 : OAI21X1 port map( A => n172, B => n380, C => n345, Y => n346);
   U567 : OAI21X1 port map( A => n347, B => n346, C => n27, Y => n350);
   U568 : NAND2X1 port map( A => n376, B => n205, Y => n348);
   U571 : NAND3X1 port map( A => n351, B => n350, C => n348, Y => n352);
   U572 : NAND2X1 port map( A => n16, B => n352, Y => n357);
   U573 : AND2X2 port map( A => currentPlainKey_5_port, B => n187, Y => n353);
   U574 : AOI21X1 port map( A => n195, B => n370, C => n353, Y => n355);
   U575 : NAND3X1 port map( A => n360, B => n357, C => n355, Y => n1606);
   U576 : AOI22X1 port map( A => currentPlainKey_6_port, B => n186, C => n376, 
                           D => n192, Y => n375);
   U577 : NAND2X1 port map( A => n400, B => n205, Y => n369);
   U578 : NAND2X1 port map( A => n2, B => n1474, Y => n392);
   U579 : INVX2 port map( A => n392, Y => n465);
   U582 : NAND2X1 port map( A => n465, B => n1132, Y => n364);
   U583 : NAND2X1 port map( A => n41, B => n153, Y => n394);
   U584 : INVX2 port map( A => n394, Y => n361);
   U585 : NAND2X1 port map( A => n1754, B => n361, Y => n363);
   U586 : AOI21X1 port map( A => n364, B => n363, C => n362, Y => n366);
   U587 : OAI22X1 port map( A => n160, B => n380, C => n1765, D => n168, Y => 
                           n365);
   U588 : OAI21X1 port map( A => n366, B => n365, C => n27, Y => n368);
   U589 : NAND2X1 port map( A => n422, B => n178, Y => n367);
   U590 : NAND3X1 port map( A => n369, B => n368, C => n367, Y => n373);
   U591 : MUX2X1 port map( B => n373, A => n219, S => n370, Y => n374);
   U592 : NAND2X1 port map( A => n375, B => n374, Y => n1607);
   U593 : AOI22X1 port map( A => currentPlainKey_7_port, B => n186, C => n376, 
                           D => n208, Y => n391);
   U594 : NAND2X1 port map( A => n422, B => n205, Y => n383);
   U596 : NOR2X1 port map( A => n1765, B => n161, Y => n378);
   U597 : OAI22X1 port map( A => n173, B => n392, C => n1758, D => n394, Y => 
                           n377);
   U600 : OAI21X1 port map( A => n378, B => n377, C => n418, Y => n382);
   U601 : INVX2 port map( A => n380, Y => n437);
   U602 : NAND2X1 port map( A => n437, B => n178, Y => n381);
   U603 : NAND3X1 port map( A => n383, B => n382, C => n381, Y => n385);
   U604 : NAND2X1 port map( A => n27, B => n385, Y => n390);
   U605 : NAND2X1 port map( A => n400, B => n197, Y => n387);
   U606 : NAND3X1 port map( A => n391, B => n390, C => n387, Y => n1608);
   U607 : AOI22X1 port map( A => currentPlainKey_8_port, B => n187, C => n422, 
                           D => n192, Y => n406);
   U608 : NAND2X1 port map( A => n184, B => n1472, Y => n399);
   U611 : OAI22X1 port map( A => n160, B => n392, C => n1771, D => n168, Y => 
                           n396);
   U612 : NAND2X1 port map( A => n2, B => n7, Y => n444);
   U613 : NAND2X1 port map( A => n1771, B => n444, Y => n427);
   U614 : INVX2 port map( A => n427, Y => n481);
   U615 : NAND2X1 port map( A => n1761, B => n481, Y => n393);
   U616 : OAI22X1 port map( A => n133, B => n444, C => n394, D => n393, Y => 
                           n395);
   U617 : OAI21X1 port map( A => n396, B => n395, C => n418, Y => n398);
   U618 : NAND2X1 port map( A => n437, B => n205, Y => n397);
   U619 : NAND3X1 port map( A => n399, B => n398, C => n397, Y => n404);
   U620 : MUX2X1 port map( B => n404, A => n219, S => n400, Y => n405);
   U621 : NAND2X1 port map( A => n406, B => n405, Y => n1609);
   U622 : NAND2X1 port map( A => n437, B => n197, Y => n425);
   U623 : NAND2X1 port map( A => n465, B => n178, Y => n414);
   U625 : NOR2X1 port map( A => n1771, B => n161, Y => n411);
   U626 : INVX2 port map( A => n1764, Y => n407);
   U629 : NAND3X1 port map( A => n481, B => n153, C => n407, Y => n408);
   U630 : OAI21X1 port map( A => n173, B => n444, C => n408, Y => n409);
   U631 : OAI21X1 port map( A => n411, B => n409, C => n41, Y => n413);
   U632 : NAND2X1 port map( A => n206, B => n1472, Y => n412);
   U633 : NAND3X1 port map( A => n414, B => n413, C => n412, Y => n416);
   U634 : NAND2X1 port map( A => n418, B => n416, Y => n424);
   U635 : AND2X2 port map( A => currentPlainKey_9_port, B => n187, Y => n419);
   U636 : AOI21X1 port map( A => n422, B => n209, C => n419, Y => n423);
   U637 : NAND3X1 port map( A => n425, B => n424, C => n423, Y => n1610);
   U640 : AOI22X1 port map( A => currentPlainKey_10_port, B => n185, C => n192,
                           D => n1472, Y => n440);
   U641 : NAND2X1 port map( A => n184, B => n1471, Y => n436);
   U642 : NAND2X1 port map( A => n81, B => n917, Y => n455);
   U643 : INVX2 port map( A => n455, Y => n526);
   U644 : NAND2X1 port map( A => n526, B => n1132, Y => n429);
   U645 : NAND2X1 port map( A => n33, B => n153, Y => n457);
   U646 : INVX2 port map( A => n457, Y => n426);
   U647 : NAND2X1 port map( A => n1767, B => n426, Y => n428);
   U648 : AOI21X1 port map( A => n429, B => n428, C => n427, Y => n431);
   U649 : OAI22X1 port map( A => n160, B => n444, C => n1777, D => n168, Y => 
                           n430);
   U650 : OAI21X1 port map( A => n431, B => n430, C => n41, Y => n435);
   U651 : NAND2X1 port map( A => n465, B => n205, Y => n432);
   U652 : NAND3X1 port map( A => n436, B => n435, C => n432, Y => n438);
   U654 : MUX2X1 port map( B => n438, A => n219, S => n437, Y => n439);
   U655 : NAND2X1 port map( A => n440, B => n439, Y => n1611);
   U656 : AOI22X1 port map( A => currentPlainKey_11_port, B => n186, C => n208,
                           D => n1472, Y => n454);
   U657 : NAND2X1 port map( A => n206, B => n1471, Y => n448);
   U660 : NOR2X1 port map( A => n1777, B => n161, Y => n443);
   U661 : OAI22X1 port map( A => n173, B => n455, C => n1770, D => n457, Y => 
                           n441);
   U662 : OAI21X1 port map( A => n443, B => n441, C => n481, Y => n446);
   U663 : INVX2 port map( A => n444, Y => n498);
   U664 : NAND2X1 port map( A => n498, B => n178, Y => n445);
   U665 : NAND3X1 port map( A => n448, B => n446, C => n445, Y => n450);
   U666 : NAND2X1 port map( A => n41, B => n450, Y => n453);
   U667 : NAND2X1 port map( A => n465, B => n197, Y => n452);
   U668 : NAND3X1 port map( A => n454, B => n453, C => n452, Y => n1612);
   U671 : AOI22X1 port map( A => currentPlainKey_12_port, B => n186, C => n192,
                           D => n1471, Y => n468);
   U673 : NAND2X1 port map( A => n184, B => n1470, Y => n462);
   U674 : OAI22X1 port map( A => n158, B => n455, C => n1783, D => n168, Y => 
                           n459);
   U675 : NAND2X1 port map( A => n81, B => n8, Y => n507);
   U676 : NAND2X1 port map( A => n1783, B => n507, Y => n487);
   U677 : INVX2 port map( A => n487, Y => n541);
   U678 : NAND2X1 port map( A => n1773, B => n541, Y => n456);
   U679 : OAI22X1 port map( A => n133, B => n507, C => n457, D => n456, Y => 
                           n458);
   U680 : OAI21X1 port map( A => n459, B => n458, C => n481, Y => n461);
   U681 : NAND2X1 port map( A => n498, B => n205, Y => n460);
   U682 : NAND3X1 port map( A => n462, B => n461, C => n460, Y => n466);
   U683 : MUX2X1 port map( B => n466, A => n219, S => n465, Y => n467);
   U684 : NAND2X1 port map( A => n468, B => n467, Y => n1613);
   U685 : NAND2X1 port map( A => n498, B => n197, Y => n485);
   U687 : NAND2X1 port map( A => n526, B => n178, Y => n479);
   U688 : NOR2X1 port map( A => n1783, B => n161, Y => n473);
   U691 : INVX2 port map( A => n1776, Y => n469);
   U692 : NAND3X1 port map( A => n541, B => n153, C => n469, Y => n471);
   U693 : OAI21X1 port map( A => n173, B => n507, C => n471, Y => n472);
   U694 : OAI21X1 port map( A => n473, B => n472, C => n33, Y => n476);
   U695 : NAND2X1 port map( A => n206, B => n1470, Y => n474);
   U696 : NAND3X1 port map( A => n479, B => n476, C => n474, Y => n480);
   U697 : NAND2X1 port map( A => n481, B => n480, Y => n484);
   U698 : AND2X2 port map( A => currentPlainKey_13_port, B => n185, Y => n482);
   U699 : AOI21X1 port map( A => n209, B => n1471, C => n482, Y => n483);
   U702 : NAND3X1 port map( A => n485, B => n484, C => n483, Y => n1614);
   U703 : AOI22X1 port map( A => currentPlainKey_14_port, B => n187, C => n192,
                           D => n1470, Y => n501);
   U704 : NAND2X1 port map( A => n184, B => n1469, Y => n496);
   U705 : NAND2X1 port map( A => n81, B => n20, Y => n515);
   U706 : INVX2 port map( A => n515, Y => n590);
   U707 : NAND2X1 port map( A => n590, B => n1132, Y => n489);
   U708 : NAND2X1 port map( A => n35, B => n153, Y => n519);
   U709 : INVX2 port map( A => n519, Y => n486);
   U710 : NAND2X1 port map( A => n1779, B => n486, Y => n488);
   U711 : AOI21X1 port map( A => n489, B => n488, C => n487, Y => n493);
   U712 : OAI22X1 port map( A => n158, B => n507, C => n1789, D => n168, Y => 
                           n492);
   U713 : OAI21X1 port map( A => n493, B => n492, C => n33, Y => n495);
   U714 : NAND2X1 port map( A => n526, B => n205, Y => n494);
   U716 : NAND3X1 port map( A => n496, B => n495, C => n494, Y => n499);
   U717 : MUX2X1 port map( B => n499, A => n219, S => n498, Y => n500);
   U720 : NAND2X1 port map( A => n501, B => n500, Y => n1615);
   U721 : AOI22X1 port map( A => currentPlainKey_15_port, B => n186, C => n208,
                           D => n1470, Y => n514);
   U722 : NAND2X1 port map( A => n206, B => n1469, Y => n510);
   U723 : NOR2X1 port map( A => n1789, B => n160, Y => n506);
   U724 : OAI22X1 port map( A => n173, B => n515, C => n1782, D => n519, Y => 
                           n503);
   U725 : OAI21X1 port map( A => n506, B => n503, C => n541, Y => n509);
   U726 : INVX2 port map( A => n507, Y => n561);
   U727 : NAND2X1 port map( A => n561, B => n178, Y => n508);
   U728 : NAND3X1 port map( A => n510, B => n509, C => n508, Y => n511);
   U731 : NAND2X1 port map( A => n33, B => n511, Y => n513);
   U732 : NAND2X1 port map( A => n526, B => n197, Y => n512);
   U733 : NAND3X1 port map( A => n514, B => n513, C => n512, Y => n1616);
   U734 : AOI22X1 port map( A => currentPlainKey_16_port, B => n186, C => n193,
                           D => n1469, Y => n530);
   U735 : NAND2X1 port map( A => n184, B => n1468, Y => n525);
   U736 : OAI22X1 port map( A => n158, B => n515, C => n1795_port, D => n172, Y
                           => n521);
   U737 : NAND2X1 port map( A => n81, B => n23, Y => n568);
   U738 : NAND2X1 port map( A => n1795_port, B => n568, Y => n550);
   U739 : INVX2 port map( A => n550, Y => n604);
   U740 : NAND2X1 port map( A => n1785, B => n604, Y => n516);
   U741 : OAI22X1 port map( A => n135, B => n568, C => n519, D => n516, Y => 
                           n520);
   U742 : OAI21X1 port map( A => n521, B => n520, C => n541, Y => n523);
   U743 : NAND2X1 port map( A => n561, B => n205, Y => n522);
   U745 : NAND3X1 port map( A => n525, B => n523, C => n522, Y => n527);
   U746 : MUX2X1 port map( B => n527, A => n219, S => n526, Y => n528);
   U749 : NAND2X1 port map( A => n530, B => n528, Y => n1617);
   U750 : NAND2X1 port map( A => n561, B => n197, Y => n548);
   U751 : NAND2X1 port map( A => n590, B => n178, Y => n539);
   U752 : NOR2X1 port map( A => n1795_port, B => n160, Y => n536);
   U753 : INVX2 port map( A => n1788, Y => n533);
   U754 : NAND3X1 port map( A => n604, B => n153, C => n533, Y => n534);
   U755 : OAI21X1 port map( A => n173, B => n568, C => n534, Y => n535);
   U756 : OAI21X1 port map( A => n536, B => n535, C => n35, Y => n538);
   U757 : NAND2X1 port map( A => n206, B => n1468, Y => n537);
   U760 : NAND3X1 port map( A => n539, B => n538, C => n537, Y => n540);
   U761 : NAND2X1 port map( A => n541, B => n540, Y => n547);
   U762 : AND2X2 port map( A => currentPlainKey_17_port, B => n186, Y => n542);
   U763 : AOI21X1 port map( A => n209, B => n1469, C => n542, Y => n543);
   U764 : NAND3X1 port map( A => n548, B => n547, C => n543, Y => n1618);
   U765 : AOI22X1 port map( A => currentPlainKey_18_port, B => n186, C => n192,
                           D => n1468, Y => n565);
   U766 : NAND2X1 port map( A => n184, B => n1467, Y => n559);
   U767 : NAND2X1 port map( A => n4, B => n119, Y => n578);
   U768 : INVX2 port map( A => n578, Y => n650);
   U769 : NAND2X1 port map( A => n650, B => n1132, Y => n552);
   U770 : NAND2X1 port map( A => n43, B => n153, Y => n580);
   U771 : INVX2 port map( A => n580, Y => n549);
   U772 : NAND2X1 port map( A => n1791, B => n549, Y => n551);
   U774 : AOI21X1 port map( A => n552, B => n551, C => n550, Y => n555);
   U775 : OAI22X1 port map( A => n158, B => n568, C => n1801, D => n168, Y => 
                           n554);
   U778 : OAI21X1 port map( A => n555, B => n554, C => n35, Y => n557);
   U779 : NAND2X1 port map( A => n590, B => n205, Y => n556);
   U780 : NAND3X1 port map( A => n559, B => n557, C => n556, Y => n563);
   U781 : MUX2X1 port map( B => n563, A => n217, S => n561, Y => n564);
   U782 : NAND2X1 port map( A => n565, B => n564, Y => n1619);
   U783 : AOI22X1 port map( A => currentPlainKey_19_port, B => n186, C => n208,
                           D => n1468, Y => n577);
   U784 : NAND2X1 port map( A => n206, B => n1467, Y => n571);
   U785 : NOR2X1 port map( A => n1801, B => n160, Y => n567);
   U786 : OAI22X1 port map( A => n71, B => n578, C => n1794_port, D => n580, Y 
                           => n566);
   U789 : OAI21X1 port map( A => n567, B => n566, C => n604, Y => n570);
   U790 : INVX2 port map( A => n568, Y => n622);
   U791 : NAND2X1 port map( A => n622, B => n180, Y => n569);
   U792 : NAND3X1 port map( A => n571, B => n570, C => n569, Y => n572);
   U793 : NAND2X1 port map( A => n35, B => n572, Y => n576);
   U794 : NAND2X1 port map( A => n590, B => n197, Y => n573);
   U795 : NAND3X1 port map( A => n577, B => n576, C => n573, Y => n1620);
   U796 : AOI22X1 port map( A => currentPlainKey_20_port, B => n186, C => n193,
                           D => n1467, Y => n593);
   U797 : NAND2X1 port map( A => n184, B => n1466, Y => n587);
   U798 : OAI22X1 port map( A => n158, B => n578, C => n1807, D => n172, Y => 
                           n583);
   U799 : NAND2X1 port map( A => n4, B => n1477, Y => n630);
   U800 : NAND2X1 port map( A => n1807, B => n630, Y => n611);
   U801 : INVX2 port map( A => n611, Y => n665);
   U802 : NAND2X1 port map( A => n1797_port, B => n665, Y => n579);
   U804 : OAI22X1 port map( A => n135, B => n630, C => n580, D => n579, Y => 
                           n582);
   U805 : OAI21X1 port map( A => n583, B => n582, C => n604, Y => n585);
   U808 : NAND2X1 port map( A => n622, B => n205, Y => n584);
   U809 : NAND3X1 port map( A => n587, B => n585, C => n584, Y => n591);
   U810 : MUX2X1 port map( B => n591, A => n217, S => n590, Y => n592);
   U811 : NAND2X1 port map( A => n593, B => n592, Y => n1621);
   U812 : NAND2X1 port map( A => n622, B => n197, Y => n609);
   U813 : NAND2X1 port map( A => n650, B => n180, Y => n600);
   U814 : NOR2X1 port map( A => n1807, B => n160, Y => n597);
   U815 : INVX2 port map( A => n1800, Y => n594);
   U816 : NAND3X1 port map( A => n665, B => n153, C => n594, Y => n595);
   U819 : OAI21X1 port map( A => n173, B => n630, C => n595, Y => n596);
   U820 : OAI21X1 port map( A => n597, B => n596, C => n43, Y => n599);
   U821 : NAND2X1 port map( A => n205, B => n1466, Y => n598);
   U822 : NAND3X1 port map( A => n600, B => n599, C => n598, Y => n603);
   U823 : NAND2X1 port map( A => n604, B => n603, Y => n607);
   U824 : AND2X2 port map( A => currentPlainKey_21_port, B => n187, Y => n605);
   U825 : AOI21X1 port map( A => n209, B => n1467, C => n605, Y => n606);
   U826 : NAND3X1 port map( A => n609, B => n607, C => n606, Y => n1622);
   U827 : AOI22X1 port map( A => currentPlainKey_22_port, B => n186, C => n193,
                           D => n1466, Y => n625);
   U828 : NAND2X1 port map( A => n183, B => n1465, Y => n621);
   U829 : NAND2X1 port map( A => n4, B => n1474, Y => n639);
   U830 : INVX2 port map( A => n639, Y => n710);
   U831 : NAND2X1 port map( A => n710, B => n1132, Y => n614);
   U833 : NAND2X1 port map( A => n45, B => n153, Y => n644);
   U834 : INVX2 port map( A => n644, Y => n610);
   U837 : NAND2X1 port map( A => n1803, B => n610, Y => n612);
   U838 : AOI21X1 port map( A => n614, B => n612, C => n611, Y => n618);
   U839 : OAI22X1 port map( A => n158, B => n630, C => n1814, D => n172, Y => 
                           n617);
   U840 : OAI21X1 port map( A => n618, B => n617, C => n43, Y => n620);
   U841 : NAND2X1 port map( A => n650, B => n205, Y => n619);
   U842 : NAND3X1 port map( A => n621, B => n620, C => n619, Y => n623);
   U843 : MUX2X1 port map( B => n623, A => n217, S => n622, Y => n624);
   U844 : NAND2X1 port map( A => n625, B => n624, Y => n1623);
   U845 : AOI22X1 port map( A => currentPlainKey_23_port, B => n186, C => n208,
                           D => n1466, Y => n638);
   U848 : NAND2X1 port map( A => n205, B => n1465, Y => n633);
   U849 : NOR2X1 port map( A => n1814, B => n160, Y => n627);
   U850 : OAI22X1 port map( A => n71, B => n639, C => n1806, D => n644, Y => 
                           n626);
   U851 : OAI21X1 port map( A => n627, B => n626, C => n665, Y => n632);
   U852 : INVX2 port map( A => n630, Y => n682);
   U853 : NAND2X1 port map( A => n682, B => n180, Y => n631);
   U854 : NAND3X1 port map( A => n633, B => n632, C => n631, Y => n634);
   U855 : NAND2X1 port map( A => n43, B => n634, Y => n637);
   U856 : NAND2X1 port map( A => n650, B => n197, Y => n636);
   U857 : NAND3X1 port map( A => n638, B => n637, C => n636, Y => n1624);
   U858 : AOI22X1 port map( A => currentPlainKey_24_port, B => n186, C => n193,
                           D => n1465, Y => n653);
   U859 : NAND2X1 port map( A => n183, B => n1464, Y => n649);
   U860 : OAI22X1 port map( A => n158, B => n639, C => n1820, D => n172, Y => 
                           n646);
   U862 : NAND2X1 port map( A => n4, B => n7, Y => n690);
   U863 : NAND2X1 port map( A => n1820, B => n690, Y => n674);
   U866 : INVX2 port map( A => n674, Y => n728);
   U867 : NAND2X1 port map( A => n1810, B => n728, Y => n641);
   U868 : OAI22X1 port map( A => n135, B => n690, C => n644, D => n641, Y => 
                           n645);
   U869 : OAI21X1 port map( A => n646, B => n645, C => n665, Y => n648);
   U870 : NAND2X1 port map( A => n682, B => n205, Y => n647);
   U871 : NAND3X1 port map( A => n649, B => n648, C => n647, Y => n651);
   U872 : MUX2X1 port map( B => n651, A => n217, S => n650, Y => n652);
   U873 : NAND2X1 port map( A => n653, B => n652, Y => n1625);
   U874 : NAND2X1 port map( A => n682, B => n195, Y => n670);
   U877 : NAND2X1 port map( A => n710, B => n180, Y => n662);
   U878 : NOR2X1 port map( A => n1820, B => n160, Y => n659);
   U879 : INVX2 port map( A => n1813, Y => n654);
   U880 : NAND3X1 port map( A => n728, B => n153, C => n654, Y => n657);
   U881 : OAI21X1 port map( A => n173, B => n690, C => n657, Y => n658);
   U882 : OAI21X1 port map( A => n659, B => n658, C => n45, Y => n661);
   U883 : NAND2X1 port map( A => n206, B => n1464, Y => n660);
   U884 : NAND3X1 port map( A => n662, B => n661, C => n660, Y => n663);
   U885 : NAND2X1 port map( A => n665, B => n663, Y => n668);
   U886 : AND2X2 port map( A => currentPlainKey_25_port, B => n187, Y => n666);
   U887 : AOI21X1 port map( A => n209, B => n1465, C => n666, Y => n667);
   U888 : NAND3X1 port map( A => n670, B => n668, C => n667, Y => n1626);
   U889 : AOI22X1 port map( A => currentPlainKey_26_port, B => n186, C => n193,
                           D => n1464, Y => n687);
   U891 : NAND2X1 port map( A => n183, B => n1463, Y => n681);
   U892 : NAND2X1 port map( A => n83, B => n917, Y => n702);
   U893 : INVX2 port map( A => n702, Y => n773);
   U894 : NAND2X1 port map( A => n773, B => n1132, Y => n676);
   U897 : NAND2X1 port map( A => n37, B => n153, Y => n704);
   U898 : INVX2 port map( A => n704, Y => n672);
   U899 : NAND2X1 port map( A => n1816, B => n672, Y => n675);
   U900 : AOI21X1 port map( A => n676, B => n675, C => n674, Y => n678);
   U901 : OAI22X1 port map( A => n158, B => n690, C => n1826, D => n172, Y => 
                           n677);
   U902 : OAI21X1 port map( A => n678, B => n677, C => n45, Y => n680);
   U903 : NAND2X1 port map( A => n710, B => n205, Y => n679);
   U904 : NAND3X1 port map( A => n681, B => n680, C => n679, Y => n683);
   U905 : MUX2X1 port map( B => n683, A => n217, S => n682, Y => n684);
   U908 : NAND2X1 port map( A => n687, B => n684, Y => n1627);
   U910 : AOI22X1 port map( A => currentPlainKey_27_port, B => n186, C => n208,
                           D => n1464, Y => n701);
   U911 : NAND2X1 port map( A => n206, B => n1463, Y => n694_port);
   U912 : NOR2X1 port map( A => n1826, B => n161, Y => n689);
   U913 : OAI22X1 port map( A => n71, B => n702, C => n1819, D => n704, Y => 
                           n688);
   U914 : OAI21X1 port map( A => n689, B => n688, C => n728, Y => n693);
   U915 : INVX2 port map( A => n690, Y => n744);
   U916 : NAND2X1 port map( A => n744, B => n178, Y => n691);
   U917 : NAND3X1 port map( A => n694_port, B => n693, C => n691, Y => n695);
   U918 : NAND2X1 port map( A => n45, B => n695, Y => n698);
   U919 : NAND2X1 port map( A => n710, B => n195, Y => n696);
   U920 : NAND3X1 port map( A => n701, B => n698, C => n696, Y => n1628);
   U921 : AOI22X1 port map( A => currentPlainKey_28_port, B => n185, C => n193,
                           D => n1463, Y => n715);
   U922 : NAND2X1 port map( A => n183, B => n1462, Y => n709);
   U924 : OAI22X1 port map( A => n158, B => n702, C => n1832, D => n172, Y => 
                           n706);
   U925 : NAND2X1 port map( A => n83, B => n8, Y => n752);
   U928 : NAND2X1 port map( A => n1832, B => n752, Y => n734);
   U929 : INVX2 port map( A => n734, Y => n789);
   U930 : NAND2X1 port map( A => n1822, B => n789, Y => n703);
   U931 : OAI22X1 port map( A => n135, B => n752, C => n704, D => n703, Y => 
                           n705);
   U932 : OAI21X1 port map( A => n706, B => n705, C => n728, Y => n708);
   U933 : NAND2X1 port map( A => n744, B => n205, Y => n707);
   U934 : NAND3X1 port map( A => n709, B => n708, C => n707, Y => n711);
   U935 : MUX2X1 port map( B => n711, A => n217, S => n710, Y => n714);
   U936 : NAND2X1 port map( A => n715, B => n714, Y => n1629);
   U939 : NAND2X1 port map( A => n744, B => n195, Y => n732);
   U940 : NAND2X1 port map( A => n773, B => n180, Y => n723);
   U941 : NOR2X1 port map( A => n1832, B => n160, Y => n720);
   U942 : INVX2 port map( A => n1825, Y => n716);
   U943 : NAND3X1 port map( A => n789, B => n153, C => n716, Y => n717);
   U944 : OAI21X1 port map( A => n173, B => n752, C => n717, Y => n718);
   U945 : OAI21X1 port map( A => n720, B => n718, C => n37, Y => n722);
   U946 : NAND2X1 port map( A => n205, B => n1462, Y => n721);
   U947 : NAND3X1 port map( A => n723, B => n722, C => n721, Y => n725);
   U948 : NAND2X1 port map( A => n728, B => n725, Y => n731);
   U949 : AND2X2 port map( A => currentPlainKey_29_port, B => n187, Y => n729);
   U950 : AOI21X1 port map( A => n209, B => n1463, C => n729, Y => n730);
   U951 : NAND3X1 port map( A => n732, B => n731, C => n730, Y => n1630);
   U953 : AOI22X1 port map( A => currentPlainKey_30_port, B => n185, C => n195,
                           D => n1462, Y => n748);
   U954 : NAND2X1 port map( A => n183, B => n1461, Y => n743);
   U957 : NAND2X1 port map( A => n83, B => n20, Y => n762);
   U958 : INVX2 port map( A => n762, Y => n834);
   U959 : NAND2X1 port map( A => n834, B => n1132, Y => n736);
   U960 : NAND2X1 port map( A => n39, B => n153, Y => n764);
   U961 : INVX2 port map( A => n764, Y => n733);
   U962 : NAND2X1 port map( A => n1828, B => n733, Y => n735);
   U963 : AOI21X1 port map( A => n736, B => n735, C => n734, Y => n738);
   U964 : OAI22X1 port map( A => n158, B => n752, C => n1838, D => n71, Y => 
                           n737);
   U965 : OAI21X1 port map( A => n738, B => n737, C => n37, Y => n742);
   U968 : NAND2X1 port map( A => n773, B => n203, Y => n741);
   U969 : NAND3X1 port map( A => n743, B => n742, C => n741, Y => n745);
   U970 : MUX2X1 port map( B => n745, A => n217, S => n744, Y => n747);
   U971 : NAND2X1 port map( A => n748, B => n747, Y => n1631);
   U972 : AOI22X1 port map( A => currentPlainKey_31_port, B => n185, C => n208,
                           D => n1462, Y => n761);
   U973 : NAND2X1 port map( A => n206, B => n1461, Y => n757);
   U974 : NOR2X1 port map( A => n1838, B => n160, Y => n750);
   U975 : OAI22X1 port map( A => n71, B => n762, C => n1831, D => n764, Y => 
                           n749);
   U976 : OAI21X1 port map( A => n750, B => n749, C => n789, Y => n756);
   U977 : INVX2 port map( A => n752, Y => n806);
   U978 : NAND2X1 port map( A => n806, B => n181, Y => n755);
   U979 : NAND3X1 port map( A => n757, B => n756, C => n755, Y => n758);
   U980 : NAND2X1 port map( A => n37, B => n758, Y => n760);
   U982 : NAND2X1 port map( A => n773, B => n195, Y => n759);
   U983 : NAND3X1 port map( A => n761, B => n760, C => n759, Y => n1632);
   U986 : AOI22X1 port map( A => currentPlainKey_32_port, B => n185, C => n195,
                           D => n1461, Y => n777);
   U987 : NAND2X1 port map( A => n183, B => n1460, Y => n772);
   U988 : OAI22X1 port map( A => n158, B => n762, C => n1844, D => n172, Y => 
                           n769);
   U989 : NAND2X1 port map( A => n83, B => n23, Y => n815);
   U990 : NAND2X1 port map( A => n1844, B => n815, Y => n795);
   U991 : INVX2 port map( A => n795, Y => n849);
   U992 : NAND2X1 port map( A => n1834, B => n849, Y => n763);
   U993 : OAI22X1 port map( A => n135, B => n815, C => n764, D => n763, Y => 
                           n765);
   U994 : OAI21X1 port map( A => n769, B => n765, C => n789, Y => n771);
   U997 : NAND2X1 port map( A => n806, B => n203, Y => n770);
   U998 : NAND3X1 port map( A => n772, B => n771, C => n770, Y => n774);
   U999 : MUX2X1 port map( B => n774, A => n217, S => n773, Y => n776);
   U1000 : NAND2X1 port map( A => n777, B => n776, Y => n1633);
   U1001 : NAND2X1 port map( A => n806, B => n195, Y => n793);
   U1002 : NAND2X1 port map( A => n834, B => n181, Y => n787);
   U1003 : NOR2X1 port map( A => n1844, B => n160, Y => n783);
   U1004 : INVX2 port map( A => n1837, Y => n778);
   U1005 : NAND3X1 port map( A => n849, B => n153, C => n778, Y => n779);
   U1006 : OAI21X1 port map( A => n173, B => n815, C => n779, Y => n781);
   U1007 : OAI21X1 port map( A => n783, B => n781, C => n39, Y => n786);
   U1008 : NAND2X1 port map( A => n206, B => n1460, Y => n785);
   U1009 : NAND3X1 port map( A => n787, B => n786, C => n785, Y => n788);
   U1011 : NAND2X1 port map( A => n789, B => n788, Y => n792);
   U1012 : AND2X2 port map( A => currentPlainKey_33_port, B => n187, Y => n790)
                           ;
   U1013 : AOI21X1 port map( A => n209, B => n1461, C => n790, Y => n791);
   U1016 : NAND3X1 port map( A => n793, B => n792, C => n791, Y => n1634);
   U1017 : AOI22X1 port map( A => currentPlainKey_34_port, B => n185, C => n193
                           , D => n1460, Y => n812);
   U1018 : NAND2X1 port map( A => n183, B => n1459, Y => n805);
   U1019 : NAND2X1 port map( A => n1, B => n119, Y => n825);
   U1020 : INVX2 port map( A => n825, Y => n897);
   U1021 : NAND2X1 port map( A => n897, B => n1132, Y => n799);
   U1022 : NAND2X1 port map( A => n47, B => n153, Y => n827);
   U1023 : INVX2 port map( A => n827, Y => n794);
   U1024 : NAND2X1 port map( A => n1840, B => n794, Y => n798);
   U1027 : AOI21X1 port map( A => n799, B => n798, C => n795, Y => n801);
   U1028 : OAI22X1 port map( A => n158, B => n815, C => n1850, D => n172, Y => 
                           n800);
   U1029 : OAI21X1 port map( A => n801, B => n800, C => n39, Y => n804);
   U1030 : NAND2X1 port map( A => n834, B => n203, Y => n802);
   U1031 : NAND3X1 port map( A => n805, B => n804, C => n802, Y => n807);
   U1032 : MUX2X1 port map( B => n807, A => n217, S => n806, Y => n809);
   U1033 : NAND2X1 port map( A => n812, B => n809, Y => n1635);
   U1034 : AOI22X1 port map( A => currentPlainKey_35_port, B => n185, C => n209
                           , D => n1460, Y => n822);
   U1035 : NAND2X1 port map( A => n206, B => n1459, Y => n818);
   U1036 : NOR2X1 port map( A => n1850, B => n160, Y => n814);
   U1037 : OAI22X1 port map( A => n71, B => n825, C => n1843, D => n827, Y => 
                           n813);
   U1038 : OAI21X1 port map( A => n814, B => n813, C => n849, Y => n817);
   U1039 : INVX2 port map( A => n815, Y => n869);
   U1040 : NAND2X1 port map( A => n869, B => n180, Y => n816);
   U1042 : NAND3X1 port map( A => n818, B => n817, C => n816, Y => n819);
   U1043 : NAND2X1 port map( A => n39, B => n819, Y => n821);
   U1047 : NAND2X1 port map( A => n834, B => n195, Y => n820);
   U1048 : NAND3X1 port map( A => n822, B => n821, C => n820, Y => n1636);
   U1049 : AOI22X1 port map( A => currentPlainKey_36_port, B => n185, C => n195
                           , D => n1459, Y => n840);
   U1050 : NAND2X1 port map( A => n183, B => n1458, Y => n833);
   U1051 : OAI22X1 port map( A => n156, B => n825, C => n1856, D => n172, Y => 
                           n829);
   U1052 : NAND2X1 port map( A => n1, B => n1477, Y => n875);
   U1053 : NAND2X1 port map( A => n1856, B => n875, Y => n858);
   U1054 : INVX2 port map( A => n858, Y => n911);
   U1055 : NAND2X1 port map( A => n1846, B => n911, Y => n826);
   U1056 : OAI22X1 port map( A => n135, B => n875, C => n827, D => n826, Y => 
                           n828);
   U1060 : OAI21X1 port map( A => n829, B => n828, C => n849, Y => n832);
   U1061 : NAND2X1 port map( A => n869, B => n203, Y => n831);
   U1062 : NAND3X1 port map( A => n833, B => n832, C => n831, Y => n836);
   U1063 : MUX2X1 port map( B => n836, A => n217, S => n834, Y => n839);
   U1064 : NAND2X1 port map( A => n840, B => n839, Y => n1637);
   U1065 : NAND2X1 port map( A => n869, B => n195, Y => n855);
   U1066 : NAND2X1 port map( A => n897, B => n181, Y => n847);
   U1067 : NOR2X1 port map( A => n1856, B => n161, Y => n844);
   U1068 : INVX2 port map( A => n1849, Y => n841);
   U1069 : NAND3X1 port map( A => n911, B => n153, C => n841, Y => n842);
   U1070 : OAI21X1 port map( A => n168, B => n875, C => n842, Y => n843);
   U1071 : OAI21X1 port map( A => n844, B => n843, C => n47, Y => n846);
   U1072 : NAND2X1 port map( A => n206, B => n1458, Y => n845);
   U1073 : NAND3X1 port map( A => n847, B => n846, C => n845, Y => n848);
   U1075 : NAND2X1 port map( A => n849, B => n848, Y => n854);
   U1076 : AND2X2 port map( A => currentPlainKey_37_port, B => n186, Y => n852)
                           ;
   U1080 : AOI21X1 port map( A => n210, B => n1459, C => n852, Y => n853);
   U1081 : NAND3X1 port map( A => n855, B => n854, C => n853, Y => n1638);
   U1082 : AOI22X1 port map( A => currentPlainKey_38_port, B => n185, C => n193
                           , D => n1458, Y => n872);
   U1083 : NAND2X1 port map( A => n183, B => n1457, Y => n868);
   U1084 : NAND2X1 port map( A => n1, B => n1474, Y => n885);
   U1085 : INVX2 port map( A => n885, Y => n958);
   U1086 : NAND2X1 port map( A => n958, B => n1132, Y => n860);
   U1087 : NAND2X1 port map( A => n49, B => n153, Y => n888);
   U1088 : INVX2 port map( A => n888, Y => n856);
   U1089 : NAND2X1 port map( A => n1852, B => n856, Y => n859);
   U1093 : AOI21X1 port map( A => n860, B => n859, C => n858, Y => n863);
   U1094 : OAI22X1 port map( A => n156, B => n875, C => n1863, D => n172, Y => 
                           n861);
   U1095 : OAI21X1 port map( A => n863, B => n861, C => n47, Y => n867);
   U1096 : NAND2X1 port map( A => n897, B => n203, Y => n866);
   U1097 : NAND3X1 port map( A => n868, B => n867, C => n866, Y => n870);
   U1098 : MUX2X1 port map( B => n870, A => n217, S => n869, Y => n871);
   U1099 : NAND2X1 port map( A => n872, B => n871, Y => n1639);
   U1100 : AOI22X1 port map( A => currentPlainKey_39_port, B => n185, C => n208
                           , D => n1458, Y => n884);
   U1101 : NAND2X1 port map( A => n206, B => n1457, Y => n880);
   U1102 : NOR2X1 port map( A => n1863, B => n161, Y => n874);
   U1103 : OAI22X1 port map( A => n173, B => n885, C => n1855, D => n888, Y => 
                           n873);
   U1104 : OAI21X1 port map( A => n874, B => n873, C => n911, Y => n879);
   U1105 : INVX2 port map( A => n875, Y => n930);
   U1106 : NAND2X1 port map( A => n930, B => n181, Y => n876);
   U1107 : NAND3X1 port map( A => n880, B => n879, C => n876, Y => n881);
   U1108 : NAND2X1 port map( A => n47, B => n881, Y => n883);
   U1109 : NAND2X1 port map( A => n897, B => n195, Y => n882);
   U1110 : NAND3X1 port map( A => n884, B => n883, C => n882, Y => n1640);
   U1114 : AOI22X1 port map( A => currentPlainKey_40_port, B => n185, C => n193
                           , D => n1457, Y => n900);
   U1115 : NAND2X1 port map( A => n183, B => n1456, Y => n896);
   U1116 : OAI22X1 port map( A => n156, B => n885, C => n1869, D => n172, Y => 
                           n890);
   U1117 : NAND2X1 port map( A => n1, B => n7, Y => n938);
   U1118 : NAND2X1 port map( A => n1869, B => n938, Y => n920);
   U1119 : INVX2 port map( A => n920, Y => n974);
   U1120 : NAND2X1 port map( A => n1859, B => n974, Y => n887);
   U1121 : OAI22X1 port map( A => n135, B => n938, C => n888, D => n887, Y => 
                           n889);
   U1122 : OAI21X1 port map( A => n890, B => n889, C => n911, Y => n894);
   U1123 : NAND2X1 port map( A => n930, B => n203, Y => n892);
   U1124 : NAND3X1 port map( A => n896, B => n894, C => n892, Y => n898);
   U1125 : MUX2X1 port map( B => n898, A => n217, S => n897, Y => n899);
   U1129 : NAND2X1 port map( A => n900, B => n899, Y => n1641);
   U1130 : NAND2X1 port map( A => n930, B => n195, Y => n916);
   U1131 : NAND2X1 port map( A => n958, B => n180, Y => n909);
   U1132 : NOR2X1 port map( A => n1869, B => n161, Y => n904);
   U1133 : INVX2 port map( A => n1862, Y => n901);
   U1134 : NAND3X1 port map( A => n974, B => n153, C => n901, Y => n902);
   U1135 : OAI21X1 port map( A => n173, B => n938, C => n902, Y => n903);
   U1136 : OAI21X1 port map( A => n904, B => n903, C => n49, Y => n906);
   U1137 : NAND2X1 port map( A => n206, B => n1456, Y => n905);
   U1138 : NAND3X1 port map( A => n909, B => n906, C => n905, Y => n910);
   U1139 : NAND2X1 port map( A => n911, B => n910, Y => n915);
   U1140 : AND2X2 port map( A => currentPlainKey_41_port, B => n185, Y => n912)
                           ;
   U1141 : AOI21X1 port map( A => n210, B => n1457, C => n912, Y => n913);
   U1142 : NAND3X1 port map( A => n916, B => n915, C => n913, Y => n1642);
   U1143 : AOI22X1 port map( A => currentPlainKey_42_port, B => n185, C => n193
                           , D => n1456, Y => n933);
   U1144 : NAND2X1 port map( A => n183, B => n1455, Y => n929);
   U1145 : NAND2X1 port map( A => n79, B => n917, Y => n950);
   U1146 : INVX2 port map( A => n950, Y => n1021);
   U1147 : NAND2X1 port map( A => n1021, B => n1132, Y => n924);
   U1148 : NAND2X1 port map( A => n31, B => n153, Y => n952);
   U1149 : INVX2 port map( A => n952, Y => n918);
   U1150 : NAND2X1 port map( A => n1865, B => n918, Y => n923);
   U1151 : AOI21X1 port map( A => n924, B => n923, C => n920, Y => n926);
   U1152 : OAI22X1 port map( A => n156, B => n938, C => n1875, D => n172, Y => 
                           n925);
   U1153 : OAI21X1 port map( A => n926, B => n925, C => n49, Y => n928);
   U1158 : NAND2X1 port map( A => n958, B => n203, Y => n927);
   U1159 : NAND3X1 port map( A => n929, B => n928, C => n927, Y => n931);
   U1160 : MUX2X1 port map( B => n931, A => n210, S => n930, Y => n932);
   U1161 : NAND2X1 port map( A => n933, B => n932, Y => n1643);
   U1162 : AOI22X1 port map( A => currentPlainKey_43_port, B => n185, C => n209
                           , D => n1456, Y => n947);
   U1163 : NAND2X1 port map( A => n206, B => n1455, Y => n942);
   U1164 : NOR2X1 port map( A => n1875, B => n161, Y => n937);
   U1165 : OAI22X1 port map( A => n173, B => n950, C => n1868, D => n952, Y => 
                           n936);
   U1166 : OAI21X1 port map( A => n937, B => n936, C => n974, Y => n940);
   U1167 : INVX2 port map( A => n938, Y => n993);
   U1168 : NAND2X1 port map( A => n993, B => n181, Y => n939);
   U1169 : NAND3X1 port map( A => n942, B => n940, C => n939, Y => n943);
   U1170 : NAND2X1 port map( A => n49, B => n943, Y => n945);
   U1171 : NAND2X1 port map( A => n958, B => n195, Y => n944);
   U1172 : NAND3X1 port map( A => n947, B => n945, C => n944, Y => n1644);
   U1173 : AOI22X1 port map( A => currentPlainKey_44_port, B => n185, C => n193
                           , D => n1455, Y => n963);
   U1174 : NAND2X1 port map( A => n181, B => n1454, Y => n957);
   U1175 : OAI22X1 port map( A => n156, B => n950, C => n1881, D => n168, Y => 
                           n954);
   U1176 : NAND2X1 port map( A => n79, B => n8, Y => n999);
   U1177 : NAND2X1 port map( A => n1881, B => n999, Y => n982);
   U1178 : INVX2 port map( A => n982, Y => n1036);
   U1179 : NAND2X1 port map( A => n1871, B => n1036, Y => n951);
   U1180 : OAI22X1 port map( A => n135, B => n999, C => n952, D => n951, Y => 
                           n953);
   U1181 : OAI21X1 port map( A => n954, B => n953, C => n974, Y => n956);
   U1188 : NAND2X1 port map( A => n993, B => n203, Y => n955);
   U1191 : NAND3X1 port map( A => n957, B => n956, C => n955, Y => n959);
   U1192 : MUX2X1 port map( B => n959, A => n210, S => n958, Y => n960);
   U1193 : NAND2X1 port map( A => n963, B => n960, Y => n1645);
   U1194 : NAND2X1 port map( A => n993, B => n197, Y => n980);
   U1195 : NAND2X1 port map( A => n1021, B => n180, Y => n971);
   U1196 : NOR2X1 port map( A => n1881, B => n161, Y => n967);
   U1197 : INVX2 port map( A => n1874, Y => n964);
   U1198 : NAND3X1 port map( A => n1036, B => n153, C => n964, Y => n965);
   U1200 : OAI21X1 port map( A => n172, B => n999, C => n965, Y => n966);
   U1201 : OAI21X1 port map( A => n967, B => n966, C => n31, Y => n970);
   U1202 : NAND2X1 port map( A => n206, B => n1454, Y => n969);
   U1203 : NAND3X1 port map( A => n971, B => n970, C => n969, Y => n972);
   U1204 : NAND2X1 port map( A => n974, B => n972, Y => n979);
   U1205 : AND2X2 port map( A => currentPlainKey_45_port, B => n187, Y => n977)
                           ;
   U1206 : AOI21X1 port map( A => n209, B => n1455, C => n977, Y => n978);
   U1207 : NAND3X1 port map( A => n980, B => n979, C => n978, Y => n1646);
   U1208 : AOI22X1 port map( A => currentPlainKey_46_port, B => n187, C => n193
                           , D => n1454, Y => n996);
   U1209 : NAND2X1 port map( A => n181, B => n1453, Y => n992);
   U1210 : NAND2X1 port map( A => n20, B => n79, Y => n1010);
   U1211 : INVX2 port map( A => n1010, Y => n1079);
   U1212 : NAND2X1 port map( A => n1079, B => n1132, Y => n984);
   U1213 : NAND2X1 port map( A => n29, B => n153, Y => n1013);
   U1214 : INVX2 port map( A => n1013, Y => n981);
   U1215 : NAND2X1 port map( A => n1877, B => n981, Y => n983);
   U1216 : AOI21X1 port map( A => n984, B => n983, C => n982, Y => n986);
   U1217 : OAI22X1 port map( A => n156, B => n999, C => n1888, D => n168, Y => 
                           n985);
   U1218 : OAI21X1 port map( A => n986, B => n985, C => n31, Y => n991);
   U1219 : NAND2X1 port map( A => n1021, B => n205, Y => n987);
   U1221 : NAND3X1 port map( A => n992, B => n991, C => n987, Y => n994);
   U1222 : MUX2X1 port map( B => n994, A => n210, S => n993, Y => n995);
   U1223 : NAND2X1 port map( A => n996, B => n995, Y => n1647);
   U1224 : AOI22X1 port map( A => currentPlainKey_47_port, B => n187, C => n208
                           , D => n1454, Y => n1009);
   U1225 : NAND2X1 port map( A => n206, B => n1453, Y => n1003);
   U1226 : NOR2X1 port map( A => n1888, B => n161, Y => n998);
   U1227 : OAI22X1 port map( A => n71, B => n1010, C => n1880, D => n1013, Y =>
                           n997);
   U1228 : OAI21X1 port map( A => n998, B => n997, C => n1036, Y => n1001);
   U1229 : INVX2 port map( A => n999, Y => n1053);
   U1230 : NAND2X1 port map( A => n1053, B => n180, Y => n1000);
   U1231 : NAND3X1 port map( A => n1003, B => n1001, C => n1000, Y => n1005);
   U1232 : NAND2X1 port map( A => n31, B => n1005, Y => n1008);
   U1233 : NAND2X1 port map( A => n1021, B => n197, Y => n1007);
   U1234 : NAND3X1 port map( A => n1009, B => n1008, C => n1007, Y => n1648);
   U1235 : AOI22X1 port map( A => currentPlainKey_48_port, B => n185, C => n193
                           , D => n1453, Y => n1024);
   U1236 : NAND2X1 port map( A => n181, B => n1452, Y => n1020);
   U1237 : OAI22X1 port map( A => n156, B => n1010, C => n1896, D => n168, Y =>
                           n1015);
   U1238 : NAND2X1 port map( A => n79, B => n23, Y => n1059);
   U1239 : NAND2X1 port map( A => n1896, B => n1059, Y => n1043);
   U1240 : INVX2 port map( A => n1043, Y => n1093);
   U1241 : NAND2X1 port map( A => n1883, B => n1093, Y => n1012);
   U1242 : OAI22X1 port map( A => n135, B => n1059, C => n1013, D => n1012, Y 
                           => n1014);
   U1243 : OAI21X1 port map( A => n1015, B => n1014, C => n1036, Y => n1017);
   U1244 : NAND2X1 port map( A => n1053, B => n203, Y => n1016);
   U1245 : NAND3X1 port map( A => n1020, B => n1017, C => n1016, Y => n1022);
   U1246 : MUX2X1 port map( B => n1022, A => n210, S => n1021, Y => n1023);
   U1247 : NAND2X1 port map( A => n1024, B => n1023, Y => n1649);
   U1248 : NAND2X1 port map( A => n1053, B => n197, Y => n1041);
   U1249 : NAND2X1 port map( A => n1079, B => n180, Y => n1032);
   U1250 : NOR2X1 port map( A => n1896, B => n161, Y => n1028);
   U1251 : INVX2 port map( A => n1887, Y => n1025);
   U1252 : NAND3X1 port map( A => n1093, B => n153, C => n1025, Y => n1026);
   U1253 : OAI21X1 port map( A => n168, B => n1059, C => n1026, Y => n1027);
   U1254 : OAI21X1 port map( A => n1028, B => n1027, C => n29, Y => n1030);
   U1255 : NAND2X1 port map( A => n206, B => n1452, Y => n1029);
   U1256 : NAND3X1 port map( A => n1032, B => n1030, C => n1029, Y => n1035);
   U1257 : NAND2X1 port map( A => n1036, B => n1035, Y => n1040);
   U1258 : AND2X2 port map( A => currentPlainKey_49_port, B => n187, Y => n1037
                           );
   U1259 : AOI21X1 port map( A => n209, B => n1453, C => n1037, Y => n1039);
   U1260 : NAND3X1 port map( A => n1041, B => n1040, C => n1039, Y => n1650);
   U1261 : AOI22X1 port map( A => currentPlainKey_50_port, B => n186, C => n192
                           , D => n1452, Y => n1056);
   U1262 : NAND2X1 port map( A => n183, B => n1451, Y => n1052);
   U1263 : NAND2X1 port map( A => n5, B => n119, Y => n1069);
   U1264 : INVX2 port map( A => n1069, Y => n1140);
   U1265 : NAND2X1 port map( A => n1140, B => n1132, Y => n1045);
   U1266 : NAND2X1 port map( A => n51, B => n153, Y => n1071);
   U1267 : INVX2 port map( A => n1071, Y => n1042);
   U1268 : NAND2X1 port map( A => n1891, B => n1042, Y => n1044);
   U1269 : AOI21X1 port map( A => n1045, B => n1044, C => n1043, Y => n1049);
   U1270 : OAI22X1 port map( A => n158, B => n1059, C => n1903, D => n168, Y =>
                           n1048);
   U1271 : OAI21X1 port map( A => n1049, B => n1048, C => n29, Y => n1051);
   U1272 : NAND2X1 port map( A => n1079, B => n203, Y => n1050);
   U1275 : NAND3X1 port map( A => n1052, B => n1051, C => n1050, Y => n1054);
   U1276 : MUX2X1 port map( B => n1054, A => n210, S => n1053, Y => n1055);
   U1277 : NAND2X1 port map( A => n1056, B => n1055, Y => n1651);
   U1278 : AOI22X1 port map( A => currentPlainKey_51_port, B => n187, C => n208
                           , D => n1452, Y => n1068);
   U1279 : NAND2X1 port map( A => n207, B => n1451, Y => n1064);
   U1280 : NOR2X1 port map( A => n1903, B => n161, Y => n1058);
   U1281 : OAI22X1 port map( A => n173, B => n1069, C => n1895, D => n1071, Y 
                           => n1057);
   U1282 : OAI21X1 port map( A => n1058, B => n1057, C => n1093, Y => n1061);
   U1283 : INVX2 port map( A => n1059, Y => n1114);
   U1284 : NAND2X1 port map( A => n1114, B => n180, Y => n1060);
   U1285 : NAND3X1 port map( A => n1064, B => n1061, C => n1060, Y => n1065);
   U1286 : NAND2X1 port map( A => n29, B => n1065, Y => n1067);
   U1287 : NAND2X1 port map( A => n1079, B => n197, Y => n1066);
   U1288 : NAND3X1 port map( A => n1068, B => n1067, C => n1066, Y => n1652);
   U1289 : AOI22X1 port map( A => currentPlainKey_52_port, B => n187, C => n192
                           , D => n1451, Y => n1082);
   U1290 : NAND2X1 port map( A => n181, B => n1450, Y => n1076);
   U1291 : OAI22X1 port map( A => n156, B => n1069, C => n1910, D => n168, Y =>
                           n1073);
   U1292 : NAND2X1 port map( A => n5, B => n1477, Y => n1118);
   U1293 : NAND2X1 port map( A => n1910, B => n1118, Y => n1099);
   U1294 : INVX2 port map( A => n1099, Y => n1153);
   U1295 : NAND2X1 port map( A => n1898, B => n1153, Y => n1070);
   U1296 : OAI22X1 port map( A => n1118, B => n133, C => n1071, D => n1070, Y 
                           => n1072);
   U1297 : OAI21X1 port map( A => n1073, B => n1072, C => n1093, Y => n1075);
   U1298 : NAND2X1 port map( A => n1114, B => n203, Y => n1074);
   U1299 : NAND3X1 port map( A => n1076, B => n1075, C => n1074, Y => n1080);
   U1300 : MUX2X1 port map( B => n1080, A => n210, S => n1079, Y => n1081);
   U1301 : NAND2X1 port map( A => n1082, B => n1081, Y => n1653);
   U1302 : NAND2X1 port map( A => n1114, B => n197, Y => n1097);
   U1303 : NAND2X1 port map( A => n1140, B => n180, Y => n1091);
   U1304 : NOR2X1 port map( A => n1910, B => n161, Y => n1086);
   U1306 : INVX2 port map( A => n1902, Y => n1083);
   U1307 : NAND3X1 port map( A => n1153, B => n153, C => n1083, Y => n1084);
   U1308 : OAI21X1 port map( A => n173, B => n1118, C => n1084, Y => n1085);
   U1309 : OAI21X1 port map( A => n1086, B => n1085, C => n51, Y => n1088);
   U1310 : NAND2X1 port map( A => n206, B => n1450, Y => n1087);
   U1311 : NAND3X1 port map( A => n1091, B => n1088, C => n1087, Y => n1092);
   U1312 : NAND2X1 port map( A => n1093, B => n1092, Y => n1096);
   U1313 : AND2X2 port map( A => currentPlainKey_53_port, B => n187, Y => n1094
                           );
   U1316 : AOI21X1 port map( A => n209, B => n1451, C => n1094, Y => n1095);
   U1317 : NAND3X1 port map( A => n1097, B => n1096, C => n1095, Y => n1654);
   U1318 : AOI22X1 port map( A => currentPlainKey_54_port, B => n185, C => n192
                           , D => n1450, Y => n1117);
   U1319 : NAND2X1 port map( A => n181, B => n1449, Y => n1113);
   U1320 : NAND2X1 port map( A => n5, B => n1474, Y => n1121);
   U1321 : NAND2X1 port map( A => n1921, B => n1121, Y => n1134);
   U1322 : INVX2 port map( A => n1134, Y => n1174);
   U1323 : NAND3X1 port map( A => n1905, B => n153, C => n1174, Y => n1102);
   U1324 : INVX2 port map( A => n1121, Y => n1190);
   U1325 : NAND2X1 port map( A => n1132, B => n1190, Y => n1100);
   U1326 : AOI21X1 port map( A => n1102, B => n1100, C => n1099, Y => n1110);
   U1327 : OAI22X1 port map( A => n1921, B => n71, C => n156, D => n1118, Y => 
                           n1109);
   U1328 : OAI21X1 port map( A => n1110, B => n1109, C => n51, Y => n1112);
   U1329 : NAND2X1 port map( A => n1140, B => n203, Y => n1111);
   U1330 : NAND3X1 port map( A => n1113, B => n1112, C => n1111, Y => n1115);
   U1331 : MUX2X1 port map( B => n1115, A => n210, S => n1114, Y => n1116);
   U1332 : NAND2X1 port map( A => n1117, B => n1116, Y => n1655);
   U1333 : NAND2X1 port map( A => n1140, B => n197, Y => n1131);
   U1334 : INVX2 port map( A => n1118, Y => n1165);
   U1335 : NAND2X1 port map( A => n1165, B => n178, Y => n1126);
   U1336 : NOR2X1 port map( A => n1921, B => n161, Y => n1123);
   U1337 : INVX2 port map( A => n1909, Y => n1119);
   U1338 : NAND3X1 port map( A => n1174, B => n11, C => n1119, Y => n1120);
   U1339 : OAI21X1 port map( A => n1121, B => n71, C => n1120, Y => n1122);
   U1340 : OAI21X1 port map( A => n1123, B => n1122, C => n1153, Y => n1125);
   U1341 : NAND2X1 port map( A => n207, B => n1449, Y => n1124);
   U1342 : NAND3X1 port map( A => n1126, B => n1125, C => n1124, Y => n1127);
   U1343 : NAND2X1 port map( A => n51, B => n1127, Y => n1130);
   U1344 : AND2X2 port map( A => currentPlainKey_55_port, B => n187, Y => n1128
                           );
   U1345 : AOI21X1 port map( A => n209, B => n1450, C => n1128, Y => n1129);
   U1346 : NAND3X1 port map( A => n1131, B => n1130, C => n1129, Y => n1656);
   U1347 : AOI22X1 port map( A => currentPlainKey_56_port, B => n186, C => n192
                           , D => n1449, Y => n1145);
   U1348 : NAND2X1 port map( A => n181, B => n1448, Y => n1139);
   U1349 : NAND2X1 port map( A => n5, B => n7, Y => n1170);
   U1350 : NAND3X1 port map( A => n1098, B => n1170, C => n1931, Y => n1146);
   U1351 : INVX2 port map( A => n1146, Y => n1196);
   U1352 : INVX2 port map( A => n1170, Y => n1266);
   U1353 : AOI22X1 port map( A => n1915, B => n1196, C => n1132, D => n1266, Y 
                           => n1135);
   U1354 : AOI22X1 port map( A => n166, B => n1190, C => n175, D => n1447, Y =>
                           n1133);
   U1355 : OAI21X1 port map( A => n1135, B => n1134, C => n1133, Y => n1136);
   U1356 : NAND2X1 port map( A => n1153, B => n1136, Y => n1138);
   U1357 : NAND2X1 port map( A => n1165, B => n203, Y => n1137);
   U1358 : NAND3X1 port map( A => n1139, B => n1138, C => n1137, Y => n1141);
   U1359 : MUX2X1 port map( B => n1141, A => n210, S => n1140, Y => n1142);
   U1360 : NAND2X1 port map( A => n1145, B => n1142, Y => n1657);
   U1361 : AOI22X1 port map( A => currentPlainKey_57_port, B => n187, C => n208
                           , D => n1449, Y => n1156);
   U1362 : NAND2X1 port map( A => n207, B => n1448, Y => n1151);
   U1363 : NOR2X1 port map( A => n1920, B => n1146, Y => n1148);
   U1364 : OAI22X1 port map( A => n1931, B => n156, C => n1170, D => n168, Y =>
                           n1147);
   U1365 : OAI21X1 port map( A => n1148, B => n1147, C => n1174, Y => n1150);
   U1366 : NAND2X1 port map( A => n1190, B => n178, Y => n1149);
   U1367 : NAND3X1 port map( A => n1151, B => n1150, C => n1149, Y => n1152);
   U1368 : NAND2X1 port map( A => n1153, B => n1152, Y => n1155);
   U1369 : NAND2X1 port map( A => n1165, B => n197, Y => n1154);
   U1370 : NAND3X1 port map( A => n1156, B => n1155, C => n1154, Y => n1658);
   U1371 : AOI22X1 port map( A => currentPlainKey_58_port, B => n187, C => n192
                           , D => n1448, Y => n1168);
   U1372 : NAND2X1 port map( A => n181, B => n1447, Y => n1164);
   U1373 : NAND2X1 port map( A => n1196, B => n1969, Y => n1183);
   U1374 : INVX2 port map( A => n1925, Y => n1157);
   U1375 : NOR2X1 port map( A => n1183, B => n1157, Y => n1161);
   U1376 : OAI22X1 port map( A => n1969, B => n71, C => n1170, D => n156, Y => 
                           n1159);
   U1377 : OAI21X1 port map( A => n1161, B => n1159, C => n1174, Y => n1163);
   U1378 : NAND2X1 port map( A => n1190, B => n203, Y => n1162);
   U1379 : NAND3X1 port map( A => n1164, B => n1163, C => n1162, Y => n1166);
   U1380 : MUX2X1 port map( B => n1166, A => n210, S => n1165, Y => n1167);
   U1381 : NAND2X1 port map( A => n1168, B => n1167, Y => n1659);
   U1382 : AOI22X1 port map( A => currentPlainKey_59_port, B => n187, C => n208
                           , D => n1448, Y => n1180);
   U1383 : OAI22X1 port map( A => n1931, B => n1171, C => n1170, D => n1169, Y 
                           => n1176);
   U1384 : INVX2 port map( A => n1930, Y => n1173);
   U1385 : NAND3X1 port map( A => RCV_DATA(3), B => n1446, C => n1196, Y => 
                           n1172);
   U1386 : OAI21X1 port map( A => n1183, B => n1173, C => n1172, Y => n1175);
   U1387 : OAI21X1 port map( A => n1176, B => n1175, C => n1174, Y => n1179);
   U1388 : NAND2X1 port map( A => n1190, B => n197, Y => n1177);
   U1389 : NAND3X1 port map( A => n1180, B => n1179, C => n1177, Y => n1660);
   U1390 : AOI22X1 port map( A => currentPlainKey_60_port, B => n185, C => n192
                           , D => n1447, Y => n1193);
   U1391 : NAND2X1 port map( A => n183, B => n1446, Y => n1189);
   U1392 : AOI22X1 port map( A => n1493, B => RCV_DATA(3), C => n1445, D => 
                           RCV_DATA(2), Y => n1182);
   U1393 : OAI21X1 port map( A => n222, B => n1963, C => n1182, Y => n1185);
   U1394 : INVX2 port map( A => n1183, Y => n1184);
   U1395 : OAI21X1 port map( A => n55, B => n1185, C => n1184, Y => n1188);
   U1396 : NAND2X1 port map( A => n207, B => n1266, Y => n1187);
   U1397 : NAND3X1 port map( A => n1189, B => n1188, C => n1187, Y => n1191);
   U1398 : MUX2X1 port map( B => n1191, A => n210, S => n1190, Y => n1192);
   U1399 : NAND2X1 port map( A => n1193, B => n1192, Y => n1661);
   U1400 : AOI22X1 port map( A => currentPlainKey_61_port, B => n187, C => n208
                           , D => n1447, Y => n1263);
   U1401 : NAND2X1 port map( A => n1446, B => RCV_DATA(5), Y => n1194);
   U1402 : NAND2X1 port map( A => n1944, B => n1194, Y => n1195);
   U1403 : NAND2X1 port map( A => n1196, B => n1195, Y => n1262);
   U1404 : NAND2X1 port map( A => n1266, B => n197, Y => n1261);
   U1405 : NAND3X1 port map( A => n1263, B => n1262, C => n1261, Y => n1662);
   U1406 : AND2X2 port map( A => n187, B => currentPlainKey_62_port, Y => n1264
                           );
   U1407 : AOI21X1 port map( A => n195, B => n1446, C => n1264, Y => n1359);
   U1408 : NOR2X1 port map( A => n1446, B => n99, Y => n1265);
   U1409 : OAI21X1 port map( A => n1954, B => n1953, C => n1265, Y => n1268);
   U1410 : MUX2X1 port map( B => n1268, A => n1267, S => n1266, Y => n1357);
   U1411 : INVX2 port map( A => n1357, Y => n1358);
   U1412 : NAND2X1 port map( A => n1359, B => n1358, Y => n1663);
   U1413 : NAND2X1 port map( A => n186, B => currentPlainKey_63_port, Y => 
                           n1370);
   U1414 : NAND2X1 port map( A => n197, B => n1493, Y => n1366);
   U1415 : NOR2X1 port map( A => n1445, B => n99, Y => n1363);
   U1416 : INVX2 port map( A => n1968, Y => n1362);
   U1417 : OAI21X1 port map( A => n203, B => n1363, C => n1362, Y => n1365);
   U1418 : NAND2X1 port map( A => n1366, B => n1365, Y => n1368);
   U1419 : MUX2X1 port map( B => n1368, A => n217, S => n1446, Y => n1369);
   U1420 : NAND2X1 port map( A => n1370, B => n1369, Y => n1664);
   U1421 : NAND2X1 port map( A => n1371, B => n1414, Y => n1382);
   U1422 : INVX2 port map( A => n1382, Y => n1372);
   U1423 : NAND3X1 port map( A => n1372, B => n233, C => n1426, Y => n1380);
   U1424 : INVX2 port map( A => n1380, Y => n1378);
   U1425 : NAND2X1 port map( A => n1378, B => keyCount_3_port, Y => n1381);
   U1426 : NAND2X1 port map( A => address_0_port, B => n1380, Y => n1373);
   U1427 : NAND2X1 port map( A => n1381, B => n1373, Y => n1600);
   U1428 : NAND2X1 port map( A => address_1_port, B => n1380, Y => n1374);
   U1429 : NAND2X1 port map( A => n1381, B => n1374, Y => n1599);
   U1430 : NAND2X1 port map( A => address_2_port, B => n1380, Y => n1375);
   U1431 : NAND2X1 port map( A => n1381, B => n1375, Y => n1598);
   U1432 : MUX2X1 port map( B => address_3_port, A => keyCount_0_port, S => 
                           n1378, Y => n1376);
   U1433 : NAND2X1 port map( A => n1381, B => n1376, Y => n1597);
   U1434 : MUX2X1 port map( B => address_4_port, A => keyCount_1_port, S => 
                           n1378, Y => n1377);
   U1435 : NAND2X1 port map( A => n1381, B => n1377, Y => n1596);
   U1436 : MUX2X1 port map( B => address_5_port, A => keyCount_2_port, S => 
                           n1378, Y => n1379);
   U1437 : NAND2X1 port map( A => n1381, B => n1379, Y => n1595);
   U1438 : OAI21X1 port map( A => n1499, B => n1378, C => n1381, Y => n1594);
   U1439 : OAI21X1 port map( A => n1491, B => n1378, C => n1381, Y => n1593);
   U1440 : OAI21X1 port map( A => n1383, B => n1382, C => parityError, Y => 
                           n1386);
   U1441 : OAI21X1 port map( A => n2037, B => n2036, C => n1384, Y => n1385);
   U1442 : NAND2X1 port map( A => n1386, B => n1385, Y => nextParityError);
   U1443 : NOR2X1 port map( A => keyCount_0_port, B => n1438, Y => n1387);
   U1444 : NOR2X1 port map( A => n1387, B => n1442, Y => n1390);
   U1445 : INVX2 port map( A => n1444, Y => n1388);
   U1446 : NAND2X1 port map( A => keyCount_0_port, B => n1388, Y => n1389);
   U1447 : MUX2X1 port map( B => n1390, A => n1389, S => n1490, Y => n1583);
   U1448 : NAND2X1 port map( A => n1391, B => CLR_RBUFF_port, Y => n1405);
   U1449 : INVX2 port map( A => n1405, Y => n1400);
   U1450 : NAND2X1 port map( A => N1799, B => n1400, Y => n1392);
   U1451 : OAI21X1 port map( A => n1489, B => n1393, C => n1392, Y => n1592);
   U1452 : NAND2X1 port map( A => N1798, B => n1400, Y => n1394);
   U1453 : OAI21X1 port map( A => n1488, B => n1395, C => n1394, Y => n1591);
   U1454 : NAND2X1 port map( A => N1797, B => n1400, Y => n1396);
   U1455 : OAI21X1 port map( A => n1487, B => n1395, C => n1396, Y => n1590);
   U1456 : NAND2X1 port map( A => N1796, B => n1400, Y => n1397);
   U1457 : OAI21X1 port map( A => n1486, B => n1393, C => n1397, Y => n1589);
   U1458 : NAND2X1 port map( A => N1795, B => n1400, Y => n1398);
   U1459 : OAI21X1 port map( A => n1485, B => n1399, C => n1398, Y => n1588);
   U1460 : NAND2X1 port map( A => N1794, B => n1400, Y => n1401);
   U1461 : OAI21X1 port map( A => n1484, B => n1399, C => n1401, Y => n1587);
   U1462 : INVX2 port map( A => N1793, Y => n1402);
   U1463 : OAI22X1 port map( A => n1483, B => n1393, C => n1405, D => n1402, Y 
                           => n1586);
   U1464 : INVX2 port map( A => N1792, Y => n1404);
   U1465 : OAI22X1 port map( A => n1482, B => n1395, C => n1405, D => n1404, Y 
                           => n1585);
   U1466 : AOI21X1 port map( A => N694, B => RBUF_FULL, C => n1730, Y => n1407)
                           ;
   U1467 : NAND2X1 port map( A => n1407, B => n1406, Y => n1410);
   U1468 : NAND2X1 port map( A => n1408, B => n115, Y => n1409);
   U1469 : NAND2X1 port map( A => n1409, B => n1424, Y => n1431);
   U1470 : NAND2X1 port map( A => n1410, B => n1431, Y => n1421);
   U1471 : INVX2 port map( A => n1421, Y => n1412);
   U1472 : OAI21X1 port map( A => n1412, B => n115, C => n1411, Y => n1579);
   U1473 : AND2X2 port map( A => n1425, B => n1426, Y => n1418);
   U1474 : OAI21X1 port map( A => OE, B => SBE, C => n1406, Y => n1417);
   U1475 : OAI22X1 port map( A => RBUF_FULL, B => n1414, C => n1413, D => n1431
                           , Y => n1415);
   U1476 : AOI21X1 port map( A => n1420, B => n1433, C => n1415, Y => n1416);
   U1477 : NAND3X1 port map( A => n1418, B => n1417, C => n1416, Y => n1581);
   U1478 : AOI21X1 port map( A => state_1_port, B => n1421, C => n1420, Y => 
                           n1422);
   U1479 : NAND2X1 port map( A => n113, B => n1422, Y => n1582);
   U1480 : INVX2 port map( A => RBUF_FULL, Y => n1423);
   U1481 : AOI21X1 port map( A => n1425, B => n1424, C => n1423, Y => n1430);
   U1482 : NAND2X1 port map( A => n1570, B => n1576, Y => n1428);
   U1483 : OAI21X1 port map( A => n1428, B => n1427, C => n1426, Y => n1429);
   U1484 : NOR2X1 port map( A => n1430, B => n1429, Y => n1437);
   U1485 : INVX2 port map( A => n1731, Y => n1433);
   U1486 : OAI22X1 port map( A => n1438, B => n1433, C => n1432, D => n1431, Y 
                           => n1434);
   U1487 : NOR2X1 port map( A => n1435, B => n1434, Y => n1436);
   U1488 : NAND2X1 port map( A => n1437, B => n1436, Y => n1580);
   U1489 : NOR2X1 port map( A => keyCount_2_port, B => n1438, Y => n1440);
   U1490 : OAI21X1 port map( A => n1440, B => n1439, C => keyCount_3_port, Y =>
                           n1441);
   U1491 : OAI21X1 port map( A => n1731, B => n1444, C => n1441, Y => n1578);
   U1492 : NAND2X1 port map( A => n1442, B => keyCount_0_port, Y => n1443);
   U1493 : OAI21X1 port map( A => keyCount_0_port, B => n1444, C => n1443, Y =>
                           n1577);
   U1494 : INVX2 port map( A => keyCount_3_port, Y => N694);
   U1495 : INVX2 port map( A => keyCount_0_port, Y => n1479);
   U1496 : INVX2 port map( A => keyCount_2_port, Y => n1480);
   U1497 : INVX2 port map( A => parityAccumulator_0_port, Y => n1482);
   U1498 : INVX2 port map( A => parityAccumulator_1_port, Y => n1483);
   U1499 : INVX2 port map( A => parityAccumulator_2_port, Y => n1484);
   U1500 : INVX2 port map( A => parityAccumulator_3_port, Y => n1485);
   U1501 : INVX2 port map( A => parityAccumulator_4_port, Y => n1486);
   U1502 : INVX2 port map( A => parityAccumulator_5_port, Y => n1487);
   U1503 : INVX2 port map( A => parityAccumulator_6_port, Y => n1488);
   U1504 : INVX2 port map( A => parityAccumulator_7_port, Y => n1489);
   U1505 : INVX2 port map( A => keyCount_1_port, Y => n1490);
   U1506 : INVX2 port map( A => address_7_port, Y => n1491);
   U1507 : INVX2 port map( A => n1945, Y => n1492);
   U1508 : INVX2 port map( A => n1967, Y => n1493);
   U1509 : INVX2 port map( A => n1963, Y => n1494);
   U1510 : INVX2 port map( A => n1962, Y => n1495);
   U1511 : INVX2 port map( A => n1959, Y => n1496);
   U1512 : INVX2 port map( A => n1957, Y => n1497);
   U1513 : INVX2 port map( A => address_6_port, Y => n1499);
   U1514 : INVX2 port map( A => n1923, Y => n1500);
   U1515 : INVX2 port map( A => n1927, Y => n1501);
   U1516 : INVX2 port map( A => n1938, Y => n1502);
   U1517 : INVX2 port map( A => n1956, Y => n1503);
   U1518 : INVX2 port map( A => address_5_port, Y => n1504);
   U1519 : INVX2 port map( A => address_4_port, Y => n1505);
   U1520 : INVX2 port map( A => currentPlainKey_63_port, Y => n1506);
   U1521 : INVX2 port map( A => currentPlainKey_62_port, Y => n1507);
   U1522 : INVX2 port map( A => currentPlainKey_61_port, Y => n1508);
   U1523 : INVX2 port map( A => currentPlainKey_60_port, Y => n1509);
   U1524 : INVX2 port map( A => currentPlainKey_59_port, Y => n1510);
   U1525 : INVX2 port map( A => currentPlainKey_58_port, Y => n1511);
   U1526 : INVX2 port map( A => currentPlainKey_57_port, Y => n1512);
   U1527 : INVX2 port map( A => currentPlainKey_56_port, Y => n1513);
   U1528 : INVX2 port map( A => currentPlainKey_55_port, Y => n1514);
   U1529 : INVX2 port map( A => currentPlainKey_54_port, Y => n1515);
   U1530 : INVX2 port map( A => currentPlainKey_53_port, Y => n1516);
   U1531 : INVX2 port map( A => currentPlainKey_52_port, Y => n1517);
   U1532 : INVX2 port map( A => currentPlainKey_51_port, Y => n1518);
   U1533 : INVX2 port map( A => currentPlainKey_50_port, Y => n1519);
   U1534 : INVX2 port map( A => currentPlainKey_49_port, Y => n1520);
   U1535 : INVX2 port map( A => currentPlainKey_48_port, Y => n1521);
   U1536 : INVX2 port map( A => currentPlainKey_47_port, Y => n1522);
   U1537 : INVX2 port map( A => currentPlainKey_46_port, Y => n1523);
   U1538 : INVX2 port map( A => currentPlainKey_45_port, Y => n1524);
   U1539 : INVX2 port map( A => currentPlainKey_44_port, Y => n1525);
   U1540 : INVX2 port map( A => currentPlainKey_43_port, Y => n1526);
   U1541 : INVX2 port map( A => currentPlainKey_42_port, Y => n1527);
   U1542 : INVX2 port map( A => currentPlainKey_41_port, Y => n1528);
   U1543 : INVX2 port map( A => currentPlainKey_40_port, Y => n1529);
   U1544 : INVX2 port map( A => currentPlainKey_39_port, Y => n1530);
   U1545 : INVX2 port map( A => currentPlainKey_38_port, Y => n1531);
   U1546 : INVX2 port map( A => currentPlainKey_37_port, Y => n1532);
   U1547 : INVX2 port map( A => currentPlainKey_36_port, Y => n1533);
   U1548 : INVX2 port map( A => currentPlainKey_35_port, Y => n1534);
   U1549 : INVX2 port map( A => currentPlainKey_34_port, Y => n1535);
   U1550 : INVX2 port map( A => currentPlainKey_33_port, Y => n1536);
   U1551 : INVX2 port map( A => currentPlainKey_32_port, Y => n1537);
   U1552 : INVX2 port map( A => currentPlainKey_31_port, Y => n1538);
   U1553 : INVX2 port map( A => currentPlainKey_30_port, Y => n1539);
   U1554 : INVX2 port map( A => currentPlainKey_29_port, Y => n1540);
   U1555 : INVX2 port map( A => currentPlainKey_28_port, Y => n1541);
   U1556 : INVX2 port map( A => currentPlainKey_27_port, Y => n1542);
   U1557 : INVX2 port map( A => currentPlainKey_26_port, Y => n1543);
   U1558 : INVX2 port map( A => currentPlainKey_25_port, Y => n1544);
   U1559 : INVX2 port map( A => currentPlainKey_24_port, Y => n1545);
   U1560 : INVX2 port map( A => currentPlainKey_23_port, Y => n1546);
   U1561 : INVX2 port map( A => currentPlainKey_22_port, Y => n1547);
   U1562 : INVX2 port map( A => currentPlainKey_21_port, Y => n1548);
   U1563 : INVX2 port map( A => currentPlainKey_20_port, Y => n1549);
   U1564 : INVX2 port map( A => currentPlainKey_19_port, Y => n1550);
   U1565 : INVX2 port map( A => currentPlainKey_18_port, Y => n1551);
   U1566 : INVX2 port map( A => currentPlainKey_17_port, Y => n1552);
   U1567 : INVX2 port map( A => currentPlainKey_16_port, Y => n1553);
   U1568 : INVX2 port map( A => currentPlainKey_15_port, Y => n1554);
   U1569 : INVX2 port map( A => currentPlainKey_14_port, Y => n1555);
   U1570 : INVX2 port map( A => currentPlainKey_13_port, Y => n1556);
   U1571 : INVX2 port map( A => currentPlainKey_12_port, Y => n1557);
   U1572 : INVX2 port map( A => currentPlainKey_11_port, Y => n1558);
   U1573 : INVX2 port map( A => currentPlainKey_10_port, Y => n1559);
   U1574 : INVX2 port map( A => currentPlainKey_9_port, Y => n1560);
   U1575 : INVX2 port map( A => currentPlainKey_8_port, Y => n1561);
   U1576 : INVX2 port map( A => currentPlainKey_7_port, Y => n1562);
   U1577 : INVX2 port map( A => currentPlainKey_6_port, Y => n1563);
   U1578 : INVX2 port map( A => currentPlainKey_5_port, Y => n1564);
   U1579 : INVX2 port map( A => currentPlainKey_4_port, Y => n1565);
   U1580 : INVX2 port map( A => currentPlainKey_0_port, Y => n1569);
   U1581 : INVX2 port map( A => SBE, Y => n1570);
   U1582 : INVX2 port map( A => OE, Y => n1576);

end SYN_keyb;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_sr_10bit_0 is

   port( CLK, RST, SHIFT_STROBE, SERIAL_IN : in std_logic;  LOAD_DATA : out 
         std_logic_vector (7 downto 0);  STOP_DATA : out std_logic_vector (1 
         downto 0));

end uart_sr_10bit_0;

architecture SYN_dataflow of uart_sr_10bit_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal LOAD_DATA_7_port, LOAD_DATA_6_port, LOAD_DATA_5_port, 
      LOAD_DATA_4_port, LOAD_DATA_3_port, LOAD_DATA_2_port, LOAD_DATA_1_port, 
      LOAD_DATA_0_port, STOP_DATA_1_port, STOP_DATA_0_port, n1, n2, n4, n5, n6,
      n7, n8, n9, n10, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, 
      n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45 : 
      std_logic;

begin
   LOAD_DATA <= ( LOAD_DATA_7_port, LOAD_DATA_6_port, LOAD_DATA_5_port, 
      LOAD_DATA_4_port, LOAD_DATA_3_port, LOAD_DATA_2_port, LOAD_DATA_1_port, 
      LOAD_DATA_0_port );
   STOP_DATA <= ( STOP_DATA_1_port, STOP_DATA_0_port );
   
   U2 : OAI21X1 port map( A => n32, B => n13, C => n45, Y => n43);
   U3 : NAND2X1 port map( A => LOAD_DATA_0_port, B => n13, Y => n45);
   U4 : OAI22X1 port map( A => n13, B => n31, C => SHIFT_STROBE, D => n32, Y =>
                           n42);
   U6 : OAI22X1 port map( A => n13, B => n29, C => SHIFT_STROBE, D => n31, Y =>
                           n41);
   U8 : OAI22X1 port map( A => n13, B => n27, C => SHIFT_STROBE, D => n29, Y =>
                           n40);
   U10 : OAI22X1 port map( A => n13, B => n25, C => SHIFT_STROBE, D => n27, Y 
                           => n39);
   U12 : OAI22X1 port map( A => n13, B => n23, C => SHIFT_STROBE, D => n25, Y 
                           => n38);
   U14 : OAI22X1 port map( A => n13, B => n21, C => SHIFT_STROBE, D => n23, Y 
                           => n37);
   U16 : OAI22X1 port map( A => n13, B => n19, C => SHIFT_STROBE, D => n21, Y 
                           => n36);
   U18 : OAI22X1 port map( A => n13, B => n17, C => SHIFT_STROBE, D => n19, Y 
                           => n35);
   U22 : OAI21X1 port map( A => SHIFT_STROBE, B => n17, C => n44, Y => n34);
   U23 : NAND2X1 port map( A => SERIAL_IN, B => SHIFT_STROBE, Y => n44);
   present_val_reg_9_inst : DFFSR port map( D => n34, CLK => CLK, R => n15, S 
                           => n11, Q => STOP_DATA_1_port);
   present_val_reg_8_inst : DFFSR port map( D => n35, CLK => CLK, R => n15, S 
                           => n10, Q => STOP_DATA_0_port);
   present_val_reg_7_inst : DFFSR port map( D => n36, CLK => CLK, R => n15, S 
                           => n9, Q => LOAD_DATA_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n37, CLK => CLK, R => n15, S 
                           => n8, Q => LOAD_DATA_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n38, CLK => CLK, R => n15, S 
                           => n7, Q => LOAD_DATA_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n39, CLK => CLK, R => n15, S 
                           => n6, Q => LOAD_DATA_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n40, CLK => CLK, R => n15, S 
                           => n5, Q => LOAD_DATA_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n41, CLK => CLK, R => n15, S 
                           => n4, Q => LOAD_DATA_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n42, CLK => CLK, R => n15, S 
                           => n2, Q => LOAD_DATA_1_port);
   present_val_reg_0_inst : DFFSR port map( D => n43, CLK => CLK, R => n15, S 
                           => n1, Q => LOAD_DATA_0_port);
   n1 <= '1';
   n2 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   U24 : INVX2 port map( A => RST, Y => n15);
   U25 : INVX2 port map( A => SHIFT_STROBE, Y => n13);
   U26 : INVX2 port map( A => STOP_DATA_1_port, Y => n17);
   U27 : INVX2 port map( A => STOP_DATA_0_port, Y => n19);
   U28 : INVX2 port map( A => LOAD_DATA_7_port, Y => n21);
   U29 : INVX2 port map( A => LOAD_DATA_6_port, Y => n23);
   U30 : INVX2 port map( A => LOAD_DATA_5_port, Y => n25);
   U31 : INVX2 port map( A => LOAD_DATA_4_port, Y => n27);
   U32 : INVX2 port map( A => LOAD_DATA_3_port, Y => n29);
   U33 : INVX2 port map( A => LOAD_DATA_2_port, Y => n31);
   U34 : INVX2 port map( A => LOAD_DATA_1_port, Y => n32);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_sb_check_0 is

   port( RST, CLK, SBC_CLR, SBC_EN : in std_logic;  STOP_DATA : in 
         std_logic_vector (1 downto 0);  SB_DETECT, SBE : out std_logic);

end uart_sb_check_0;

architecture SYN_behavioral of uart_sb_check_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal SBE_prime, sb_detect_flag, n1, n2, n3, n4, n5, n6, n10, n11, n12 : 
      std_logic;

begin
   
   U6 : OR2X2 port map( A => SBC_CLR, B => STOP_DATA(0), Y => n12);
   U10 : NOR2X1 port map( A => n12, B => n11, Y => sb_detect_flag);
   U11 : NAND2X1 port map( A => STOP_DATA(1), B => SBC_EN, Y => n11);
   U12 : NOR2X1 port map( A => n6, B => n10, Y => SBE_prime);
   U13 : OAI21X1 port map( A => STOP_DATA(0), B => n4, C => n5, Y => n10);
   SBE_reg : DFFSR port map( D => SBE_prime, CLK => CLK, R => n3, S => n2, Q =>
                           SBE);
   SB_DETECT_reg : DFFSR port map( D => sb_detect_flag, CLK => CLK, R => n3, S 
                           => n1, Q => SB_DETECT);
   n1 <= '1';
   n2 <= '1';
   U5 : INVX2 port map( A => RST, Y => n3);
   U7 : INVX2 port map( A => STOP_DATA(1), Y => n4);
   U8 : INVX2 port map( A => SBC_CLR, Y => n5);
   U9 : INVX2 port map( A => SBC_EN, Y => n6);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_buf_full_0 is

   port( CLK, RST, CLR_RBUF, SET_RBUF_FULL : in std_logic;  RBUF_FULL : out 
         std_logic);

end uart_rcv_buf_full_0;

architecture SYN_Behavioral of uart_rcv_buf_full_0 is

   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal RBUF_FULL_port, n2, n4, n5 : std_logic;

begin
   RBUF_FULL <= RBUF_FULL_port;
   
   U3 : NOR2X1 port map( A => RST, B => CLR_RBUF, Y => n5);
   U4 : OR2X2 port map( A => RBUF_FULL_port, B => SET_RBUF_FULL, Y => n4);
   Q_int_reg : DFFSR port map( D => n4, CLK => CLK, R => n5, S => n2, Q => 
                           RBUF_FULL_port);
   n2 <= '1';

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_buf_0 is

   port( CLK, RST, LOAD_RBUF : in std_logic;  LOAD_DATA : in std_logic_vector 
         (7 downto 0);  RCV_DATA : out std_logic_vector (7 downto 0));

end uart_rcv_buf_0;

architecture SYN_Behavioral of uart_rcv_buf_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, n2, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35 : std_logic;

begin
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   U3 : AOI22X1 port map( A => n17, B => LOAD_DATA(0), C => RCV_DATA_0_port, D 
                           => n27, Y => n35);
   U5 : AOI22X1 port map( A => LOAD_DATA(1), B => n17, C => RCV_DATA_1_port, D 
                           => n27, Y => n34);
   U7 : AOI22X1 port map( A => LOAD_DATA(2), B => n17, C => RCV_DATA_2_port, D 
                           => n27, Y => n33);
   U9 : AOI22X1 port map( A => LOAD_DATA(3), B => n17, C => RCV_DATA_3_port, D 
                           => n27, Y => n32);
   U11 : AOI22X1 port map( A => LOAD_DATA(4), B => n17, C => RCV_DATA_4_port, D
                           => n27, Y => n31);
   U13 : AOI22X1 port map( A => LOAD_DATA(5), B => n17, C => RCV_DATA_5_port, D
                           => n27, Y => n30);
   U15 : AOI22X1 port map( A => LOAD_DATA(6), B => n17, C => RCV_DATA_6_port, D
                           => n27, Y => n29);
   U18 : AOI22X1 port map( A => LOAD_DATA(7), B => n17, C => RCV_DATA_7_port, D
                           => n27, Y => n28);
   Q_int_reg_0_inst : DFFSR port map( D => n26, CLK => CLK, R => n18, S => n16,
                           Q => RCV_DATA_0_port);
   Q_int_reg_7_inst : DFFSR port map( D => n19, CLK => CLK, R => n18, S => n15,
                           Q => RCV_DATA_7_port);
   Q_int_reg_6_inst : DFFSR port map( D => n20, CLK => CLK, R => n18, S => n14,
                           Q => RCV_DATA_6_port);
   Q_int_reg_5_inst : DFFSR port map( D => n21, CLK => CLK, R => n18, S => n13,
                           Q => RCV_DATA_5_port);
   Q_int_reg_4_inst : DFFSR port map( D => n22, CLK => CLK, R => n18, S => n12,
                           Q => RCV_DATA_4_port);
   Q_int_reg_1_inst : DFFSR port map( D => n25, CLK => CLK, R => n18, S => n11,
                           Q => RCV_DATA_1_port);
   Q_int_reg_2_inst : DFFSR port map( D => n24, CLK => CLK, R => n18, S => n10,
                           Q => RCV_DATA_2_port);
   Q_int_reg_3_inst : DFFSR port map( D => n23, CLK => CLK, R => n18, S => n2, 
                           Q => RCV_DATA_3_port);
   n2 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   U17 : INVX2 port map( A => RST, Y => n18);
   U19 : BUFX2 port map( A => LOAD_RBUF, Y => n17);
   U20 : INVX2 port map( A => n28, Y => n19);
   U21 : INVX2 port map( A => n29, Y => n20);
   U22 : INVX2 port map( A => n30, Y => n21);
   U23 : INVX2 port map( A => n31, Y => n22);
   U24 : INVX2 port map( A => n32, Y => n23);
   U25 : INVX2 port map( A => n33, Y => n24);
   U26 : INVX2 port map( A => n34, Y => n25);
   U27 : INVX2 port map( A => n35, Y => n26);
   U28 : INVX2 port map( A => n17, Y => n27);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcu_0 is

   port( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT : in std_logic;  RBUF_LOAD
         , TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR : out 
         std_logic);

end uart_rcu_0;

architecture SYN_rcub of uart_rcu_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal RBUF_LOAD_port, TIMER_TRIG_port, CHK_ERROR_port, SET_RBUF_FULL_port, 
      SBC_EN_port, SBC_CLR_port, state_2_port, state_1_port, state_0_port, 
      timerRunning, count_7_port, count_6_port, count_5_port, count_4_port, 
      count_3_port, count_2_port, count_1_port, count_0_port, nextCount_7_port,
      nextCount_6_port, nextCount_5_port, nextCount_4_port, nextCount_3_port, 
      nextCount_2_port, nextCount_1_port, nextCount_0_port, nextState_1_port, 
      nextState_0_port, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, 
      N35, N36, N37, N38, N99, add_46_carry_3_port, add_46_carry_4_port, 
      add_46_carry_5_port, add_46_carry_6_port, add_46_carry_7_port, n1, n2, n3
      , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n22, n23, n24_port, n25_port, n26_port, n27_port, n28_port, 
      n29_port, n30_port, n31_port, n32_port, n33_port, n34_port, n35_port, 
      n36_port, n37_port, n38_port, n39, n40, n41, n42, n43, n44, n45, n46, n47
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99_port, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114 : std_logic;

begin
   RBUF_LOAD <= RBUF_LOAD_port;
   TIMER_TRIG <= TIMER_TRIG_port;
   CHK_ERROR <= CHK_ERROR_port;
   SET_RBUF_FULL <= SET_RBUF_FULL_port;
   SBC_EN <= SBC_EN_port;
   SBC_CLR <= SBC_CLR_port;
   
   nextCount_reg_0_inst : DFFSR port map( D => N31, CLK => CLK, R => n114, S =>
                           n27_port, Q => nextCount_0_port);
   n114 <= '1';
   U33 : AND2X2 port map( A => N30, B => timerRunning, Y => N38);
   U34 : AND2X2 port map( A => N29, B => timerRunning, Y => N37);
   U35 : AND2X2 port map( A => N28, B => timerRunning, Y => N36);
   U36 : AND2X2 port map( A => N27, B => timerRunning, Y => N35);
   U37 : AND2X2 port map( A => N26, B => timerRunning, Y => N34);
   U38 : AND2X2 port map( A => N25, B => timerRunning, Y => N33);
   U39 : AND2X2 port map( A => N24, B => timerRunning, Y => N32);
   U54 : OAI21X1 port map( A => n112, B => n43, C => n111, Y => n113);
   U55 : OAI21X1 port map( A => n44, B => n42, C => n43, Y => n111);
   U56 : NAND2X1 port map( A => n110, B => n109, Y => n87);
   U57 : OAI21X1 port map( A => n108, B => n107, C => timerRunning, Y => n109);
   U58 : NAND2X1 port map( A => n106, B => n105, Y => n107);
   U59 : NAND2X1 port map( A => n104, B => n105, Y => n86);
   U60 : NAND3X1 port map( A => n35_port, B => n110, C => CHK_ERROR_port, Y => 
                           n104);
   U61 : OAI21X1 port map( A => n103, B => n47, C => n102, Y => n85);
   U62 : NAND2X1 port map( A => n105, B => n101, Y => n103);
   U63 : NAND2X1 port map( A => n100, B => n38_port, Y => n105);
   U64 : NAND3X1 port map( A => n99_port, B => n98, C => n97, Y => n84);
   U65 : NAND3X1 port map( A => n34_port, B => n110, C => SET_RBUF_FULL_port, Y
                           => n97);
   U66 : NAND2X1 port map( A => n101, B => n98, Y => n108);
   U67 : NAND3X1 port map( A => nextState_0_port, B => nextState_1_port, C => 
                           n100, Y => n98);
   U68 : NAND3X1 port map( A => n36_port, B => n38_port, C => n100, Y => 
                           n99_port);
   U69 : OAI21X1 port map( A => n96, B => n45, C => n110, Y => n83);
   U70 : OAI21X1 port map( A => n96, B => n46, C => n110, Y => n82);
   U71 : NAND2X1 port map( A => n101, B => n102, Y => n96);
   U72 : NAND3X1 port map( A => nextState_1_port, B => n36_port, C => n39, Y =>
                           n102);
   U73 : NAND2X1 port map( A => n95, B => n106, Y => n81);
   U74 : NAND3X1 port map( A => nextState_1_port, B => n36_port, C => n100, Y 
                           => n106);
   U75 : NAND3X1 port map( A => n101, B => n110, C => RBUF_LOAD_port, Y => n95)
                           ;
   U76 : NAND3X1 port map( A => nextState_0_port, B => n38_port, C => n39, Y =>
                           n110);
   U77 : NAND3X1 port map( A => n36_port, B => n38_port, C => n39, Y => n101);
   U78 : OAI21X1 port map( A => n40, B => n43, C => n94, Y => n100);
   U79 : NAND3X1 port map( A => state_0_port, B => n43, C => state_1_port, Y =>
                           n94);
   U80 : NAND2X1 port map( A => n93, B => n92, Y => n112);
   U81 : OAI21X1 port map( A => n91, B => n92, C => n93, Y => nextState_1_port)
                           ;
   U82 : NOR2X1 port map( A => N99, B => state_2_port, Y => n91);
   U83 : OAI21X1 port map( A => state_2_port, B => n90, C => n93, Y => 
                           nextState_0_port);
   U84 : NAND2X1 port map( A => state_1_port, B => n44, Y => n93);
   U85 : AOI21X1 port map( A => START_BIT, B => n44, C => n89, Y => n90);
   U86 : OAI21X1 port map( A => N99, B => n92, C => n88, Y => n89);
   U87 : NAND2X1 port map( A => SB_DETECT, B => state_1_port, Y => n88);
   U88 : NAND2X1 port map( A => state_0_port, B => n42, Y => n92);
   U89 : NAND2X1 port map( A => n37_port, B => timerRunning, Y => N31);
   count_reg_7_inst : DFFSR port map( D => nextCount_7_port, CLK => CLK, R => 
                           n27_port, S => n26_port, Q => count_7_port);
   count_reg_6_inst : DFFSR port map( D => nextCount_6_port, CLK => CLK, R => 
                           n27_port, S => n25_port, Q => count_6_port);
   count_reg_5_inst : DFFSR port map( D => nextCount_5_port, CLK => CLK, R => 
                           n27_port, S => n24_port, Q => count_5_port);
   count_reg_4_inst : DFFSR port map( D => nextCount_4_port, CLK => CLK, R => 
                           n27_port, S => n23, Q => count_4_port);
   count_reg_3_inst : DFFSR port map( D => nextCount_3_port, CLK => CLK, R => 
                           n27_port, S => n22, Q => count_3_port);
   count_reg_2_inst : DFFSR port map( D => nextCount_2_port, CLK => CLK, R => 
                           n27_port, S => n20, Q => count_2_port);
   count_reg_1_inst : DFFSR port map( D => nextCount_1_port, CLK => CLK, R => 
                           n27_port, S => n19, Q => count_1_port);
   count_reg_0_inst : DFFSR port map( D => nextCount_0_port, CLK => CLK, R => 
                           n27_port, S => n18, Q => count_0_port);
   nextCount_reg_2_inst : DFFSR port map( D => N33, CLK => CLK, R => n27_port, 
                           S => n17, Q => nextCount_2_port);
   nextCount_reg_1_inst : DFFSR port map( D => N32, CLK => CLK, R => n27_port, 
                           S => n16, Q => nextCount_1_port);
   state_reg_2_inst : DFFSR port map( D => n41, CLK => CLK, R => n27_port, S =>
                           n15, Q => state_2_port);
   nextCount_reg_3_inst : DFFSR port map( D => N34, CLK => CLK, R => n27_port, 
                           S => n14, Q => nextCount_3_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n27_port, S => n13, Q => state_1_port);
   nextCount_reg_4_inst : DFFSR port map( D => N35, CLK => CLK, R => n27_port, 
                           S => n12, Q => nextCount_4_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n27_port, S => n11, Q => state_0_port);
   nextCount_reg_5_inst : DFFSR port map( D => N36, CLK => CLK, R => n27_port, 
                           S => n10, Q => nextCount_5_port);
   nextCount_reg_6_inst : DFFSR port map( D => N37, CLK => CLK, R => n27_port, 
                           S => n9, Q => nextCount_6_port);
   RBUF_LOAD_reg : DFFSR port map( D => n81, CLK => CLK, R => n27_port, S => n8
                           , Q => RBUF_LOAD_port);
   timerRunning_reg : DFFSR port map( D => n87, CLK => CLK, R => n27_port, S =>
                           n7, Q => timerRunning);
   TIMER_TRIG_reg : DFFSR port map( D => n82, CLK => CLK, R => n27_port, S => 
                           n6, Q => TIMER_TRIG_port);
   SBC_CLR_reg : DFFSR port map( D => n83, CLK => CLK, R => n27_port, S => n5, 
                           Q => SBC_CLR_port);
   SBC_EN_reg : DFFSR port map( D => n85, CLK => CLK, R => n27_port, S => n4, Q
                           => SBC_EN_port);
   nextCount_reg_7_inst : DFFSR port map( D => N38, CLK => CLK, R => n27_port, 
                           S => n3, Q => nextCount_7_port);
   SET_RBUF_FULL_reg : DFFSR port map( D => n84, CLK => CLK, R => n27_port, S 
                           => n2, Q => SET_RBUF_FULL_port);
   CHK_ERROR_reg : DFFSR port map( D => n86, CLK => CLK, R => n27_port, S => n1
                           , Q => CHK_ERROR_port);
   U3 : INVX4 port map( A => RST, Y => n27_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   n18 <= '1';
   n19 <= '1';
   n20 <= '1';
   n22 <= '1';
   n23 <= '1';
   n24_port <= '1';
   n25_port <= '1';
   n26_port <= '1';
   U30 : XOR2X1 port map( A => count_7_port, B => add_46_carry_7_port, Y => N30
                           );
   U31 : AND2X1 port map( A => count_6_port, B => add_46_carry_6_port, Y => 
                           add_46_carry_7_port);
   U32 : XOR2X1 port map( A => add_46_carry_6_port, B => count_6_port, Y => N29
                           );
   U40 : AND2X1 port map( A => count_5_port, B => add_46_carry_5_port, Y => 
                           add_46_carry_6_port);
   U41 : XOR2X1 port map( A => add_46_carry_5_port, B => count_5_port, Y => N28
                           );
   U42 : AND2X1 port map( A => count_4_port, B => add_46_carry_4_port, Y => 
                           add_46_carry_5_port);
   U43 : XOR2X1 port map( A => add_46_carry_4_port, B => count_4_port, Y => N27
                           );
   U44 : AND2X1 port map( A => count_3_port, B => add_46_carry_3_port, Y => 
                           add_46_carry_4_port);
   U45 : XOR2X1 port map( A => add_46_carry_3_port, B => count_3_port, Y => N26
                           );
   U46 : AND2X1 port map( A => count_2_port, B => count_1_port, Y => 
                           add_46_carry_3_port);
   U47 : XOR2X1 port map( A => count_1_port, B => count_2_port, Y => N25);
   U48 : INVX2 port map( A => count_1_port, Y => N24);
   U49 : OAI21X1 port map( A => count_0_port, B => count_1_port, C => 
                           count_2_port, Y => n28_port);
   U50 : NOR2X1 port map( A => n33_port, B => n28_port, Y => n29_port);
   U51 : OAI21X1 port map( A => n29_port, B => count_4_port, C => count_6_port,
                           Y => n30_port);
   U52 : OAI21X1 port map( A => n32_port, B => n30_port, C => n31_port, Y => 
                           N99);
   U53 : INVX2 port map( A => count_7_port, Y => n31_port);
   U90 : INVX2 port map( A => count_5_port, Y => n32_port);
   U91 : INVX2 port map( A => count_3_port, Y => n33_port);
   U92 : INVX2 port map( A => n108, Y => n34_port);
   U93 : INVX2 port map( A => n103, Y => n35_port);
   U94 : INVX2 port map( A => nextState_0_port, Y => n36_port);
   U95 : INVX2 port map( A => count_0_port, Y => n37_port);
   U96 : INVX2 port map( A => nextState_1_port, Y => n38_port);
   U97 : INVX2 port map( A => n100, Y => n39);
   U98 : INVX2 port map( A => n112, Y => n40);
   U99 : INVX2 port map( A => n113, Y => n41);
   U100 : INVX2 port map( A => state_1_port, Y => n42);
   U101 : INVX2 port map( A => state_2_port, Y => n43);
   U102 : INVX2 port map( A => state_0_port, Y => n44);
   U103 : INVX2 port map( A => SBC_CLR_port, Y => n45);
   U104 : INVX2 port map( A => TIMER_TRIG_port, Y => n46);
   U105 : INVX2 port map( A => SBC_EN_port, Y => n47);

end SYN_rcub;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_error_0 is

   port( RST, CLK, RBUF_FULL, CHK_ERROR : in std_logic;  OE : out std_logic);

end uart_error_0;

architecture SYN_behavioral of uart_error_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal OE_prime, n1, n2 : std_logic;

begin
   
   U5 : AND2X2 port map( A => RBUF_FULL, B => CHK_ERROR, Y => OE_prime);
   OE_reg : DFFSR port map( D => OE_prime, CLK => CLK, R => n2, S => n1, Q => 
                           OE);
   n1 <= '1';
   U4 : INVX2 port map( A => RST, Y => n2);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_edge_detector_0 is

   port( CLK, RST, SERIAL_IN : in std_logic;  START_BIT : out std_logic);

end uart_edge_detector_0;

architecture SYN_Behavioral of uart_edge_detector_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal Q_int, Q_int2, n1, n2, n4, n5 : std_logic;

begin
   
   Q_int_reg : DFFSR port map( D => SERIAL_IN, CLK => CLK, R => n2, S => n5, Q 
                           => Q_int);
   n5 <= '1';
   U7 : NOR2X1 port map( A => Q_int, B => n4, Y => START_BIT);
   Q_int2_reg : DFFSR port map( D => Q_int, CLK => CLK, R => n2, S => n1, Q => 
                           Q_int2);
   n1 <= '1';
   U4 : INVX2 port map( A => RST, Y => n2);
   U6 : INVX2 port map( A => Q_int2, Y => n4);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_timer_0 is

   port( CLK, RST, SENDING : in std_logic;  SHIFT_ENABLE_R, SHIFT_ENABLE_E : 
         out std_logic);

end tx_timer_0;

architecture SYN_moore of tx_timer_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_3_port, count_2_port, count_1_port, count_0_port, state, 
      nextcount_3_port, nextcount_2_port, nextcount_1_port, nextcount_0_port, 
      nxt_SHIFT_ENABLE_E, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n20, 
      n21, n22, n23, n24, n25, n26, n27 : std_logic;

begin
   SHIFT_ENABLE_R <= nxt_SHIFT_ENABLE_E;
   
   U14 : NOR2X1 port map( A => n27, B => n26, Y => nextcount_3_port);
   U15 : XNOR2X1 port map( A => count_3_port, B => n25, Y => n27);
   U16 : NOR2X1 port map( A => n24, B => n9, Y => n25);
   U17 : AOI21X1 port map( A => n23, B => state, C => n11, Y => 
                           nextcount_2_port);
   U18 : XNOR2X1 port map( A => n24, B => n9, Y => n23);
   U19 : NAND2X1 port map( A => count_1_port, B => count_0_port, Y => n24);
   U20 : NOR2X1 port map( A => n22, B => n26, Y => nextcount_1_port);
   U21 : NAND3X1 port map( A => SENDING, B => n21, C => state, Y => n26);
   U22 : XNOR2X1 port map( A => count_0_port, B => count_1_port, Y => n22);
   U23 : OAI21X1 port map( A => count_0_port, B => n11, C => state, Y => 
                           nextcount_0_port);
   U24 : NOR2X1 port map( A => n21, B => n20, Y => nxt_SHIFT_ENABLE_E);
   U25 : NAND3X1 port map( A => count_3_port, B => SENDING, C => state, Y => 
                           n20);
   U26 : NAND3X1 port map( A => n10, B => n9, C => n8, Y => n21);
   state_reg : DFFSR port map( D => SENDING, CLK => CLK, R => n7, S => n6, Q =>
                           state);
   count_reg_2_inst : DFFSR port map( D => nextcount_2_port, CLK => CLK, R => 
                           n7, S => n5, Q => count_2_port);
   count_reg_0_inst : DFFSR port map( D => nextcount_0_port, CLK => CLK, R => 
                           n7, S => n4, Q => count_0_port);
   count_reg_3_inst : DFFSR port map( D => nextcount_3_port, CLK => CLK, R => 
                           n7, S => n3, Q => count_3_port);
   count_reg_1_inst : DFFSR port map( D => nextcount_1_port, CLK => CLK, R => 
                           n7, S => n2, Q => count_1_port);
   SHIFT_ENABLE_E_reg : DFFSR port map( D => nxt_SHIFT_ENABLE_E, CLK => CLK, R 
                           => n7, S => n1, Q => SHIFT_ENABLE_E);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   U9 : INVX2 port map( A => RST, Y => n7);
   U10 : INVX2 port map( A => count_0_port, Y => n8);
   U11 : INVX2 port map( A => count_2_port, Y => n9);
   U12 : INVX2 port map( A => count_1_port, Y => n10);
   U13 : INVX2 port map( A => SENDING, Y => n11);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_tcu_0 is

   port( clk, rst, p_ready, t_bitstuff : in std_logic;  PRGA_OUT : in 
         std_logic_vector (7 downto 0);  prga_opcode : in std_logic_vector (1 
         downto 0);  t_crc : in std_logic_vector (15 downto 0);  sending, EOP, 
         next_byte : out std_logic;  send_data : out std_logic_vector (7 downto
         0);  t_strobe : out std_logic);

end tx_tcu_0;

architecture SYN_behavioral of tx_tcu_0 is

   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component tx_tcu_0_DW01_inc_0
      port( A : in std_logic_vector (6 downto 0);  SUM : out std_logic_vector 
            (6 downto 0));
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal send_data_7_port, send_data_6_port, send_data_5_port, 
      send_data_4_port, send_data_3_port, send_data_2_port, send_data_1_port, 
      send_data_0_port, state_2_port, state_1_port, state_0_port, count_5_port,
      count_4_port, count_3_port, count_2_port, count_1_port, count_0_port, 
      nextstate_2_port, nextstate_1_port, nextstate_0_port, flop_data_7_port, 
      flop_data_6_port, flop_data_5_port, flop_data_4_port, flop_data_3_port, 
      flop_data_2_port, flop_data_1_port, flop_data_0_port, 
      current_send_data_7_port, current_send_data_6_port, 
      current_send_data_5_port, current_send_data_4_port, 
      current_send_data_3_port, current_send_data_2_port, 
      current_send_data_1_port, current_send_data_0_port, N59, N60, N61, N62, 
      N63, N64, N65, N84, N85, N86, N87, N88, N89, N90, N188, r81_carry_1_port,
      r81_carry_2_port, r81_carry_3_port, r81_carry_4_port, r81_carry_5_port, 
      r81_carry_6_port, r81_B_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59_port, n60_port, n61_port, n62_port, n63_port, 
      n64_port, n65_port, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83, n84_port, n85_port, n86_port, 
      n87_port, n88_port, n89_port, n90_port, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188_port, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198 : std_logic;

begin
   send_data <= ( send_data_7_port, send_data_6_port, send_data_5_port, 
      send_data_4_port, send_data_3_port, send_data_2_port, send_data_1_port, 
      send_data_0_port );
   
   flop_data_reg_7_inst : DFFPOSX1 port map( D => n152, CLK => clk, Q => 
                           flop_data_7_port);
   current_send_data_reg_7_inst : DFFPOSX1 port map( D => n183, CLK => clk, Q 
                           => current_send_data_7_port);
   flop_data_reg_6_inst : DFFPOSX1 port map( D => n153, CLK => clk, Q => 
                           flop_data_6_port);
   current_send_data_reg_6_inst : DFFPOSX1 port map( D => n184, CLK => clk, Q 
                           => current_send_data_6_port);
   flop_data_reg_5_inst : DFFPOSX1 port map( D => n154, CLK => clk, Q => 
                           flop_data_5_port);
   current_send_data_reg_5_inst : DFFPOSX1 port map( D => n185, CLK => clk, Q 
                           => current_send_data_5_port);
   flop_data_reg_4_inst : DFFPOSX1 port map( D => n155, CLK => clk, Q => 
                           flop_data_4_port);
   current_send_data_reg_4_inst : DFFPOSX1 port map( D => n186, CLK => clk, Q 
                           => current_send_data_4_port);
   flop_data_reg_3_inst : DFFPOSX1 port map( D => n156, CLK => clk, Q => 
                           flop_data_3_port);
   current_send_data_reg_3_inst : DFFPOSX1 port map( D => n187, CLK => clk, Q 
                           => current_send_data_3_port);
   flop_data_reg_2_inst : DFFPOSX1 port map( D => n157, CLK => clk, Q => 
                           flop_data_2_port);
   current_send_data_reg_2_inst : DFFPOSX1 port map( D => n188_port, CLK => clk
                           , Q => current_send_data_2_port);
   flop_data_reg_1_inst : DFFPOSX1 port map( D => n174, CLK => clk, Q => 
                           flop_data_1_port);
   current_send_data_reg_1_inst : DFFPOSX1 port map( D => n189, CLK => clk, Q 
                           => current_send_data_1_port);
   flop_data_reg_0_inst : DFFPOSX1 port map( D => n175, CLK => clk, Q => 
                           flop_data_0_port);
   current_send_data_reg_0_inst : DFFPOSX1 port map( D => n190, CLK => clk, Q 
                           => current_send_data_0_port);
   send_data_reg_7_inst : DFFPOSX1 port map( D => n191, CLK => clk, Q => 
                           send_data_7_port);
   send_data_reg_6_inst : DFFPOSX1 port map( D => n192, CLK => clk, Q => 
                           send_data_6_port);
   send_data_reg_5_inst : DFFPOSX1 port map( D => n193, CLK => clk, Q => 
                           send_data_5_port);
   send_data_reg_4_inst : DFFPOSX1 port map( D => n194, CLK => clk, Q => 
                           send_data_4_port);
   send_data_reg_3_inst : DFFPOSX1 port map( D => n195, CLK => clk, Q => 
                           send_data_3_port);
   send_data_reg_2_inst : DFFPOSX1 port map( D => n196, CLK => clk, Q => 
                           send_data_2_port);
   send_data_reg_1_inst : DFFPOSX1 port map( D => n197, CLK => clk, Q => 
                           send_data_1_port);
   send_data_reg_0_inst : DFFPOSX1 port map( D => n198, CLK => clk, Q => 
                           send_data_0_port);
   r80 : tx_tcu_0_DW01_inc_0 port map( A(6) => N188, A(5) => count_5_port, A(4)
                           => count_4_port, A(3) => count_3_port, A(2) => 
                           count_2_port, A(1) => count_1_port, A(0) => 
                           count_0_port, SUM(6) => N65, SUM(5) => N64, SUM(4) 
                           => N63, SUM(3) => N62, SUM(2) => N61, SUM(1) => N60,
                           SUM(0) => N59);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n15, S => n10, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n15, S => n9, Q => state_1_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n15, S => n8, Q => state_0_port);
   count_reg_3_inst : DFFSR port map( D => n180, CLK => clk, R => n15, S => n7,
                           Q => count_3_port);
   count_reg_2_inst : DFFSR port map( D => n181, CLK => clk, R => n15, S => n6,
                           Q => count_2_port);
   count_reg_1_inst : DFFSR port map( D => n182, CLK => clk, R => n15, S => n5,
                           Q => count_1_port);
   count_reg_0_inst : DFFSR port map( D => n176, CLK => clk, R => n15, S => n4,
                           Q => count_0_port);
   count_reg_4_inst : DFFSR port map( D => n179, CLK => clk, R => n15, S => n3,
                           Q => count_4_port);
   count_reg_5_inst : DFFSR port map( D => n178, CLK => clk, R => n15, S => n2,
                           Q => count_5_port);
   count_reg_6_inst : DFFSR port map( D => n177, CLK => clk, R => n15, S => n1,
                           Q => N188);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   U13 : INVX2 port map( A => n12, Y => n15);
   U14 : BUFX2 port map( A => rst, Y => n13);
   U15 : BUFX2 port map( A => rst, Y => n12);
   U16 : BUFX2 port map( A => rst, Y => n14);
   U17 : INVX2 port map( A => N188, Y => n11);
   U18 : XOR2X1 port map( A => N188, B => r81_carry_6_port, Y => N90);
   U19 : AND2X1 port map( A => count_5_port, B => r81_carry_5_port, Y => 
                           r81_carry_6_port);
   U20 : XOR2X1 port map( A => r81_carry_5_port, B => count_5_port, Y => N89);
   U21 : AND2X1 port map( A => count_4_port, B => r81_carry_4_port, Y => 
                           r81_carry_5_port);
   U22 : XOR2X1 port map( A => r81_carry_4_port, B => count_4_port, Y => N88);
   U23 : AND2X1 port map( A => count_3_port, B => r81_carry_3_port, Y => 
                           r81_carry_4_port);
   U24 : XOR2X1 port map( A => r81_carry_3_port, B => count_3_port, Y => N87);
   U25 : AND2X1 port map( A => count_2_port, B => r81_carry_2_port, Y => 
                           r81_carry_3_port);
   U26 : XOR2X1 port map( A => r81_carry_2_port, B => count_2_port, Y => N86);
   U27 : AND2X1 port map( A => count_1_port, B => r81_carry_1_port, Y => 
                           r81_carry_2_port);
   U28 : XOR2X1 port map( A => r81_carry_1_port, B => count_1_port, Y => N85);
   U29 : AND2X1 port map( A => count_0_port, B => r81_B_0_port, Y => 
                           r81_carry_1_port);
   U30 : XOR2X1 port map( A => r81_B_0_port, B => count_0_port, Y => N84);
   U31 : NOR2X1 port map( A => n16, B => n17, Y => t_strobe);
   U32 : NAND2X1 port map( A => n18, B => n19, Y => n17);
   U33 : NAND2X1 port map( A => n11, B => n20, Y => n16);
   U34 : OR2X1 port map( A => n21, B => n22, Y => sending);
   U35 : OAI21X1 port map( A => N188, B => n23, C => n24, Y => n22);
   U36 : NAND3X1 port map( A => n25, B => n26, C => n27, Y => n21);
   U37 : NAND3X1 port map( A => n28, B => n27, C => n29, Y => nextstate_2_port)
                           ;
   U38 : AOI22X1 port map( A => n30, B => p_ready, C => n31, D => n32, Y => n29
                           );
   U39 : NOR2X1 port map( A => state_1_port, B => state_0_port, Y => n30);
   U40 : NAND3X1 port map( A => n33, B => n34, C => n35, Y => nextstate_1_port)
                           ;
   U41 : AOI22X1 port map( A => n36, B => n18, C => n31, D => n37, Y => n35);
   U42 : INVX1 port map( A => n38, Y => n36);
   U43 : NAND3X1 port map( A => n39, B => n40, C => p_ready, Y => n33);
   U44 : NAND3X1 port map( A => n41, B => n28, C => n42, Y => nextstate_0_port)
                           ;
   U45 : AOI21X1 port map( A => n18, B => n38, C => n43, Y => n42);
   U46 : OAI21X1 port map( A => n44, B => n27, C => n45, Y => n43);
   U47 : NAND3X1 port map( A => p_ready, B => n37, C => n31, Y => n45);
   U48 : AND2X1 port map( A => n46, B => n47, Y => n31);
   U49 : INVX1 port map( A => n48, Y => n44);
   U50 : NAND3X1 port map( A => n19, B => n11, C => count_0_port, Y => n38);
   U51 : INVX1 port map( A => n49, Y => n28);
   U52 : AND2X1 port map( A => n26, B => n25, Y => n41);
   U53 : OAI21X1 port map( A => n50, B => n51, C => n52, Y => next_byte);
   U54 : MUX2X1 port map( B => n53, A => n54, S => n55, Y => n152);
   U55 : INVX1 port map( A => n56, Y => n153);
   U56 : MUX2X1 port map( B => PRGA_OUT(6), A => flop_data_6_port, S => n55, Y 
                           => n56);
   U57 : INVX1 port map( A => n57, Y => n154);
   U58 : MUX2X1 port map( B => PRGA_OUT(5), A => flop_data_5_port, S => n55, Y 
                           => n57);
   U59 : INVX1 port map( A => n58, Y => n155);
   U60 : MUX2X1 port map( B => PRGA_OUT(4), A => flop_data_4_port, S => n55, Y 
                           => n58);
   U61 : INVX1 port map( A => n59_port, Y => n156);
   U62 : MUX2X1 port map( B => PRGA_OUT(3), A => flop_data_3_port, S => n55, Y 
                           => n59_port);
   U63 : INVX1 port map( A => n60_port, Y => n157);
   U64 : MUX2X1 port map( B => PRGA_OUT(2), A => flop_data_2_port, S => n55, Y 
                           => n60_port);
   U65 : INVX1 port map( A => n61_port, Y => n174);
   U66 : MUX2X1 port map( B => PRGA_OUT(1), A => flop_data_1_port, S => n55, Y 
                           => n61_port);
   U67 : INVX1 port map( A => n62_port, Y => n175);
   U68 : MUX2X1 port map( B => PRGA_OUT(0), A => flop_data_0_port, S => n55, Y 
                           => n62_port);
   U69 : NAND3X1 port map( A => n63_port, B => n23, C => n64_port, Y => n55);
   U70 : AND2X1 port map( A => n24, B => n52, Y => n64_port);
   U71 : MUX2X1 port map( B => n65_port, A => n66, S => n40, Y => n52);
   U72 : NOR2X1 port map( A => p_ready, B => n67, Y => n66);
   U73 : NOR2X1 port map( A => n14, B => n65_port, Y => n63_port);
   U74 : INVX1 port map( A => t_bitstuff, Y => r81_B_0_port);
   U75 : OAI21X1 port map( A => n20, B => n68, C => n69, Y => n176);
   U76 : AOI22X1 port map( A => N59, B => n70, C => N84, D => n71, Y => n69);
   U77 : OAI21X1 port map( A => n11, B => n68, C => n72, Y => n177);
   U78 : AOI22X1 port map( A => N65, B => n70, C => N90, D => n71, Y => n72);
   U79 : OAI21X1 port map( A => n73, B => n68, C => n74, Y => n178);
   U80 : AOI22X1 port map( A => N64, B => n70, C => N89, D => n71, Y => n74);
   U81 : OAI21X1 port map( A => n75, B => n68, C => n76, Y => n179);
   U82 : AOI22X1 port map( A => N63, B => n70, C => N88, D => n71, Y => n76);
   U83 : OAI21X1 port map( A => n77, B => n68, C => n78, Y => n180);
   U84 : AOI22X1 port map( A => N62, B => n70, C => N87, D => n71, Y => n78);
   U85 : OAI21X1 port map( A => n79, B => n68, C => n80, Y => n181);
   U86 : AOI22X1 port map( A => N61, B => n70, C => N86, D => n71, Y => n80);
   U87 : OAI21X1 port map( A => n81, B => n68, C => n82, Y => n182);
   U88 : AOI22X1 port map( A => N60, B => n70, C => N85, D => n71, Y => n82);
   U89 : OAI21X1 port map( A => n32, B => n51, C => n34, Y => n71);
   U90 : OR2X1 port map( A => n25, B => n48, Y => n34);
   U91 : NAND3X1 port map( A => state_0_port, B => n83, C => state_1_port, Y =>
                           n25);
   U92 : INVX1 port map( A => n37, Y => n32);
   U93 : NAND2X1 port map( A => n48, B => n50, Y => n37);
   U94 : AND2X1 port map( A => prga_opcode(1), B => prga_opcode(0), Y => n50);
   U95 : AND2X1 port map( A => n68, B => n84_port, Y => n70);
   U96 : OAI21X1 port map( A => n48, B => n27, C => n85_port, Y => n84_port);
   U97 : NOR2X1 port map( A => n18, B => n49, Y => n85_port);
   U98 : NOR2X1 port map( A => n86_port, B => n87_port, Y => n48);
   U99 : NAND3X1 port map( A => count_4_port, B => count_1_port, C => 
                           count_5_port, Y => n87_port);
   U100 : NAND3X1 port map( A => count_0_port, B => count_3_port, C => n88_port
                           , Y => n86_port);
   U101 : NOR2X1 port map( A => N188, B => n79, Y => n88_port);
   U102 : NAND2X1 port map( A => n18, B => t_bitstuff, Y => n68);
   U103 : INVX1 port map( A => count_1_port, Y => n81);
   U104 : OAI21X1 port map( A => n89_port, B => n90_port, C => n91, Y => n183);
   U105 : INVX1 port map( A => current_send_data_7_port, Y => n90_port);
   U106 : OAI21X1 port map( A => n89_port, B => n92, C => n93, Y => n184);
   U107 : INVX1 port map( A => current_send_data_6_port, Y => n92);
   U108 : OAI21X1 port map( A => n89_port, B => n94, C => n95, Y => n185);
   U109 : INVX1 port map( A => current_send_data_5_port, Y => n94);
   U110 : OAI21X1 port map( A => n89_port, B => n96, C => n97, Y => n186);
   U111 : INVX1 port map( A => current_send_data_4_port, Y => n96);
   U112 : OAI21X1 port map( A => n89_port, B => n98, C => n99, Y => n187);
   U113 : INVX1 port map( A => current_send_data_3_port, Y => n98);
   U114 : OAI21X1 port map( A => n89_port, B => n100, C => n101, Y => n188_port
                           );
   U115 : INVX1 port map( A => current_send_data_2_port, Y => n100);
   U116 : OAI21X1 port map( A => n89_port, B => n102, C => n103, Y => n189);
   U117 : INVX1 port map( A => current_send_data_1_port, Y => n102);
   U118 : OAI21X1 port map( A => n89_port, B => n104, C => n105, Y => n190);
   U119 : INVX1 port map( A => current_send_data_0_port, Y => n104);
   U120 : AOI21X1 port map( A => state_0_port, B => state_1_port, C => n13, Y 
                           => n89_port);
   U121 : NAND2X1 port map( A => n106, B => n91, Y => n191);
   U122 : NOR2X1 port map( A => n107, B => n108, Y => n91);
   U123 : OAI21X1 port map( A => n53, B => n109, C => n110, Y => n108);
   U124 : NAND2X1 port map( A => t_crc(15), B => n111, Y => n110);
   U125 : INVX1 port map( A => n112, Y => n109);
   U126 : INVX1 port map( A => PRGA_OUT(7), Y => n53);
   U127 : OAI22X1 port map( A => n54, B => n113, C => n114, D => n115, Y => 
                           n107);
   U128 : NAND2X1 port map( A => n116, B => state_0_port, Y => n115);
   U129 : OAI21X1 port map( A => N188, B => t_crc(7), C => n15, Y => n114);
   U130 : INVX1 port map( A => n117, Y => n113);
   U131 : INVX1 port map( A => flop_data_7_port, Y => n54);
   U132 : AOI22X1 port map( A => n118, B => current_send_data_7_port, C => 
                           send_data_7_port, D => n12, Y => n106);
   U133 : NAND2X1 port map( A => n119, B => n93, Y => n192);
   U134 : AND2X1 port map( A => n120, B => n121, Y => n93);
   U135 : AOI22X1 port map( A => t_crc(6), B => n122, C => n117, D => 
                           flop_data_6_port, Y => n121);
   U136 : AOI22X1 port map( A => t_crc(14), B => n111, C => n112, D => 
                           PRGA_OUT(6), Y => n120);
   U137 : AOI22X1 port map( A => n118, B => current_send_data_6_port, C => 
                           send_data_6_port, D => n12, Y => n119);
   U138 : NAND2X1 port map( A => n123, B => n95, Y => n193);
   U139 : AND2X1 port map( A => n124, B => n125, Y => n95);
   U140 : AOI22X1 port map( A => t_crc(5), B => n122, C => n117, D => 
                           flop_data_5_port, Y => n125);
   U141 : AOI22X1 port map( A => t_crc(13), B => n111, C => n112, D => 
                           PRGA_OUT(5), Y => n124);
   U142 : AOI22X1 port map( A => n118, B => current_send_data_5_port, C => 
                           send_data_5_port, D => n13, Y => n123);
   U143 : NAND2X1 port map( A => n126, B => n97, Y => n194);
   U144 : AND2X1 port map( A => n127, B => n128, Y => n97);
   U145 : AOI22X1 port map( A => t_crc(4), B => n122, C => n117, D => 
                           flop_data_4_port, Y => n128);
   U146 : AOI22X1 port map( A => t_crc(12), B => n111, C => n112, D => 
                           PRGA_OUT(4), Y => n127);
   U147 : AOI22X1 port map( A => n118, B => current_send_data_4_port, C => 
                           send_data_4_port, D => n13, Y => n126);
   U148 : NAND2X1 port map( A => n129, B => n99, Y => n195);
   U149 : AND2X1 port map( A => n130, B => n131, Y => n99);
   U150 : AOI22X1 port map( A => t_crc(3), B => n122, C => n117, D => 
                           flop_data_3_port, Y => n131);
   U151 : AOI22X1 port map( A => t_crc(11), B => n111, C => n112, D => 
                           PRGA_OUT(3), Y => n130);
   U152 : AOI22X1 port map( A => n118, B => current_send_data_3_port, C => 
                           send_data_3_port, D => n13, Y => n129);
   U153 : NAND2X1 port map( A => n132, B => n101, Y => n196);
   U154 : AND2X1 port map( A => n133, B => n134, Y => n101);
   U155 : AOI22X1 port map( A => t_crc(2), B => n122, C => n117, D => 
                           flop_data_2_port, Y => n134);
   U156 : AOI22X1 port map( A => t_crc(10), B => n111, C => n112, D => 
                           PRGA_OUT(2), Y => n133);
   U157 : AOI22X1 port map( A => n118, B => current_send_data_2_port, C => 
                           send_data_2_port, D => n13, Y => n132);
   U158 : NAND2X1 port map( A => n135, B => n103, Y => n197);
   U159 : AND2X1 port map( A => n136, B => n137, Y => n103);
   U160 : AOI22X1 port map( A => t_crc(1), B => n122, C => n117, D => 
                           flop_data_1_port, Y => n137);
   U161 : AOI22X1 port map( A => t_crc(9), B => n111, C => n112, D => 
                           PRGA_OUT(1), Y => n136);
   U162 : AOI22X1 port map( A => n118, B => current_send_data_1_port, C => 
                           send_data_1_port, D => n13, Y => n135);
   U163 : NAND2X1 port map( A => n138, B => n105, Y => n198);
   U164 : AND2X1 port map( A => n139, B => n140, Y => n105);
   U165 : AOI22X1 port map( A => t_crc(0), B => n122, C => n117, D => 
                           flop_data_0_port, Y => n140);
   U166 : NOR2X1 port map( A => n24, B => n13, Y => n117);
   U167 : NOR2X1 port map( A => n46, B => n18, Y => n24);
   U168 : NOR2X1 port map( A => n40, B => n67, Y => n18);
   U169 : INVX1 port map( A => n39, Y => n67);
   U170 : NOR2X1 port map( A => state_1_port, B => state_2_port, Y => n39);
   U171 : INVX1 port map( A => n51, Y => n46);
   U172 : INVX1 port map( A => n141, Y => n122);
   U173 : NAND3X1 port map( A => n116, B => state_0_port, C => n142, Y => n141)
                           ;
   U174 : NOR2X1 port map( A => n14, B => N188, Y => n142);
   U175 : AOI22X1 port map( A => t_crc(8), B => n111, C => n112, D => 
                           PRGA_OUT(0), Y => n139);
   U176 : NOR2X1 port map( A => n26, B => n13, Y => n112);
   U177 : NAND2X1 port map( A => n65_port, B => n40, Y => n26);
   U178 : NOR2X1 port map( A => n83, B => n143, Y => n65_port);
   U179 : INVX1 port map( A => state_1_port, Y => n143);
   U180 : NOR2X1 port map( A => n27, B => n14, Y => n111);
   U181 : NAND2X1 port map( A => n116, B => n40, Y => n27);
   U182 : AOI22X1 port map( A => n118, B => current_send_data_0_port, C => 
                           send_data_0_port, D => n12, Y => n138);
   U183 : INVX1 port map( A => n144, Y => n118);
   U184 : NAND3X1 port map( A => state_0_port, B => n15, C => state_1_port, Y 
                           => n144);
   U185 : OAI21X1 port map( A => n51, B => n47, C => n145, Y => EOP);
   U186 : NAND3X1 port map( A => N188, B => n146, C => n49, Y => n145);
   U187 : NOR2X1 port map( A => n23, B => n147, Y => n49);
   U188 : OAI21X1 port map( A => n148, B => n149, C => state_0_port, Y => n147)
                           ;
   U189 : NAND3X1 port map( A => count_2_port, B => N188, C => count_3_port, Y 
                           => n149);
   U190 : NAND3X1 port map( A => n75, B => n73, C => n150, Y => n148);
   U191 : NOR2X1 port map( A => count_1_port, B => count_0_port, Y => n150);
   U192 : INVX1 port map( A => count_5_port, Y => n73);
   U193 : INVX1 port map( A => count_4_port, Y => n75);
   U194 : INVX1 port map( A => n116, Y => n23);
   U195 : NOR2X1 port map( A => n83, B => state_1_port, Y => n116);
   U196 : NAND3X1 port map( A => n19, B => n20, C => N188, Y => n47);
   U197 : INVX1 port map( A => count_0_port, Y => n20);
   U198 : NOR2X1 port map( A => n146, B => count_1_port, Y => n19);
   U199 : NAND3X1 port map( A => n79, B => n77, C => n151, Y => n146);
   U200 : NOR2X1 port map( A => count_5_port, B => count_4_port, Y => n151);
   U201 : INVX1 port map( A => count_3_port, Y => n77);
   U202 : INVX1 port map( A => count_2_port, Y => n79);
   U203 : NAND3X1 port map( A => n40, B => n83, C => state_1_port, Y => n51);
   U204 : INVX1 port map( A => state_2_port, Y => n83);
   U205 : INVX1 port map( A => state_0_port, Y => n40);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_shiftreg_0 is

   port( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe : in std_logic;  
         send_data : in std_logic_vector (7 downto 0);  d_encode : out 
         std_logic);

end tx_shiftreg_0;

architecture SYN_dataflow of tx_shiftreg_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal d_encode_port, present_val_7_port, present_val_6_port, 
      present_val_5_port, present_val_4_port, present_val_3_port, 
      present_val_2_port, present_val_1_port, count_2_port, count_1_port, 
      count_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n11, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83 : std_logic;

begin
   d_encode <= d_encode_port;
   
   count_reg_0_inst : DFFSR port map( D => n55, CLK => clk, R => n81, S => n14,
                           Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => n57, CLK => clk, R => n82, S => n14,
                           Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n56, CLK => clk, R => n83, S => n14,
                           Q => count_2_port);
   n83 <= '1';
   n82 <= '1';
   n81 <= '1';
   U30 : OAI21X1 port map( A => n13, B => n54, C => n79, Y => n65);
   U31 : AOI22X1 port map( A => send_data(0), B => n17, C => present_val_1_port
                           , D => n15, Y => n79);
   U32 : OAI21X1 port map( A => n13, B => n21, C => n78, Y => n64);
   U33 : NAND2X1 port map( A => send_data(7), B => n17, Y => n78);
   U34 : OAI21X1 port map( A => n13, B => n22, C => n77, Y => n63);
   U35 : AOI22X1 port map( A => send_data(6), B => n17, C => present_val_7_port
                           , D => n15, Y => n77);
   U36 : OAI21X1 port map( A => n13, B => n23, C => n76, Y => n62);
   U37 : AOI22X1 port map( A => send_data(5), B => n17, C => present_val_6_port
                           , D => n15, Y => n76);
   U38 : OAI21X1 port map( A => n13, B => n24, C => n75, Y => n61);
   U39 : AOI22X1 port map( A => send_data(4), B => n17, C => present_val_5_port
                           , D => n15, Y => n75);
   U40 : OAI21X1 port map( A => n13, B => n25, C => n74, Y => n60);
   U41 : AOI22X1 port map( A => send_data(3), B => n17, C => present_val_4_port
                           , D => n15, Y => n74);
   U42 : OAI21X1 port map( A => n13, B => n26, C => n73, Y => n59);
   U43 : AOI22X1 port map( A => send_data(2), B => n17, C => present_val_3_port
                           , D => n15, Y => n73);
   U44 : OAI21X1 port map( A => n27, B => n13, C => n72, Y => n58);
   U45 : AOI22X1 port map( A => send_data(1), B => n17, C => present_val_2_port
                           , D => n15, Y => n72);
   U46 : OAI21X1 port map( A => n71, B => n70, C => n69, Y => n57);
   U47 : OAI21X1 port map( A => n18, B => n11, C => count_1_port, Y => n69);
   U48 : NAND2X1 port map( A => count_0_port, B => n19, Y => n70);
   U49 : OAI21X1 port map( A => n17, B => n20, C => n68, Y => n56);
   U50 : NAND3X1 port map( A => count_1_port, B => count_0_port, C => n15, Y =>
                           n68);
   U51 : OAI22X1 port map( A => n18, B => n13, C => count_0_port, D => n71, Y 
                           => n55);
   U52 : NAND2X1 port map( A => n13, B => n67, Y => n71);
   U53 : OAI21X1 port map( A => t_bitstuff, B => n16, C => n67, Y => n80);
   U54 : NAND3X1 port map( A => SHIFT_ENABLE_R, B => count_0_port, C => n66, Y 
                           => n67);
   U55 : NOR2X1 port map( A => n19, B => n20, Y => n66);
   present_val_reg_7_inst : DFFSR port map( D => n64, CLK => clk, R => n14, S 
                           => n8, Q => present_val_7_port);
   present_val_reg_1_inst : DFFSR port map( D => n58, CLK => clk, R => n14, S 
                           => n7, Q => present_val_1_port);
   present_val_reg_6_inst : DFFSR port map( D => n63, CLK => clk, R => n14, S 
                           => n6, Q => present_val_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n62, CLK => clk, R => n14, S 
                           => n5, Q => present_val_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n61, CLK => clk, R => n14, S 
                           => n4, Q => present_val_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n60, CLK => clk, R => n14, S 
                           => n3, Q => present_val_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n59, CLK => clk, R => n14, S 
                           => n2, Q => present_val_2_port);
   present_val_reg_0_inst : DFFSR port map( D => n65, CLK => clk, R => n14, S 
                           => n1, Q => d_encode_port);
   U3 : INVX4 port map( A => n11, Y => n13);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   U15 : INVX2 port map( A => rst, Y => n14);
   U16 : INVX2 port map( A => n67, Y => n17);
   U17 : INVX2 port map( A => n80, Y => n11);
   U18 : INVX2 port map( A => n71, Y => n15);
   U19 : INVX2 port map( A => SHIFT_ENABLE_R, Y => n16);
   U20 : INVX2 port map( A => count_0_port, Y => n18);
   U21 : INVX2 port map( A => count_1_port, Y => n19);
   U22 : INVX2 port map( A => count_2_port, Y => n20);
   U23 : INVX2 port map( A => present_val_7_port, Y => n21);
   U24 : INVX2 port map( A => present_val_6_port, Y => n22);
   U25 : INVX2 port map( A => present_val_5_port, Y => n23);
   U26 : INVX2 port map( A => present_val_4_port, Y => n24);
   U27 : INVX2 port map( A => present_val_3_port, Y => n25);
   U28 : INVX2 port map( A => present_val_2_port, Y => n26);
   U29 : INVX2 port map( A => present_val_1_port, Y => n27);
   U56 : INVX2 port map( A => d_encode_port, Y => n54);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_encode_0 is

   port( clk, rst, SHIFT_ENABLE_E, d_encode, EOP : in std_logic;  t_bitstuff, 
         dp_tx_out, dm_tx_out : out std_logic);

end tx_encode_0;

architecture SYN_moore of tx_encode_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal DE_holdout, DE_holdout_BS, state_3_port, state_2_port, state_1_port, 
      state_0_port, nextstate_3_port, nextstate_2_port, nextstate_1_port, 
      nextstate_0_port, DE_holdout_last, DE_holdout_nxt, dm_tx_nxt, n2, n4, n7,
      n8, n10, n11, n16, n17, n21, n25, n28, n29, n30, n31, n34, n35, n42, n53,
      n54, n56, n57, n58, n59, n60, n63, n66, n67, n68, n69, n70, n71, n72, n73
      , n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, 
      n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
      n102, n103, n104 : std_logic;

begin
   
   DE_holdout_reg : DFFSR port map( D => DE_holdout_nxt, CLK => clk, R => n67, 
                           S => n16, Q => DE_holdout);
   DE_holdout_last_reg : DFFPOSX1 port map( D => n68, CLK => clk, Q => 
                           DE_holdout_last);
   dp_tx_out_reg : DFFSR port map( D => DE_holdout_nxt, CLK => clk, R => n69, S
                           => n16, Q => dp_tx_out);
   U3 : AOI21X1 port map( A => state_3_port, B => n104, C => n30, Y => 
                           nextstate_3_port);
   U4 : OAI21X1 port map( A => n103, B => n60, C => n102, Y => nextstate_2_port
                           );
   U5 : AOI21X1 port map( A => n101, B => n17, C => n34, Y => n102);
   U7 : NOR2X1 port map( A => state_2_port, B => n59, Y => n101);
   U8 : AOI21X1 port map( A => n35, B => n59, C => n99, Y => n103);
   U9 : OAI21X1 port map( A => state_1_port, B => n100, C => n98, Y => 
                           nextstate_1_port);
   U10 : AOI21X1 port map( A => state_1_port, B => n97, C => n34, Y => n98);
   U11 : OAI21X1 port map( A => state_0_port, B => n96, C => n21, Y => n97);
   U12 : NAND3X1 port map( A => SHIFT_ENABLE_E, B => n35, C => state_0_port, Y 
                           => n100);
   U14 : OAI21X1 port map( A => n58, B => n21, C => n95, Y => nextstate_0_port)
                           ;
   U15 : OAI21X1 port map( A => n94, B => n93, C => SHIFT_ENABLE_E, Y => n95);
   U16 : OAI21X1 port map( A => n31, B => n92, C => n91, Y => n93);
   U17 : NAND2X1 port map( A => n90, B => n42, Y => n92);
   U18 : NOR2X1 port map( A => state_0_port, B => n96, Y => n94);
   U19 : NAND3X1 port map( A => d_encode, B => n89, C => n88, Y => n96);
   U20 : XNOR2X1 port map( A => n54, B => n53, Y => n88);
   U22 : NOR2X1 port map( A => n31, B => SHIFT_ENABLE_E, Y => n99);
   U23 : OAI22X1 port map( A => n16, B => n54, C => rst, D => n53, Y => n68);
   U26 : OAI22X1 port map( A => n25, B => n63, C => n53, D => n87, Y => n66);
   U28 : NAND2X1 port map( A => n34, B => SHIFT_ENABLE_E, Y => n87);
   U30 : NAND3X1 port map( A => n90, B => n58, C => n89, Y => n91);
   U31 : NOR2X1 port map( A => state_3_port, B => n86, Y => t_bitstuff);
   U32 : OAI21X1 port map( A => n57, B => n56, C => n85, Y => dm_tx_nxt);
   U33 : AOI22X1 port map( A => n84, B => n90, C => n83, D => n82, Y => n85);
   U34 : NOR2X1 port map( A => n90, B => n31, Y => n83);
   U36 : NOR2X1 port map( A => EOP, B => state_3_port, Y => n89);
   U37 : NOR2X1 port map( A => EOP, B => n81, Y => n84);
   U38 : AOI22X1 port map( A => state_0_port, B => n80, C => n28, D => n58, Y 
                           => n81);
   U40 : XNOR2X1 port map( A => DE_holdout_BS, B => n78, Y => n80);
   U41 : OAI21X1 port map( A => n57, B => n56, C => n77, Y => DE_holdout_nxt);
   U42 : OAI21X1 port map( A => n76, B => n75, C => n30, Y => n77);
   U44 : OAI21X1 port map( A => n90, B => n82, C => n74, Y => n75);
   U45 : NAND3X1 port map( A => n79, B => n58, C => n90, Y => n74);
   U46 : XOR2X1 port map( A => DE_holdout, B => SHIFT_ENABLE_E, Y => n79);
   U47 : XNOR2X1 port map( A => n73, B => n53, Y => n82);
   U49 : NAND2X1 port map( A => SHIFT_ENABLE_E, B => n42, Y => n73);
   U51 : OAI21X1 port map( A => n86, B => n72, C => n71, Y => n76);
   U52 : AOI21X1 port map( A => n70, B => n29, C => state_3_port, Y => n71);
   U54 : NOR2X1 port map( A => n63, B => n86, Y => n70);
   U55 : NAND2X1 port map( A => n78, B => n63, Y => n72);
   U57 : NAND2X1 port map( A => SHIFT_ENABLE_E, B => d_encode, Y => n78);
   U58 : NAND2X1 port map( A => state_0_port, B => n90, Y => n86);
   U59 : NOR2X1 port map( A => n60, B => n59, Y => n90);
   U62 : NAND3X1 port map( A => n59, B => n60, C => n58, Y => n104);
   n69 <= '1';
   n67 <= '1';
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => clk, R => 
                           n16, S => n11, Q => state_3_port);
   dm_tx_out_reg : DFFSR port map( D => dm_tx_nxt, CLK => clk, R => n16, S => 
                           n10, Q => dm_tx_out);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n16, S => n8, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n16, S => n7, Q => state_1_port);
   DE_holdout_BS_reg : DFFSR port map( D => n66, CLK => clk, R => n16, S => n4,
                           Q => DE_holdout_BS);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n16, S => n2, Q => state_2_port);
   n2 <= '1';
   n4 <= '1';
   n7 <= '1';
   n8 <= '1';
   n10 <= '1';
   n11 <= '1';
   U29 : INVX2 port map( A => rst, Y => n16);
   U35 : INVX2 port map( A => n100, Y => n17);
   U39 : INVX2 port map( A => n99, Y => n21);
   U43 : INVX2 port map( A => n87, Y => n25);
   U48 : INVX2 port map( A => n79, Y => n28);
   U50 : INVX2 port map( A => n78, Y => n29);
   U53 : INVX2 port map( A => EOP, Y => n30);
   U56 : INVX2 port map( A => n89, Y => n31);
   U60 : INVX2 port map( A => n91, Y => n34);
   U61 : INVX2 port map( A => n96, Y => n35);
   U63 : INVX2 port map( A => d_encode, Y => n42);
   U64 : INVX2 port map( A => DE_holdout, Y => n53);
   U65 : INVX2 port map( A => DE_holdout_last, Y => n54);
   U66 : INVX2 port map( A => state_3_port, Y => n56);
   U68 : INVX2 port map( A => n104, Y => n57);
   U69 : INVX2 port map( A => state_0_port, Y => n58);
   U70 : INVX2 port map( A => state_1_port, Y => n59);
   U71 : INVX2 port map( A => state_2_port, Y => n60);
   U72 : INVX2 port map( A => DE_holdout_BS, Y => n63);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_CRC_CALC_0 is

   port( CLK, RST, EOP, T_STROBE : in std_logic;  PRGA_OPCODE : in 
         std_logic_vector (1 downto 0);  PRGA_OUT : in std_logic_vector (7 
         downto 0);  TX_CRC : out std_logic_vector (15 downto 0));

end tx_CRC_CALC_0;

architecture SYN_txcrcm of tx_CRC_CALC_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal TX_CRC_15_port, TX_CRC_14_port, TX_CRC_13_port, TX_CRC_12_port, 
      TX_CRC_11_port, TX_CRC_10_port, TX_CRC_9_port, TX_CRC_8_port, 
      TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port, TX_CRC_4_port, TX_CRC_3_port
      , TX_CRC_2_port, TX_CRC_1_port, TX_CRC_0_port, n1, n2, n3, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22
      , n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
      n37, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122 : std_logic;

begin
   TX_CRC <= ( TX_CRC_15_port, TX_CRC_14_port, TX_CRC_13_port, TX_CRC_12_port, 
      TX_CRC_11_port, TX_CRC_10_port, TX_CRC_9_port, TX_CRC_8_port, 
      TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port, TX_CRC_4_port, TX_CRC_3_port
      , TX_CRC_2_port, TX_CRC_1_port, TX_CRC_0_port );
   
   U39 : OAI22X1 port map( A => n25, B => n20, C => n122, D => n19, Y => n97);
   U40 : XNOR2X1 port map( A => n120, B => n80, Y => n122);
   U41 : OAI22X1 port map( A => n79, B => n20, C => n19, D => n37, Y => n96);
   U42 : OAI22X1 port map( A => n36, B => n20, C => n19, D => n35, Y => n95);
   U43 : OAI22X1 port map( A => n34, B => n20, C => n19, D => n33, Y => n94);
   U44 : OAI22X1 port map( A => n32, B => n20, C => n19, D => n31, Y => n93);
   U45 : OAI22X1 port map( A => n29, B => n20, C => n19, D => n28, Y => n92);
   U46 : OAI22X1 port map( A => n27, B => n20, C => n119, D => n19, Y => n91);
   U47 : XNOR2X1 port map( A => TX_CRC_1_port, B => n118, Y => n119);
   U48 : OAI22X1 port map( A => n24, B => n20, C => n117, D => n19, Y => n90);
   U49 : XOR2X1 port map( A => n116, B => n115, Y => n117);
   U50 : XNOR2X1 port map( A => TX_CRC_0_port, B => n118, Y => n116);
   U51 : OAI22X1 port map( A => n80, B => n20, C => n114, D => n19, Y => n89);
   U52 : OAI22X1 port map( A => n20, B => n37, C => n113, D => n19, Y => n88);
   U53 : XNOR2X1 port map( A => n112, B => n111, Y => n113);
   U54 : OAI22X1 port map( A => n20, B => n35, C => n110, D => n121, Y => n87);
   U55 : OAI22X1 port map( A => n20, B => n33, C => n109, D => n121, Y => n86);
   U56 : XNOR2X1 port map( A => n108, B => n107, Y => n109);
   U57 : OAI22X1 port map( A => n20, B => n31, C => n106, D => n121, Y => n85);
   U58 : OAI22X1 port map( A => n20, B => n28, C => n105, D => n121, Y => n84);
   U59 : XOR2X1 port map( A => n104, B => n103, Y => n105);
   U60 : OAI22X1 port map( A => n20, B => n26, C => n102, D => n121, Y => n83);
   U61 : XOR2X1 port map( A => n101, B => n100, Y => n102);
   U62 : XOR2X1 port map( A => n118, B => n114, Y => n101);
   U63 : OAI22X1 port map( A => n20, B => n23, C => n120, D => n121, Y => n82);
   U64 : XOR2X1 port map( A => n99, B => n98, Y => n120);
   U65 : XOR2X1 port map( A => n103, B => n118, Y => n98);
   U66 : XNOR2X1 port map( A => n25, B => PRGA_OUT(7), Y => n118);
   U67 : XNOR2X1 port map( A => n24, B => PRGA_OUT(0), Y => n103);
   U68 : XOR2X1 port map( A => n114, B => n100, Y => n99);
   U69 : XOR2X1 port map( A => n106, B => n110, Y => n100);
   U70 : XNOR2X1 port map( A => n107, B => n112, Y => n110);
   U71 : XOR2X1 port map( A => TX_CRC_12_port, B => PRGA_OUT(4), Y => n112);
   U72 : XOR2X1 port map( A => TX_CRC_11_port, B => PRGA_OUT(3), Y => n107);
   U73 : XNOR2X1 port map( A => n104, B => n30, Y => n106);
   U74 : XOR2X1 port map( A => TX_CRC_10_port, B => PRGA_OUT(2), Y => n108);
   U75 : XNOR2X1 port map( A => TX_CRC_9_port, B => PRGA_OUT(1), Y => n104);
   U76 : XNOR2X1 port map( A => n111, B => n115, Y => n114);
   U77 : XNOR2X1 port map( A => n79, B => PRGA_OUT(6), Y => n115);
   U78 : XOR2X1 port map( A => TX_CRC_13_port, B => PRGA_OUT(5), Y => n111);
   U80 : NAND3X1 port map( A => PRGA_OPCODE(0), B => n81, C => T_STROBE, Y => 
                           n121);
   current_crc_reg_6_inst : DFFSR port map( D => n88, CLK => CLK, R => n21, S 
                           => n17, Q => TX_CRC_6_port);
   current_crc_reg_5_inst : DFFSR port map( D => n87, CLK => CLK, R => n21, S 
                           => n16, Q => TX_CRC_5_port);
   current_crc_reg_4_inst : DFFSR port map( D => n86, CLK => CLK, R => n21, S 
                           => n15, Q => TX_CRC_4_port);
   current_crc_reg_3_inst : DFFSR port map( D => n85, CLK => CLK, R => n21, S 
                           => n14, Q => TX_CRC_3_port);
   current_crc_reg_2_inst : DFFSR port map( D => n84, CLK => CLK, R => n21, S 
                           => n13, Q => TX_CRC_2_port);
   current_crc_reg_1_inst : DFFSR port map( D => n83, CLK => CLK, R => n21, S 
                           => n12, Q => TX_CRC_1_port);
   current_crc_reg_0_inst : DFFSR port map( D => n82, CLK => CLK, R => n21, S 
                           => n11, Q => TX_CRC_0_port);
   current_crc_reg_15_inst : DFFSR port map( D => n97, CLK => CLK, R => n21, S 
                           => n10, Q => TX_CRC_15_port);
   current_crc_reg_14_inst : DFFSR port map( D => n96, CLK => CLK, R => n21, S 
                           => n9, Q => TX_CRC_14_port);
   current_crc_reg_13_inst : DFFSR port map( D => n95, CLK => CLK, R => n21, S 
                           => n8, Q => TX_CRC_13_port);
   current_crc_reg_12_inst : DFFSR port map( D => n94, CLK => CLK, R => n21, S 
                           => n7, Q => TX_CRC_12_port);
   current_crc_reg_11_inst : DFFSR port map( D => n93, CLK => CLK, R => n21, S 
                           => n6, Q => TX_CRC_11_port);
   current_crc_reg_10_inst : DFFSR port map( D => n92, CLK => CLK, R => n21, S 
                           => n5, Q => TX_CRC_10_port);
   current_crc_reg_9_inst : DFFSR port map( D => n91, CLK => CLK, R => n21, S 
                           => n4, Q => TX_CRC_9_port);
   current_crc_reg_8_inst : DFFSR port map( D => n90, CLK => CLK, R => n21, S 
                           => n3, Q => TX_CRC_8_port);
   current_crc_reg_7_inst : DFFSR port map( D => n89, CLK => CLK, R => n21, S 
                           => n2, Q => TX_CRC_7_port);
   U3 : AND2X2 port map( A => n19, B => n22, Y => n1);
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   U20 : INVX2 port map( A => n1, Y => n20);
   U21 : INVX2 port map( A => RST, Y => n21);
   U22 : INVX2 port map( A => n18, Y => n19);
   U23 : INVX2 port map( A => n121, Y => n18);
   U24 : INVX2 port map( A => EOP, Y => n22);
   U25 : INVX2 port map( A => TX_CRC_0_port, Y => n23);
   U26 : INVX2 port map( A => TX_CRC_8_port, Y => n24);
   U27 : INVX2 port map( A => TX_CRC_15_port, Y => n25);
   U28 : INVX2 port map( A => TX_CRC_1_port, Y => n26);
   U29 : INVX2 port map( A => TX_CRC_9_port, Y => n27);
   U30 : INVX2 port map( A => TX_CRC_2_port, Y => n28);
   U31 : INVX2 port map( A => TX_CRC_10_port, Y => n29);
   U32 : INVX2 port map( A => n108, Y => n30);
   U33 : INVX2 port map( A => TX_CRC_3_port, Y => n31);
   U34 : INVX2 port map( A => TX_CRC_11_port, Y => n32);
   U35 : INVX2 port map( A => TX_CRC_4_port, Y => n33);
   U36 : INVX2 port map( A => TX_CRC_12_port, Y => n34);
   U37 : INVX2 port map( A => TX_CRC_5_port, Y => n35);
   U38 : INVX2 port map( A => TX_CRC_13_port, Y => n36);
   U79 : INVX2 port map( A => TX_CRC_6_port, Y => n37);
   U81 : INVX2 port map( A => TX_CRC_14_port, Y => n79);
   U82 : INVX2 port map( A => TX_CRC_7_port, Y => n80);
   U83 : INVX2 port map( A => PRGA_OPCODE(1), Y => n81);

end SYN_txcrcm;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_timer_0 is

   port( CLK, RST, D_EDGE, RCVING : in std_logic;  SHIFT_ENABLE : out std_logic
         );

end rx_timer_0;

architecture SYN_moore of rx_timer_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_3_port, count_2_port, count_1_port, count_0_port, state, 
      nextcount_3_port, nextcount_2_port, nextcount_1_port, nextcount_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n19, n20, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n33, n34 : std_logic;

begin
   
   U17 : NOR2X1 port map( A => n34, B => n33, Y => nextcount_3_port);
   U18 : AOI22X1 port map( A => n32, B => n31, C => n30, D => count_3_port, Y 
                           => n34);
   U19 : XOR2X1 port map( A => n29, B => n31, Y => n30);
   U20 : NOR2X1 port map( A => count_3_port, B => n20, Y => n32);
   U23 : NOR2X1 port map( A => n27, B => n33, Y => nextcount_1_port);
   U24 : NAND2X1 port map( A => state, B => n26, Y => nextcount_0_port);
   U25 : OAI21X1 port map( A => D_EDGE, B => n19, C => RCVING, Y => n26);
   U28 : NAND3X1 port map( A => RCVING, B => n25, C => state, Y => n33);
   U29 : OAI21X1 port map( A => n27, B => n24, C => n28, Y => n29);
   U30 : NAND2X1 port map( A => count_0_port, B => count_1_port, Y => n28);
   U31 : XOR2X1 port map( A => n24, B => n27, Y => n31);
   U32 : XNOR2X1 port map( A => count_0_port, B => count_1_port, Y => n27);
   state_reg : DFFSR port map( D => RCVING, CLK => CLK, R => n11, S => n5, Q =>
                           state);
   count_reg_2_inst : DFFSR port map( D => nextcount_2_port, CLK => CLK, R => 
                           n11, S => n4, Q => count_2_port);
   count_reg_0_inst : DFFSR port map( D => nextcount_0_port, CLK => CLK, R => 
                           n11, S => n3, Q => count_0_port);
   count_reg_3_inst : DFFSR port map( D => nextcount_3_port, CLK => CLK, R => 
                           n11, S => n2, Q => count_3_port);
   count_reg_1_inst : DFFSR port map( D => nextcount_1_port, CLK => CLK, R => 
                           n11, S => n1, Q => count_1_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   U8 : AND2X1 port map( A => n12, B => count_3_port, Y => n7);
   U9 : INVX2 port map( A => n8, Y => nextcount_2_port);
   U10 : INVX2 port map( A => RST, Y => n11);
   U11 : AND2X2 port map( A => n6, B => n7, Y => SHIFT_ENABLE);
   U12 : NOR2X1 port map( A => n31, B => n29, Y => n6);
   U13 : OAI21X1 port map( A => n9, B => n10, C => RCVING, Y => n8);
   U14 : NAND2X1 port map( A => n25, B => state, Y => n9);
   U15 : XNOR2X1 port map( A => n28, B => count_2_port, Y => n10);
   U16 : INVX2 port map( A => n33, Y => n12);
   U21 : INVX2 port map( A => count_0_port, Y => n19);
   U22 : INVX2 port map( A => n29, Y => n20);
   U26 : INVX2 port map( A => count_2_port, Y => n24);
   U27 : INVX2 port map( A => D_EDGE, Y => n25);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_shift_reg_0 is

   port( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF : in std_logic;  RCV_DATA : 
         out std_logic_vector (7 downto 0));

end rx_shift_reg_0;

architecture SYN_dataflow of rx_shift_reg_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      present_val_7_port, present_val_6_port, present_val_5_port, 
      present_val_4_port, present_val_3_port, present_val_2_port, 
      present_val_1_port, present_val_0_port, n1, n3, n5, n7, n9, n11, n13, n15
      , n17, n20, n22, n25, n28, n31, n34, n37, n40, n43, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   RCV_DATA_reg_7_inst : DFFPOSX1 port map( D => n47, CLK => CLK, Q => 
                           RCV_DATA_7_port);
   RCV_DATA_reg_6_inst : DFFPOSX1 port map( D => n49, CLK => CLK, Q => 
                           RCV_DATA_6_port);
   RCV_DATA_reg_5_inst : DFFPOSX1 port map( D => n51, CLK => CLK, Q => 
                           RCV_DATA_5_port);
   RCV_DATA_reg_4_inst : DFFPOSX1 port map( D => n53, CLK => CLK, Q => 
                           RCV_DATA_4_port);
   RCV_DATA_reg_3_inst : DFFPOSX1 port map( D => n55, CLK => CLK, Q => 
                           RCV_DATA_3_port);
   RCV_DATA_reg_2_inst : DFFPOSX1 port map( D => n57, CLK => CLK, Q => 
                           RCV_DATA_2_port);
   RCV_DATA_reg_1_inst : DFFPOSX1 port map( D => n59, CLK => CLK, Q => 
                           RCV_DATA_1_port);
   RCV_DATA_reg_0_inst : DFFPOSX1 port map( D => n61, CLK => CLK, Q => 
                           RCV_DATA_0_port);
   U2 : OAI21X1 port map( A => RST, B => n43, C => n71, Y => n61);
   U3 : NAND2X1 port map( A => RCV_DATA_0_port, B => RST, Y => n71);
   U4 : OAI22X1 port map( A => n20, B => n43, C => n70, D => n40, Y => n60);
   U6 : OAI21X1 port map( A => RST, B => n40, C => n69, Y => n59);
   U7 : NAND2X1 port map( A => RCV_DATA_1_port, B => RST, Y => n69);
   U8 : OAI22X1 port map( A => n20, B => n40, C => n70, D => n37, Y => n58);
   U10 : OAI21X1 port map( A => RST, B => n37, C => n68, Y => n57);
   U11 : NAND2X1 port map( A => RCV_DATA_2_port, B => RST, Y => n68);
   U12 : OAI22X1 port map( A => n20, B => n37, C => n70, D => n34, Y => n56);
   U14 : OAI21X1 port map( A => RST, B => n34, C => n67, Y => n55);
   U15 : NAND2X1 port map( A => RCV_DATA_3_port, B => RST, Y => n67);
   U16 : OAI22X1 port map( A => n20, B => n34, C => n70, D => n31, Y => n54);
   U18 : OAI21X1 port map( A => RST, B => n31, C => n66, Y => n53);
   U19 : NAND2X1 port map( A => RCV_DATA_4_port, B => RST, Y => n66);
   U20 : OAI22X1 port map( A => n20, B => n31, C => n70, D => n28, Y => n52);
   U22 : OAI21X1 port map( A => RST, B => n28, C => n65, Y => n51);
   U23 : NAND2X1 port map( A => RCV_DATA_5_port, B => RST, Y => n65);
   U24 : OAI22X1 port map( A => n20, B => n28, C => n70, D => n25, Y => n50);
   U26 : OAI21X1 port map( A => RST, B => n25, C => n64, Y => n49);
   U27 : NAND2X1 port map( A => RCV_DATA_6_port, B => RST, Y => n64);
   U28 : OAI22X1 port map( A => n20, B => n25, C => n70, D => n22, Y => n48);
   U30 : OAI21X1 port map( A => RST, B => n22, C => n63, Y => n47);
   U31 : NAND2X1 port map( A => RCV_DATA_7_port, B => RST, Y => n63);
   U32 : OAI21X1 port map( A => n20, B => n22, C => n62, Y => n46);
   U33 : NAND2X1 port map( A => D_ORIG, B => n20, Y => n62);
   U36 : NAND2X1 port map( A => SHIFT_ENABLE, B => n45, Y => n70);
   present_val_reg_7_inst : DFFSR port map( D => n46, CLK => CLK, R => n17, S 
                           => n15, Q => present_val_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n48, CLK => CLK, R => n17, S 
                           => n13, Q => present_val_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n50, CLK => CLK, R => n17, S 
                           => n11, Q => present_val_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n52, CLK => CLK, R => n17, S 
                           => n9, Q => present_val_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n54, CLK => CLK, R => n17, S 
                           => n7, Q => present_val_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n56, CLK => CLK, R => n17, S 
                           => n5, Q => present_val_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n58, CLK => CLK, R => n17, S 
                           => n3, Q => present_val_1_port);
   present_val_reg_0_inst : DFFSR port map( D => n60, CLK => CLK, R => n17, S 
                           => n1, Q => present_val_0_port);
   U5 : INVX2 port map( A => n70, Y => n20);
   n1 <= '1';
   n3 <= '1';
   n5 <= '1';
   n7 <= '1';
   n9 <= '1';
   n11 <= '1';
   n13 <= '1';
   n15 <= '1';
   U37 : INVX2 port map( A => RST, Y => n17);
   U38 : INVX2 port map( A => present_val_7_port, Y => n22);
   U39 : INVX2 port map( A => present_val_6_port, Y => n25);
   U40 : INVX2 port map( A => present_val_5_port, Y => n28);
   U41 : INVX2 port map( A => present_val_4_port, Y => n31);
   U42 : INVX2 port map( A => present_val_3_port, Y => n34);
   U43 : INVX2 port map( A => present_val_2_port, Y => n37);
   U44 : INVX2 port map( A => present_val_1_port, Y => n40);
   U45 : INVX2 port map( A => present_val_0_port, Y => n43);
   U46 : INVX2 port map( A => BITSTUFF, Y => n45);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_rcu_0 is

   port( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR : in std_logic
         ;  RX_CRC, RX_CHECK_CRC : in std_logic_vector (15 downto 0);  RCV_DATA
         : in std_logic_vector (7 downto 0);  RCVING, W_ENABLE, R_ERROR, 
         CRC_ERROR : out std_logic;  OPCODE : out std_logic_vector (1 downto 0)
         );

end rx_rcu_0;

architecture SYN_moore of rx_rcu_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal CRC_ERROR_port, OPCODE_1_port, OPCODE_0_port, state_3_port, 
      state_2_port, state_1_port, state_0_port, count_3_port, count_2_port, 
      count_1_port, count_0_port, nextstate_3_port, nextstate_2_port, 
      nextstate_1_port, nextstate_0_port, nxtR_ERROR, curR_ERROR, curCRC_ERROR,
      n1, n2, n3, n4, n5, n6, n7, n8, n10, n13, n17, n18, n19, n23, n24, n25, 
      n26, n28, n30, n35, n43, n44, n49, n58, n64, n68, n69, n73, n76, n82, n93
      , n101, n104, n108, n110, n112, n114, n115, n118, n124, n128, n130, n131,
      n132, n135, n141, n143, n148, n149, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297 : std_logic;

begin
   CRC_ERROR <= CRC_ERROR_port;
   OPCODE <= ( OPCODE_1_port, OPCODE_0_port );
   
   curCRC_ERROR_reg : DFFPOSX1 port map( D => n196, CLK => CLK, Q => 
                           curCRC_ERROR);
   curR_ERROR_reg : DFFPOSX1 port map( D => n197, CLK => CLK, Q => curR_ERROR);
   CRC_ERROR_reg : DFFPOSX1 port map( D => n172, CLK => CLK, Q => 
                           CRC_ERROR_port);
   U5 : OAI21X1 port map( A => EOP, B => n23, C => n294, Y => n295);
   U6 : AOI22X1 port map( A => BS_ERROR, B => n293, C => n292, D => n44, Y => 
                           n294);
   U7 : OAI21X1 port map( A => n192, B => n26, C => n291, Y => n292);
   U8 : AOI22X1 port map( A => n290, B => D_EDGE, C => n19, D => n289, Y => 
                           n291);
   U9 : OAI21X1 port map( A => n183, B => n190, C => n184, Y => n289);
   U11 : NOR2X1 port map( A => n183, B => n177, Y => n290);
   U12 : OAI21X1 port map( A => n288, B => n24, C => n287, Y => n293);
   U13 : OAI21X1 port map( A => n2, B => n286, C => n285, Y => n296);
   U15 : NAND2X1 port map( A => n178, B => n282, Y => n286);
   U16 : NAND2X1 port map( A => n281, B => n280, Y => nextstate_2_port);
   U17 : NOR2X1 port map( A => n279, B => n278, Y => n280);
   U18 : OAI21X1 port map( A => n26, B => n277, C => n283, Y => n278);
   U19 : OAI21X1 port map( A => n2, B => n276, C => n49, Y => n277);
   U20 : NAND2X1 port map( A => n179, B => n187, Y => n276);
   U21 : NAND2X1 port map( A => n275, B => n274, Y => n279);
   U22 : NOR2X1 port map( A => n273, B => n272, Y => n281);
   U23 : OAI22X1 port map( A => n171, B => n44, C => n271, D => n190, Y => n272
                           );
   U24 : OAI21X1 port map( A => n49, B => n270, C => n269, Y => n273);
   U25 : OAI21X1 port map( A => n268, B => n267, C => n266, Y => n269);
   U26 : AOI22X1 port map( A => n265, B => n264, C => n282, D => n192, Y => 
                           n270);
   U27 : NOR2X1 port map( A => D_EDGE, B => n183, Y => n265);
   U28 : OAI21X1 port map( A => n170, B => n192, C => n263, Y => 
                           nextstate_1_port);
   U30 : OAI21X1 port map( A => n260, B => n259, C => n190, Y => n262);
   U31 : OAI21X1 port map( A => n287, B => n180, C => n258, Y => n259);
   U33 : OAI21X1 port map( A => n23, B => n256, C => n175, Y => n260);
   U34 : NAND2X1 port map( A => n181, B => n192, Y => n256);
   U35 : OAI22X1 port map( A => n255, B => n254, C => n44, D => n253, Y => 
                           nextstate_0_port);
   U36 : OAI21X1 port map( A => n183, B => n28, C => n252, Y => n253);
   U37 : NAND3X1 port map( A => n190, B => n183, C => n251, Y => n252);
   U38 : OAI21X1 port map( A => n25, B => n192, C => n250, Y => n251);
   U39 : AOI22X1 port map( A => n257, B => n249, C => n248, D => n247, Y => 
                           n250);
   U42 : OAI22X1 port map( A => state_0_port, B => n184, C => n246, D => n183, 
                           Y => n254);
   U43 : AOI22X1 port map( A => EOP, B => n249, C => D_EDGE, D => n174, Y => 
                           n246);
   U45 : OAI21X1 port map( A => n35, B => n244, C => n243, Y => n255);
   U46 : NOR2X1 port map( A => n49, B => n282, Y => n243);
   U47 : AOI22X1 port map( A => n242, B => n257, C => D_EDGE, D => n249, Y => 
                           n244);
   U48 : NOR2X1 port map( A => n181, B => EOP, Y => n257);
   U50 : NOR2X1 port map( A => BS_ERROR, B => n25, Y => n242);
   U52 : AOI21X1 port map( A => CRC_ERROR_port, B => RST, C => n240, Y => n241)
                           ;
   U53 : OAI21X1 port map( A => n239, B => n238, C => n237, Y => n240);
   U54 : NAND2X1 port map( A => curCRC_ERROR, B => n236, Y => n238);
   U55 : NAND2X1 port map( A => n58, B => n44, Y => n239);
   U56 : OAI21X1 port map( A => n58, B => n189, C => n235, Y => n197);
   U57 : AOI21X1 port map( A => n297, B => n58, C => n173, Y => n235);
   U59 : NAND3X1 port map( A => n233, B => n44, C => curR_ERROR, Y => n234);
   U60 : OAI21X1 port map( A => n19, B => n183, C => n232, Y => n233);
   U61 : OAI21X1 port map( A => n178, B => n26, C => n231, Y => n297);
   U64 : OAI21X1 port map( A => n19, B => n247, C => n177, Y => n229);
   U65 : OAI21X1 port map( A => n267, B => n176, C => EOP, Y => n230);
   U69 : OAI21X1 port map( A => n227, B => n188, C => n237, Y => n196);
   U70 : NAND3X1 port map( A => n2, B => n58, C => n226, Y => n237);
   U71 : NOR2X1 port map( A => n26, B => n228, Y => n226);
   U72 : NAND3X1 port map( A => n49, B => n187, C => n179, Y => n228);
   U76 : AOI21X1 port map( A => n236, B => n44, C => RST, Y => n227);
   U77 : OAI21X1 port map( A => n183, B => n25, C => n232, Y => n236);
   U78 : NAND2X1 port map( A => n288, B => n245, Y => n232);
   U79 : NOR2X1 port map( A => D_EDGE, B => n35, Y => n245);
   U81 : OAI21X1 port map( A => n224, B => n185, C => n223, Y => n195);
   U82 : NAND3X1 port map( A => n165, B => n185, C => count_0_port, Y => n223);
   U83 : AOI21X1 port map( A => n222, B => n182, C => n221, Y => n224);
   U84 : OAI21X1 port map( A => n159, B => n186, C => n220, Y => n194);
   U85 : NAND3X1 port map( A => n219, B => n186, C => n160, Y => n220);
   U87 : OAI21X1 port map( A => n217, B => n187, C => n216, Y => n193);
   U88 : NAND3X1 port map( A => n219, B => n187, C => n215, Y => n216);
   U89 : NOR2X1 port map( A => n214, B => n186, Y => n215);
   U90 : AOI21X1 port map( A => n222, B => n186, C => n218, Y => n217);
   U91 : OAI21X1 port map( A => n160, B => n168, C => n274, Y => n218);
   U93 : NAND3X1 port map( A => count_1_port, B => count_0_port, C => n213, Y 
                           => n214);
   U95 : AOI22X1 port map( A => n221, B => count_0_port, C => n182, D => n165, 
                           Y => n212);
   U97 : NAND3X1 port map( A => n219, B => n191, C => SHIFT_ENABLE, Y => n211);
   U100 : OAI21X1 port map( A => n213, B => n168, C => n274, Y => n221);
   U101 : NAND2X1 port map( A => EOP, B => n210, Y => n274);
   U103 : NOR2X1 port map( A => n266, B => n169, Y => n222);
   U104 : NOR2X1 port map( A => n187, B => n225, Y => n266);
   U105 : NAND3X1 port map( A => n185, B => n186, C => n182, Y => n225);
   U110 : NOR2X1 port map( A => BITSTUFF, B => n164, Y => n213);
   U115 : NAND3X1 port map( A => n208, B => n166, C => n248, Y => n284);
   U117 : NAND3X1 port map( A => n207, B => n206, C => n205, Y => n247);
   U119 : NOR2X1 port map( A => RCV_DATA(6), B => RCV_DATA(5), Y => n203);
   U120 : NOR2X1 port map( A => RCV_DATA(4), B => RCV_DATA(3), Y => n204);
   U121 : NOR2X1 port map( A => RCV_DATA(2), B => RCV_DATA(1), Y => n206);
   U122 : NOR2X1 port map( A => RCV_DATA(0), B => n167, Y => n207);
   U124 : NAND3X1 port map( A => n170, B => n261, C => n271, Y => RCVING);
   U125 : NOR2X1 port map( A => n210, B => n202, Y => n271);
   U126 : OAI21X1 port map( A => n24, B => n43, C => n209, Y => n202);
   U127 : NAND3X1 port map( A => n35, B => n44, C => n288, Y => n209);
   U129 : OAI21X1 port map( A => n49, B => n26, C => n283, Y => n201);
   U130 : NAND3X1 port map( A => n35, B => n44, C => n249, Y => n283);
   U131 : NAND3X1 port map( A => n200, B => n199, C => n169, Y => OPCODE_1_port
                           );
   U133 : NAND3X1 port map( A => n23, B => n287, C => n175, Y => n210);
   U135 : NOR2X1 port map( A => n25, B => n24, Y => n268);
   U141 : NOR2X1 port map( A => n44, B => state_2_port, Y => n208);
   U144 : OAI21X1 port map( A => n183, B => n171, C => n44, Y => n199);
   U146 : NOR2X1 port map( A => n174, B => state_0_port, Y => n288);
   U148 : OAI21X1 port map( A => n198, B => n19, C => n49, Y => n200);
   U149 : NOR2X1 port map( A => state_0_port, B => n183, Y => n198);
   U150 : OAI21X1 port map( A => n44, B => n26, C => n261, Y => OPCODE_0_port);
   U151 : NAND3X1 port map( A => n49, B => n35, C => n264, Y => n261);
   U155 : NOR2X1 port map( A => n43, B => n183, Y => n282);
   U3 : OR2X2 port map( A => n297, B => n173, Y => nxtR_ERROR);
   U4 : OR2X2 port map( A => n296, B => n295, Y => nextstate_3_port);
   U14 : AND2X2 port map( A => n284, B => n283, Y => n285);
   U29 : AND2X2 port map( A => n262, B => n261, Y => n263);
   U62 : AND2X2 port map( A => n230, B => n275, Y => n231);
   U63 : OR2X2 port map( A => n24, B => n229, Y => n275);
   U99 : AND2X2 port map( A => n222, B => n274, Y => n219);
   U114 : AND2X2 port map( A => n284, B => n209, Y => n258);
   U118 : AND2X2 port map( A => n204, B => n203, Y => n205);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => CLK, R => 
                           n58, S => n17, Q => state_1_port);
   R_ERROR_reg : DFFSR port map( D => nxtR_ERROR, CLK => CLK, R => n58, S => 
                           n13, Q => R_ERROR);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => CLK, R => 
                           n58, S => n10, Q => state_0_port);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => CLK, R => 
                           n58, S => n8, Q => state_2_port);
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => CLK, R => 
                           n58, S => n7, Q => state_3_port);
   count_reg_0_inst : DFFSR port map( D => n158, CLK => CLK, R => n58, S => n6,
                           Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => n195, CLK => CLK, R => n58, S => n5,
                           Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n194, CLK => CLK, R => n58, S => n4,
                           Q => count_2_port);
   count_reg_3_inst : DFFSR port map( D => n193, CLK => CLK, R => n58, S => n3,
                           Q => count_3_port);
   U10 : AND2X2 port map( A => n183, B => n44, Y => n1);
   U32 : NAND2X1 port map( A => n154, B => n153, Y => n2);
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n10 <= '1';
   n13 <= '1';
   n17 <= '1';
   U73 : INVX2 port map( A => state_3_port, Y => n18);
   U74 : INVX2 port map( A => n18, Y => n19);
   U75 : OR2X2 port map( A => n28, B => n24, Y => n23);
   U80 : INVX2 port map( A => n23, Y => n267);
   U86 : NAND2X1 port map( A => n264, B => n1, Y => n287);
   U92 : INVX2 port map( A => state_2_port, Y => n183);
   U94 : INVX2 port map( A => n25, Y => n264);
   U96 : INVX1 port map( A => n287, Y => n176);
   U98 : OR2X2 port map( A => n44, B => state_2_port, Y => n24);
   U102 : OR2X2 port map( A => n177, B => n19, Y => n25);
   U106 : OR2X2 port map( A => n43, B => n183, Y => n26);
   U107 : OR2X1 port map( A => state_0_port, B => n19, Y => n43);
   U108 : OR2X2 port map( A => n177, B => n174, Y => n28);
   U109 : INVX1 port map( A => n28, Y => n249);
   U111 : INVX2 port map( A => n258, Y => n30);
   U112 : OR2X2 port map( A => n30, B => OPCODE_0_port, Y => W_ENABLE);
   U113 : INVX2 port map( A => RST, Y => n58);
   U116 : INVX1 port map( A => n183, Y => n35);
   U123 : INVX1 port map( A => n43, Y => n248);
   U128 : INVX2 port map( A => state_1_port, Y => n44);
   U132 : INVX1 port map( A => n44, Y => n49);
   U134 : XNOR2X1 port map( A => RX_CHECK_CRC(10), B => RX_CRC(10), Y => n76);
   U136 : XNOR2X1 port map( A => RX_CHECK_CRC(9), B => RX_CRC(9), Y => n73);
   U137 : XOR2X1 port map( A => RX_CHECK_CRC(7), B => RX_CRC(7), Y => n68);
   U138 : XOR2X1 port map( A => RX_CHECK_CRC(8), B => RX_CRC(8), Y => n64);
   U139 : NOR2X1 port map( A => n68, B => n64, Y => n69);
   U140 : NAND3X1 port map( A => n76, B => n73, C => n69, Y => n112);
   U142 : XNOR2X1 port map( A => RX_CHECK_CRC(14), B => RX_CRC(14), Y => n108);
   U143 : XNOR2X1 port map( A => RX_CHECK_CRC(13), B => RX_CRC(13), Y => n104);
   U145 : XOR2X1 port map( A => RX_CHECK_CRC(11), B => RX_CRC(11), Y => n93);
   U147 : XOR2X1 port map( A => RX_CHECK_CRC(12), B => RX_CRC(12), Y => n82);
   U152 : NOR2X1 port map( A => n93, B => n82, Y => n101);
   U153 : NAND3X1 port map( A => n108, B => n104, C => n101, Y => n110);
   U154 : NOR2X1 port map( A => n112, B => n110, Y => n154);
   U156 : NOR2X1 port map( A => n155, B => RX_CHECK_CRC(0), Y => n114);
   U157 : OAI22X1 port map( A => RX_CRC(1), B => n114, C => n114, D => n157, Y 
                           => n131);
   U158 : AND2X1 port map( A => RX_CHECK_CRC(0), B => n155, Y => n115);
   U159 : OAI22X1 port map( A => n115, B => n156, C => RX_CHECK_CRC(1), D => 
                           n115, Y => n130);
   U160 : XOR2X1 port map( A => RX_CHECK_CRC(15), B => RX_CRC(15), Y => n124);
   U161 : XOR2X1 port map( A => RX_CHECK_CRC(2), B => RX_CRC(2), Y => n118);
   U162 : NOR2X1 port map( A => n124, B => n118, Y => n128);
   U163 : NAND3X1 port map( A => n131, B => n130, C => n128, Y => n152);
   U164 : XNOR2X1 port map( A => RX_CHECK_CRC(6), B => RX_CRC(6), Y => n148);
   U165 : XNOR2X1 port map( A => RX_CHECK_CRC(5), B => RX_CRC(5), Y => n143);
   U166 : XOR2X1 port map( A => RX_CHECK_CRC(3), B => RX_CRC(3), Y => n135);
   U167 : XOR2X1 port map( A => RX_CHECK_CRC(4), B => RX_CRC(4), Y => n132);
   U168 : NOR2X1 port map( A => n135, B => n132, Y => n141);
   U169 : NAND3X1 port map( A => n148, B => n143, C => n141, Y => n149);
   U170 : NOR2X1 port map( A => n152, B => n149, Y => n153);
   U171 : INVX2 port map( A => RX_CRC(0), Y => n155);
   U172 : INVX2 port map( A => RX_CRC(1), Y => n156);
   U173 : INVX2 port map( A => RX_CHECK_CRC(1), Y => n157);
   U174 : INVX2 port map( A => n212, Y => n158);
   U175 : INVX2 port map( A => n218, Y => n159);
   U176 : INVX2 port map( A => n214, Y => n160);
   U177 : INVX2 port map( A => SHIFT_ENABLE, Y => n164);
   U178 : INVX2 port map( A => n211, Y => n165);
   U179 : INVX2 port map( A => n247, Y => n166);
   U180 : INVX2 port map( A => RCV_DATA(7), Y => n167);
   U181 : INVX2 port map( A => n222, Y => n168);
   U182 : INVX2 port map( A => n210, Y => n169);
   U183 : INVX2 port map( A => n201, Y => n170);
   U184 : INVX2 port map( A => n288, Y => n171);
   U185 : INVX2 port map( A => n241, Y => n172);
   U186 : INVX2 port map( A => n234, Y => n173);
   U187 : INVX2 port map( A => n19, Y => n174);
   U188 : INVX2 port map( A => n268, Y => n175);
   U189 : INVX2 port map( A => state_0_port, Y => n177);
   U190 : INVX2 port map( A => n228, Y => n178);
   U191 : INVX2 port map( A => n225, Y => n179);
   U192 : INVX2 port map( A => n257, Y => n180);
   U193 : INVX2 port map( A => n266, Y => n181);
   U194 : INVX2 port map( A => count_0_port, Y => n182);
   U195 : INVX2 port map( A => n245, Y => n184);
   U196 : INVX2 port map( A => count_1_port, Y => n185);
   U197 : INVX2 port map( A => count_2_port, Y => n186);
   U198 : INVX2 port map( A => count_3_port, Y => n187);
   U199 : INVX2 port map( A => curCRC_ERROR, Y => n188);
   U200 : INVX2 port map( A => curR_ERROR, Y => n189);
   U201 : INVX2 port map( A => BS_ERROR, Y => n190);
   U202 : INVX2 port map( A => BITSTUFF, Y => n191);
   U203 : INVX2 port map( A => EOP, Y => n192);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_eopdetect_0 is

   port( DP1_RX, DM1_RX : in std_logic;  EOP : out std_logic);

end rx_eopdetect_0;

architecture SYN_Behavioral of rx_eopdetect_0 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;

begin
   
   U1 : NOR2X1 port map( A => DP1_RX, B => DM1_RX, Y => EOP);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_edgedetect_0 is

   port( CLK, RST, DP1_RX : in std_logic;  D_EDGE : out std_logic);

end rx_edgedetect_0;

architecture SYN_Behavioral of rx_edgedetect_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal DP_hold1, DP_hold2, n2, n5, n6, n7 : std_logic;

begin
   
   DP_hold1_reg : DFFSR port map( D => DP1_RX, CLK => CLK, R => n6, S => n2, Q 
                           => DP_hold1);
   DP_hold2_reg : DFFSR port map( D => DP_hold1, CLK => CLK, R => n7, S => n2, 
                           Q => DP_hold2);
   n7 <= '1';
   n6 <= '1';
   U6 : NOR2X1 port map( A => RST, B => n5, Y => D_EDGE);
   U7 : XNOR2X1 port map( A => DP_hold2, B => DP_hold1, Y => n5);
   U4 : INVX2 port map( A => RST, Y => n2);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_decode_0 is

   port( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP : in std_logic;  D_ORIG, BITSTUFF,
         BS_ERROR : out std_logic);

end rx_decode_0;

architecture SYN_moore of rx_decode_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal DP_hold1, DP_hold2, state_3_port, state_2_port, state_1_port, 
      state_0_port, N29, N30, N31, N32, n2, n3, n4, n5, n6, n8, n9, n10, 
      BS_ERROR_port, n12, n13, n14, n15, n16, BITSTUFF_port, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, 
      n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76 : std_logic;

begin
   BITSTUFF <= BITSTUFF_port;
   BS_ERROR <= BS_ERROR_port;
   
   DP_hold2_reg : DFFSR port map( D => n47, CLK => CLK, R => n75, S => n6, Q =>
                           DP_hold2);
   DP_hold1_reg : DFFSR port map( D => n48, CLK => CLK, R => n76, S => n6, Q =>
                           DP_hold1);
   n76 <= '1';
   n75 <= '1';
   U10 : OR2X2 port map( A => n8, B => state_1_port, Y => n55);
   U20 : NAND2X1 port map( A => n74, B => n73, Y => n48);
   U21 : AOI22X1 port map( A => DP_hold1, B => n12, C => DP1_RX, D => n72, Y =>
                           n74);
   U22 : NAND2X1 port map( A => n71, B => n73, Y => n47);
   U23 : AOI22X1 port map( A => n10, B => DP_hold1, C => DP_hold2, D => n70, Y 
                           => n71);
   U24 : NAND2X1 port map( A => SHIFT_ENABLE, B => n72, Y => n70);
   U25 : XNOR2X1 port map( A => DP_hold1, B => DP_hold2, Y => D_ORIG);
   U26 : NOR2X1 port map( A => n69, B => EOP, Y => N32);
   U27 : AOI21X1 port map( A => n68, B => BITSTUFF_port, C => BS_ERROR_port, Y 
                           => n69);
   U28 : NAND3X1 port map( A => state_3_port, B => n16, C => n66, Y => n67);
   U29 : NOR2X1 port map( A => state_2_port, B => state_1_port, Y => n66);
   U30 : NOR2X1 port map( A => n72, B => state_3_port, Y => BITSTUFF_port);
   U31 : NOR2X1 port map( A => n65, B => n14, Y => N31);
   U32 : AOI21X1 port map( A => state_2_port, B => n64, C => n63, Y => n65);
   U33 : OAI21X1 port map( A => n62, B => n61, C => n60, Y => n63);
   U34 : NAND2X1 port map( A => state_0_port, B => n68, Y => n61);
   U35 : NAND2X1 port map( A => state_1_port, B => n15, Y => n62);
   U36 : OAI21X1 port map( A => state_1_port, B => n59, C => SHIFT_ENABLE, Y =>
                           n64);
   U37 : NOR2X1 port map( A => n58, B => n14, Y => N30);
   U38 : AOI21X1 port map( A => state_1_port, B => n57, C => n56, Y => n58);
   U39 : OAI21X1 port map( A => n16, B => n55, C => n60, Y => n56);
   U40 : NAND2X1 port map( A => n12, B => n59, Y => n60);
   U41 : NAND2X1 port map( A => n13, B => n16, Y => n72);
   U42 : OAI21X1 port map( A => n59, B => n54, C => SHIFT_ENABLE, Y => n57);
   U43 : NAND2X1 port map( A => n16, B => n15, Y => n54);
   U44 : NOR2X1 port map( A => n53, B => n14, Y => N29);
   U45 : NOR2X1 port map( A => EOP, B => state_3_port, Y => n73);
   U46 : AOI21X1 port map( A => state_0_port, B => n9, C => n52, Y => n53);
   U47 : OAI21X1 port map( A => n8, B => n51, C => n50, Y => n52);
   U48 : NAND3X1 port map( A => n13, B => n59, C => SHIFT_ENABLE, Y => n50);
   U49 : NAND2X1 port map( A => n49, B => n16, Y => n51);
   U50 : NAND2X1 port map( A => state_2_port, B => state_1_port, Y => n49);
   U51 : NOR2X1 port map( A => n59, B => n9, Y => n68);
   U52 : XOR2X1 port map( A => DP1_RX, B => DP_hold2, Y => n59);
   state_reg_3_inst : DFFSR port map( D => N32, CLK => CLK, R => n6, S => n5, Q
                           => state_3_port);
   state_reg_0_inst : DFFSR port map( D => N29, CLK => CLK, R => n6, S => n4, Q
                           => state_0_port);
   state_reg_2_inst : DFFSR port map( D => N31, CLK => CLK, R => n6, S => n3, Q
                           => state_2_port);
   state_reg_1_inst : DFFSR port map( D => N30, CLK => CLK, R => n6, S => n2, Q
                           => state_1_port);
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   U8 : INVX2 port map( A => RST, Y => n6);
   U11 : INVX2 port map( A => n68, Y => n8);
   U12 : INVX2 port map( A => SHIFT_ENABLE, Y => n9);
   U13 : INVX2 port map( A => n70, Y => n10);
   U14 : INVX2 port map( A => n67, Y => BS_ERROR_port);
   U15 : INVX2 port map( A => n72, Y => n12);
   U16 : INVX2 port map( A => n49, Y => n13);
   U17 : INVX2 port map( A => n73, Y => n14);
   U18 : INVX2 port map( A => state_2_port, Y => n15);
   U19 : INVX2 port map( A => state_0_port, Y => n16);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_accumulator_0 is

   port( CLK, RST : in std_logic;  RCV_DATA : in std_logic_vector (7 downto 0);
         W_ENABLE : in std_logic;  rx_CHECK_CRC : out std_logic_vector (15 
         downto 0));

end rx_accumulator_0;

architecture SYN_Behavioral of rx_accumulator_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, rx_CHECK_CRC_13_port, 
      rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, rx_CHECK_CRC_10_port, 
      rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, rx_CHECK_CRC_7_port, 
      rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, rx_CHECK_CRC_4_port, 
      rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, rx_CHECK_CRC_1_port, 
      rx_CHECK_CRC_0_port, n1, n2, n5, n8, n11, n14, n17, n20, n23, n26, n28, 
      n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n57
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91 : std_logic;

begin
   rx_CHECK_CRC <= ( rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, 
      rx_CHECK_CRC_13_port, rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, 
      rx_CHECK_CRC_10_port, rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, 
      rx_CHECK_CRC_7_port, rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, 
      rx_CHECK_CRC_4_port, rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, 
      rx_CHECK_CRC_1_port, rx_CHECK_CRC_0_port );
   
   U2 : OAI21X1 port map( A => n40, B => n59, C => n91, Y => n75);
   U3 : NAND2X1 port map( A => rx_CHECK_CRC_8_port, B => n40, Y => n91);
   U4 : OAI21X1 port map( A => n42, B => n59, C => n90, Y => n74);
   U5 : NAND2X1 port map( A => RCV_DATA(0), B => n42, Y => n90);
   U7 : OAI21X1 port map( A => n40, B => n57, C => n89, Y => n73);
   U8 : NAND2X1 port map( A => rx_CHECK_CRC_9_port, B => n40, Y => n89);
   U9 : OAI21X1 port map( A => n42, B => n57, C => n88, Y => n72);
   U10 : NAND2X1 port map( A => RCV_DATA(1), B => n42, Y => n88);
   U12 : OAI21X1 port map( A => n40, B => n56, C => n87, Y => n71);
   U13 : NAND2X1 port map( A => rx_CHECK_CRC_10_port, B => n40, Y => n87);
   U14 : OAI21X1 port map( A => n42, B => n56, C => n86, Y => n70);
   U15 : NAND2X1 port map( A => RCV_DATA(2), B => n42, Y => n86);
   U17 : OAI21X1 port map( A => n40, B => n54, C => n85, Y => n69);
   U18 : NAND2X1 port map( A => rx_CHECK_CRC_11_port, B => n40, Y => n85);
   U19 : OAI21X1 port map( A => n42, B => n54, C => n84, Y => n68);
   U20 : NAND2X1 port map( A => RCV_DATA(3), B => n42, Y => n84);
   U22 : OAI21X1 port map( A => n40, B => n52, C => n83, Y => n67);
   U23 : NAND2X1 port map( A => rx_CHECK_CRC_12_port, B => n40, Y => n83);
   U24 : OAI21X1 port map( A => n42, B => n52, C => n82, Y => n66);
   U25 : NAND2X1 port map( A => RCV_DATA(4), B => n42, Y => n82);
   U27 : OAI21X1 port map( A => n40, B => n50, C => n81, Y => n65);
   U28 : NAND2X1 port map( A => rx_CHECK_CRC_13_port, B => n40, Y => n81);
   U29 : OAI21X1 port map( A => n42, B => n50, C => n80, Y => n64);
   U30 : NAND2X1 port map( A => RCV_DATA(5), B => n42, Y => n80);
   U32 : OAI21X1 port map( A => n40, B => n48, C => n79, Y => n63);
   U33 : NAND2X1 port map( A => rx_CHECK_CRC_14_port, B => n40, Y => n79);
   U34 : OAI21X1 port map( A => n42, B => n48, C => n78, Y => n62);
   U35 : NAND2X1 port map( A => RCV_DATA(6), B => n42, Y => n78);
   U37 : OAI21X1 port map( A => n40, B => n46, C => n77, Y => n61);
   U38 : NAND2X1 port map( A => rx_CHECK_CRC_15_port, B => n40, Y => n77);
   U41 : OAI21X1 port map( A => n42, B => n46, C => n76, Y => n60);
   U42 : NAND2X1 port map( A => RCV_DATA(7), B => n42, Y => n76);
   present_CHECK_CRC_reg_7_inst : DFFSR port map( D => n60, CLK => CLK, R => 
                           n44, S => n38, Q => rx_CHECK_CRC_7_port);
   present_CHECK_CRC_reg_6_inst : DFFSR port map( D => n62, CLK => CLK, R => 
                           n44, S => n36, Q => rx_CHECK_CRC_6_port);
   present_CHECK_CRC_reg_5_inst : DFFSR port map( D => n64, CLK => CLK, R => 
                           n44, S => n34, Q => rx_CHECK_CRC_5_port);
   present_CHECK_CRC_reg_4_inst : DFFSR port map( D => n66, CLK => CLK, R => 
                           n44, S => n32, Q => rx_CHECK_CRC_4_port);
   present_CHECK_CRC_reg_3_inst : DFFSR port map( D => n68, CLK => CLK, R => 
                           n44, S => n30, Q => rx_CHECK_CRC_3_port);
   present_CHECK_CRC_reg_2_inst : DFFSR port map( D => n70, CLK => CLK, R => 
                           n44, S => n28, Q => rx_CHECK_CRC_2_port);
   present_CHECK_CRC_reg_1_inst : DFFSR port map( D => n72, CLK => CLK, R => 
                           n44, S => n26, Q => rx_CHECK_CRC_1_port);
   present_CHECK_CRC_reg_0_inst : DFFSR port map( D => n74, CLK => CLK, R => 
                           n44, S => n23, Q => rx_CHECK_CRC_0_port);
   present_CHECK_CRC_reg_15_inst : DFFSR port map( D => n61, CLK => CLK, R => 
                           n44, S => n20, Q => rx_CHECK_CRC_15_port);
   present_CHECK_CRC_reg_14_inst : DFFSR port map( D => n63, CLK => CLK, R => 
                           n44, S => n17, Q => rx_CHECK_CRC_14_port);
   present_CHECK_CRC_reg_13_inst : DFFSR port map( D => n65, CLK => CLK, R => 
                           n44, S => n14, Q => rx_CHECK_CRC_13_port);
   present_CHECK_CRC_reg_12_inst : DFFSR port map( D => n67, CLK => CLK, R => 
                           n44, S => n11, Q => rx_CHECK_CRC_12_port);
   present_CHECK_CRC_reg_11_inst : DFFSR port map( D => n69, CLK => CLK, R => 
                           n44, S => n8, Q => rx_CHECK_CRC_11_port);
   present_CHECK_CRC_reg_10_inst : DFFSR port map( D => n71, CLK => CLK, R => 
                           n44, S => n5, Q => rx_CHECK_CRC_10_port);
   present_CHECK_CRC_reg_9_inst : DFFSR port map( D => n73, CLK => CLK, R => 
                           n44, S => n2, Q => rx_CHECK_CRC_9_port);
   present_CHECK_CRC_reg_8_inst : DFFSR port map( D => n75, CLK => CLK, R => 
                           n44, S => n1, Q => rx_CHECK_CRC_8_port);
   n1 <= '1';
   n2 <= '1';
   n5 <= '1';
   n8 <= '1';
   n11 <= '1';
   n14 <= '1';
   n17 <= '1';
   n20 <= '1';
   n23 <= '1';
   n26 <= '1';
   n28 <= '1';
   n30 <= '1';
   n32 <= '1';
   n34 <= '1';
   n36 <= '1';
   n38 <= '1';
   U50 : INVX2 port map( A => n40, Y => n42);
   U51 : INVX2 port map( A => W_ENABLE, Y => n40);
   U52 : INVX2 port map( A => RST, Y => n44);
   U53 : INVX2 port map( A => rx_CHECK_CRC_7_port, Y => n46);
   U54 : INVX2 port map( A => rx_CHECK_CRC_6_port, Y => n48);
   U55 : INVX2 port map( A => rx_CHECK_CRC_5_port, Y => n50);
   U56 : INVX2 port map( A => rx_CHECK_CRC_4_port, Y => n52);
   U57 : INVX2 port map( A => rx_CHECK_CRC_3_port, Y => n54);
   U58 : INVX2 port map( A => rx_CHECK_CRC_2_port, Y => n56);
   U59 : INVX2 port map( A => rx_CHECK_CRC_1_port, Y => n57);
   U60 : INVX2 port map( A => rx_CHECK_CRC_0_port, Y => n59);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_CRC_CALC_0 is

   port( CLK, RST, W_ENABLE : in std_logic;  OPCODE : in std_logic_vector (1 
         downto 0);  RCV_DATA : in std_logic_vector (7 downto 0);  RX_CRC : out
         std_logic_vector (15 downto 0));

end rx_CRC_CALC_0;

architecture SYN_moore of rx_CRC_CALC_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port, current_crc_15_port, 
      current_crc_14_port, current_crc_13_port, current_crc_12_port, 
      current_crc_11_port, current_crc_10_port, current_crc_9_port, 
      current_crc_8_port, current_crc_7_port, current_crc_6_port, 
      current_crc_5_port, current_crc_4_port, current_crc_3_port, 
      current_crc_2_port, current_crc_1_port, current_crc_0_port, 
      cache_1_15_port, cache_1_14_port, cache_1_13_port, cache_1_12_port, 
      cache_1_11_port, cache_1_10_port, cache_1_9_port, cache_1_8_port, 
      cache_1_7_port, cache_1_6_port, cache_1_5_port, cache_1_4_port, 
      cache_1_3_port, cache_1_2_port, cache_1_1_port, cache_1_0_port, n1, n2, 
      n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48
      , n49, n50, n56, n60, n79, n80, n81, n82, n100, n102, n104, n106, n108, 
      n110, n112, n114, n116, n118, n120, n122, n124, n126, n128, n130, n131, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246 : std_logic;

begin
   RX_CRC <= ( RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port );
   
   cache_1_reg_0_inst : DFFPOSX1 port map( D => n173, CLK => CLK, Q => 
                           cache_1_0_port);
   cache_1_reg_8_inst : DFFPOSX1 port map( D => n174, CLK => CLK, Q => 
                           cache_1_8_port);
   cache_1_reg_15_inst : DFFPOSX1 port map( D => n175, CLK => CLK, Q => 
                           cache_1_15_port);
   cache_1_reg_1_inst : DFFPOSX1 port map( D => n176, CLK => CLK, Q => 
                           cache_1_1_port);
   cache_1_reg_9_inst : DFFPOSX1 port map( D => n177, CLK => CLK, Q => 
                           cache_1_9_port);
   cache_1_reg_2_inst : DFFPOSX1 port map( D => n178, CLK => CLK, Q => 
                           cache_1_2_port);
   cache_1_reg_10_inst : DFFPOSX1 port map( D => n179, CLK => CLK, Q => 
                           cache_1_10_port);
   cache_1_reg_3_inst : DFFPOSX1 port map( D => n180, CLK => CLK, Q => 
                           cache_1_3_port);
   cache_1_reg_11_inst : DFFPOSX1 port map( D => n181, CLK => CLK, Q => 
                           cache_1_11_port);
   cache_1_reg_4_inst : DFFPOSX1 port map( D => n182, CLK => CLK, Q => 
                           cache_1_4_port);
   cache_1_reg_12_inst : DFFPOSX1 port map( D => n183, CLK => CLK, Q => 
                           cache_1_12_port);
   cache_1_reg_5_inst : DFFPOSX1 port map( D => n184, CLK => CLK, Q => 
                           cache_1_5_port);
   cache_1_reg_13_inst : DFFPOSX1 port map( D => n185, CLK => CLK, Q => 
                           cache_1_13_port);
   cache_1_reg_6_inst : DFFPOSX1 port map( D => n186, CLK => CLK, Q => 
                           cache_1_6_port);
   cache_1_reg_14_inst : DFFPOSX1 port map( D => n187, CLK => CLK, Q => 
                           cache_1_14_port);
   cache_1_reg_7_inst : DFFPOSX1 port map( D => n188, CLK => CLK, Q => 
                           cache_1_7_port);
   cache_2_reg_15_inst : DFFPOSX1 port map( D => n189, CLK => CLK, Q => 
                           RX_CRC_15_port);
   cache_2_reg_14_inst : DFFPOSX1 port map( D => n190, CLK => CLK, Q => 
                           RX_CRC_14_port);
   cache_2_reg_13_inst : DFFPOSX1 port map( D => n191, CLK => CLK, Q => 
                           RX_CRC_13_port);
   cache_2_reg_12_inst : DFFPOSX1 port map( D => n192, CLK => CLK, Q => 
                           RX_CRC_12_port);
   cache_2_reg_11_inst : DFFPOSX1 port map( D => n193, CLK => CLK, Q => 
                           RX_CRC_11_port);
   cache_2_reg_10_inst : DFFPOSX1 port map( D => n194, CLK => CLK, Q => 
                           RX_CRC_10_port);
   cache_2_reg_9_inst : DFFPOSX1 port map( D => n195, CLK => CLK, Q => 
                           RX_CRC_9_port);
   cache_2_reg_8_inst : DFFPOSX1 port map( D => n196, CLK => CLK, Q => 
                           RX_CRC_8_port);
   cache_2_reg_7_inst : DFFPOSX1 port map( D => n197, CLK => CLK, Q => 
                           RX_CRC_7_port);
   cache_2_reg_6_inst : DFFPOSX1 port map( D => n198, CLK => CLK, Q => 
                           RX_CRC_6_port);
   cache_2_reg_5_inst : DFFPOSX1 port map( D => n199, CLK => CLK, Q => 
                           RX_CRC_5_port);
   cache_2_reg_4_inst : DFFPOSX1 port map( D => n200, CLK => CLK, Q => 
                           RX_CRC_4_port);
   cache_2_reg_3_inst : DFFPOSX1 port map( D => n201, CLK => CLK, Q => 
                           RX_CRC_3_port);
   cache_2_reg_2_inst : DFFPOSX1 port map( D => n202, CLK => CLK, Q => 
                           RX_CRC_2_port);
   cache_2_reg_1_inst : DFFPOSX1 port map( D => n203, CLK => CLK, Q => 
                           RX_CRC_1_port);
   cache_2_reg_0_inst : DFFPOSX1 port map( D => n204, CLK => CLK, Q => 
                           RX_CRC_0_port);
   U3 : OAI21X1 port map( A => n42, B => n60, C => n246, Y => n204);
   U4 : NAND2X1 port map( A => RX_CRC_0_port, B => n43, Y => n246);
   U5 : OAI21X1 port map( A => n41, B => n102, C => n245, Y => n203);
   U6 : NAND2X1 port map( A => RX_CRC_1_port, B => n43, Y => n245);
   U7 : OAI21X1 port map( A => n41, B => n110, C => n244, Y => n202);
   U8 : NAND2X1 port map( A => RX_CRC_2_port, B => n43, Y => n244);
   U9 : OAI21X1 port map( A => n41, B => n118, C => n243, Y => n201);
   U10 : NAND2X1 port map( A => RX_CRC_3_port, B => n43, Y => n243);
   U11 : OAI21X1 port map( A => n41, B => n126, C => n242, Y => n200);
   U12 : NAND2X1 port map( A => RX_CRC_4_port, B => n43, Y => n242);
   U13 : OAI21X1 port map( A => n41, B => n148, C => n241, Y => n199);
   U14 : NAND2X1 port map( A => RX_CRC_5_port, B => n42, Y => n241);
   U15 : OAI21X1 port map( A => n41, B => n152, C => n240, Y => n198);
   U16 : NAND2X1 port map( A => RX_CRC_6_port, B => n42, Y => n240);
   U17 : OAI21X1 port map( A => n41, B => n156, C => n239, Y => n197);
   U18 : NAND2X1 port map( A => RX_CRC_7_port, B => n42, Y => n239);
   U19 : OAI21X1 port map( A => n41, B => n80, C => n238, Y => n196);
   U20 : NAND2X1 port map( A => RX_CRC_8_port, B => n42, Y => n238);
   U21 : OAI21X1 port map( A => n41, B => n106, C => n237, Y => n195);
   U22 : NAND2X1 port map( A => RX_CRC_9_port, B => n42, Y => n237);
   U23 : OAI21X1 port map( A => n42, B => n114, C => n236, Y => n194);
   U24 : NAND2X1 port map( A => RX_CRC_10_port, B => n42, Y => n236);
   U25 : OAI21X1 port map( A => n42, B => n122, C => n235, Y => n193);
   U26 : NAND2X1 port map( A => RX_CRC_11_port, B => n42, Y => n235);
   U27 : OAI21X1 port map( A => n42, B => n130, C => n234, Y => n192);
   U28 : NAND2X1 port map( A => RX_CRC_12_port, B => n42, Y => n234);
   U29 : OAI21X1 port map( A => n42, B => n150, C => n233, Y => n191);
   U30 : NAND2X1 port map( A => RX_CRC_13_port, B => n43, Y => n233);
   U31 : OAI21X1 port map( A => n42, B => n154, C => n232, Y => n190);
   U32 : NAND2X1 port map( A => RX_CRC_14_port, B => n43, Y => n232);
   U33 : OAI21X1 port map( A => n42, B => n82, C => n231, Y => n189);
   U34 : NAND2X1 port map( A => RX_CRC_15_port, B => n43, Y => n231);
   U35 : OAI22X1 port map( A => n41, B => n155, C => n39, D => n156, Y => n188)
                           ;
   U37 : OAI22X1 port map( A => n41, B => n153, C => n39, D => n154, Y => n187)
                           ;
   U39 : OAI22X1 port map( A => n41, B => n151, C => n39, D => n152, Y => n186)
                           ;
   U41 : OAI22X1 port map( A => n41, B => n149, C => n39, D => n150, Y => n185)
                           ;
   U43 : OAI22X1 port map( A => n40, B => n131, C => n39, D => n148, Y => n184)
                           ;
   U45 : OAI22X1 port map( A => n40, B => n128, C => n39, D => n130, Y => n183)
                           ;
   U47 : OAI22X1 port map( A => n40, B => n124, C => n39, D => n126, Y => n182)
                           ;
   U49 : OAI22X1 port map( A => n40, B => n120, C => n39, D => n122, Y => n181)
                           ;
   U51 : OAI22X1 port map( A => n40, B => n116, C => n39, D => n118, Y => n180)
                           ;
   U53 : OAI22X1 port map( A => n40, B => n112, C => n38, D => n114, Y => n179)
                           ;
   U55 : OAI22X1 port map( A => n40, B => n108, C => n38, D => n110, Y => n178)
                           ;
   U57 : OAI22X1 port map( A => n40, B => n104, C => n38, D => n106, Y => n177)
                           ;
   U59 : OAI22X1 port map( A => n40, B => n100, C => n38, D => n102, Y => n176)
                           ;
   U61 : OAI22X1 port map( A => n40, B => n81, C => n38, D => n82, Y => n175);
   U63 : OAI22X1 port map( A => n40, B => n79, C => n38, D => n80, Y => n174);
   U65 : OAI22X1 port map( A => n40, B => n56, C => n38, D => n60, Y => n173);
   U70 : OAI22X1 port map( A => n81, B => n37, C => n228, D => n35, Y => n172);
   U71 : XOR2X1 port map( A => n227, B => current_crc_7_port, Y => n228);
   U72 : OAI22X1 port map( A => n35, B => n151, C => n153, D => n37, Y => n171)
                           ;
   U73 : OAI22X1 port map( A => n35, B => n131, C => n149, D => n229, Y => n170
                           );
   U74 : OAI22X1 port map( A => n230, B => n124, C => n128, D => n37, Y => n169
                           );
   U75 : OAI22X1 port map( A => n35, B => n116, C => n120, D => n229, Y => n168
                           );
   U77 : OAI22X1 port map( A => n230, B => n108, C => n112, D => n37, Y => n167
                           );
   U78 : OAI22X1 port map( A => n104, B => n37, C => n226, D => n230, Y => n166
                           );
   U79 : XOR2X1 port map( A => n100, B => n45, Y => n226);
   U80 : OAI22X1 port map( A => n79, B => n229, C => n225, D => n35, Y => n165)
                           ;
   U81 : XOR2X1 port map( A => n224, B => n223, Y => n225);
   U82 : XOR2X1 port map( A => n56, B => n45, Y => n224);
   U84 : OAI22X1 port map( A => n155, B => n37, C => n46, D => n230, Y => n164)
                           ;
   U86 : OAI22X1 port map( A => n151, B => n229, C => n222, D => n35, Y => n163
                           );
   U87 : XOR2X1 port map( A => n221, B => n220, Y => n222);
   U89 : OAI22X1 port map( A => n131, B => n37, C => n219, D => n230, Y => n162
                           );
   U91 : OAI22X1 port map( A => n124, B => n229, C => n218, D => n35, Y => n161
                           );
   U92 : XOR2X1 port map( A => n217, B => n216, Y => n218);
   U94 : OAI22X1 port map( A => n116, B => n37, C => n215, D => n230, Y => n160
                           );
   U96 : OAI22X1 port map( A => n108, B => n229, C => n214, D => n35, Y => n159
                           );
   U97 : XOR2X1 port map( A => n213, B => n212, Y => n214);
   U99 : OAI22X1 port map( A => n100, B => n37, C => n211, D => n230, Y => n158
                           );
   U100 : XOR2X1 port map( A => n210, B => n209, Y => n211);
   U101 : XOR2X1 port map( A => n208, B => n207, Y => n210);
   U103 : OAI22X1 port map( A => n56, B => n229, C => n227, D => n35, Y => n157
                           );
   U104 : XOR2X1 port map( A => n206, B => n205, Y => n227);
   U105 : XOR2X1 port map( A => n45, B => n212, Y => n205);
   U106 : XOR2X1 port map( A => current_crc_8_port, B => RCV_DATA(0), Y => n212
                           );
   U108 : XOR2X1 port map( A => n81, B => RCV_DATA(7), Y => n208);
   U110 : XOR2X1 port map( A => n46, B => n207, Y => n206);
   U111 : XOR2X1 port map( A => n215, B => n219, Y => n207);
   U112 : XNOR2X1 port map( A => n220, B => n216, Y => n219);
   U113 : XOR2X1 port map( A => current_crc_11_port, B => RCV_DATA(3), Y => 
                           n216);
   U114 : XNOR2X1 port map( A => n128, B => RCV_DATA(4), Y => n220);
   U116 : XOR2X1 port map( A => n213, B => n48, Y => n215);
   U118 : XOR2X1 port map( A => n112, B => RCV_DATA(2), Y => n217);
   U120 : XOR2X1 port map( A => n104, B => RCV_DATA(1), Y => n213);
   U123 : XOR2X1 port map( A => n223, B => n47, Y => n209);
   U125 : XOR2X1 port map( A => n149, B => RCV_DATA(5), Y => n221);
   U127 : XNOR2X1 port map( A => n153, B => RCV_DATA(6), Y => n223);
   U129 : OAI21X1 port map( A => n50, B => n49, C => n230, Y => n229);
   U130 : NAND3X1 port map( A => OPCODE(0), B => n49, C => W_ENABLE, Y => n230)
                           ;
   current_crc_reg_14_inst : DFFSR port map( D => n171, CLK => CLK, R => n44, S
                           => n30, Q => current_crc_14_port);
   current_crc_reg_12_inst : DFFSR port map( D => n169, CLK => CLK, R => n44, S
                           => n28, Q => current_crc_12_port);
   current_crc_reg_10_inst : DFFSR port map( D => n167, CLK => CLK, R => n44, S
                           => n26, Q => current_crc_10_port);
   current_crc_reg_13_inst : DFFSR port map( D => n170, CLK => CLK, R => n44, S
                           => n24, Q => current_crc_13_port);
   current_crc_reg_11_inst : DFFSR port map( D => n168, CLK => CLK, R => n44, S
                           => n22, Q => current_crc_11_port);
   current_crc_reg_15_inst : DFFSR port map( D => n172, CLK => CLK, R => n44, S
                           => n20, Q => current_crc_15_port);
   current_crc_reg_8_inst : DFFSR port map( D => n165, CLK => CLK, R => n44, S 
                           => n18, Q => current_crc_8_port);
   current_crc_reg_6_inst : DFFSR port map( D => n163, CLK => CLK, R => n44, S 
                           => n16, Q => current_crc_6_port);
   current_crc_reg_4_inst : DFFSR port map( D => n161, CLK => CLK, R => n44, S 
                           => n14, Q => current_crc_4_port);
   current_crc_reg_2_inst : DFFSR port map( D => n159, CLK => CLK, R => n44, S 
                           => n12, Q => current_crc_2_port);
   current_crc_reg_0_inst : DFFSR port map( D => n157, CLK => CLK, R => n44, S 
                           => n10, Q => current_crc_0_port);
   current_crc_reg_9_inst : DFFSR port map( D => n166, CLK => CLK, R => n44, S 
                           => n8, Q => current_crc_9_port);
   current_crc_reg_7_inst : DFFSR port map( D => n164, CLK => CLK, R => n44, S 
                           => n6, Q => current_crc_7_port);
   current_crc_reg_5_inst : DFFSR port map( D => n162, CLK => CLK, R => n44, S 
                           => n4, Q => current_crc_5_port);
   current_crc_reg_3_inst : DFFSR port map( D => n160, CLK => CLK, R => n44, S 
                           => n2, Q => current_crc_3_port);
   current_crc_reg_1_inst : DFFSR port map( D => n158, CLK => CLK, R => n44, S 
                           => n1, Q => current_crc_1_port);
   U36 : INVX2 port map( A => n32, Y => n38);
   n1 <= '1';
   n2 <= '1';
   n4 <= '1';
   n6 <= '1';
   n8 <= '1';
   n10 <= '1';
   n12 <= '1';
   n14 <= '1';
   n16 <= '1';
   n18 <= '1';
   n20 <= '1';
   n22 <= '1';
   n24 <= '1';
   n26 <= '1';
   n28 <= '1';
   n30 <= '1';
   U68 : INVX2 port map( A => n230, Y => n34);
   U69 : BUFX2 port map( A => n32, Y => n43);
   U76 : INVX2 port map( A => n32, Y => n39);
   U83 : OR2X2 port map( A => n35, B => RST, Y => n32);
   U85 : INVX2 port map( A => n34, Y => n35);
   U88 : INVX2 port map( A => n36, Y => n37);
   U90 : INVX2 port map( A => n229, Y => n36);
   U93 : INVX2 port map( A => RST, Y => n44);
   U95 : INVX1 port map( A => OPCODE(0), Y => n50);
   U98 : INVX1 port map( A => OPCODE(1), Y => n49);
   U102 : BUFX4 port map( A => n32, Y => n40);
   U107 : BUFX4 port map( A => n32, Y => n41);
   U109 : BUFX4 port map( A => n32, Y => n42);
   U115 : INVX2 port map( A => n208, Y => n45);
   U117 : INVX2 port map( A => n209, Y => n46);
   U119 : INVX2 port map( A => n221, Y => n47);
   U121 : INVX2 port map( A => n217, Y => n48);
   U122 : INVX2 port map( A => current_crc_0_port, Y => n56);
   U124 : INVX2 port map( A => cache_1_0_port, Y => n60);
   U126 : INVX2 port map( A => current_crc_8_port, Y => n79);
   U128 : INVX2 port map( A => cache_1_8_port, Y => n80);
   U131 : INVX2 port map( A => current_crc_15_port, Y => n81);
   U132 : INVX2 port map( A => cache_1_15_port, Y => n82);
   U133 : INVX2 port map( A => current_crc_1_port, Y => n100);
   U134 : INVX2 port map( A => cache_1_1_port, Y => n102);
   U135 : INVX2 port map( A => current_crc_9_port, Y => n104);
   U136 : INVX2 port map( A => cache_1_9_port, Y => n106);
   U137 : INVX2 port map( A => current_crc_2_port, Y => n108);
   U138 : INVX2 port map( A => cache_1_2_port, Y => n110);
   U139 : INVX2 port map( A => current_crc_10_port, Y => n112);
   U140 : INVX2 port map( A => cache_1_10_port, Y => n114);
   U141 : INVX2 port map( A => current_crc_3_port, Y => n116);
   U142 : INVX2 port map( A => cache_1_3_port, Y => n118);
   U143 : INVX2 port map( A => current_crc_11_port, Y => n120);
   U144 : INVX2 port map( A => cache_1_11_port, Y => n122);
   U145 : INVX2 port map( A => current_crc_4_port, Y => n124);
   U146 : INVX2 port map( A => cache_1_4_port, Y => n126);
   U147 : INVX2 port map( A => current_crc_12_port, Y => n128);
   U148 : INVX2 port map( A => cache_1_12_port, Y => n130);
   U149 : INVX2 port map( A => current_crc_5_port, Y => n131);
   U150 : INVX2 port map( A => cache_1_5_port, Y => n148);
   U151 : INVX2 port map( A => current_crc_13_port, Y => n149);
   U152 : INVX2 port map( A => cache_1_13_port, Y => n150);
   U153 : INVX2 port map( A => current_crc_6_port, Y => n151);
   U154 : INVX2 port map( A => cache_1_6_port, Y => n152);
   U155 : INVX2 port map( A => current_crc_14_port, Y => n153);
   U156 : INVX2 port map( A => cache_1_14_port, Y => n154);
   U157 : INVX2 port map( A => current_crc_7_port, Y => n155);
   U158 : INVX2 port map( A => cache_1_7_port, Y => n156);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RFIFO_0 is

   port( CLK, RST, W_ENABLE, R_ENABLE : in std_logic;  RCV_DATA : in 
         std_logic_vector (7 downto 0);  RCV_OPCODE : in std_logic_vector (1 
         downto 0);  DATA : out std_logic_vector (7 downto 0);  OUT_OPCODE : 
         out std_logic_vector (1 downto 0);  BYTE_COUNT : out std_logic_vector 
         (4 downto 0);  EMPTY, FULL : out std_logic);

end RFIFO_0;

architecture SYN_BRFIFO of RFIFO_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, 
      DATA_3_port, DATA_2_port, DATA_1_port, DATA_0_port, OUT_OPCODE_1_port, 
      OUT_OPCODE_0_port, EMPTY_port, FULL_port, readptr_4_port, readptr_3_port,
      readptr_2_port, readptr_1_port, readptr_0_port, writeptr_4_port, 
      writeptr_3_port, writeptr_2_port, writeptr_1_port, writeptr_0_port, state
      , N32, N33, N34, N43, N44, N45, N46, opcode_0_1_port, opcode_0_0_port, 
      opcode_1_1_port, opcode_1_0_port, opcode_2_1_port, opcode_2_0_port, 
      opcode_3_1_port, opcode_3_0_port, opcode_4_1_port, opcode_4_0_port, 
      opcode_5_1_port, opcode_5_0_port, opcode_6_1_port, opcode_6_0_port, 
      opcode_7_1_port, opcode_7_0_port, opcode_8_1_port, opcode_8_0_port, 
      opcode_9_1_port, opcode_9_0_port, opcode_10_1_port, opcode_10_0_port, 
      opcode_11_1_port, opcode_11_0_port, opcode_12_1_port, opcode_12_0_port, 
      opcode_13_1_port, opcode_13_0_port, opcode_14_1_port, opcode_14_0_port, 
      opcode_15_1_port, opcode_15_0_port, opcode_16_1_port, opcode_16_0_port, 
      opcode_17_1_port, opcode_17_0_port, opcode_18_1_port, opcode_18_0_port, 
      opcode_19_1_port, opcode_19_0_port, opcode_20_1_port, opcode_20_0_port, 
      opcode_21_1_port, opcode_21_0_port, opcode_22_1_port, opcode_22_0_port, 
      opcode_23_1_port, opcode_23_0_port, opcode_24_1_port, opcode_24_0_port, 
      opcode_25_1_port, opcode_25_0_port, opcode_26_1_port, opcode_26_0_port, 
      opcode_27_1_port, opcode_27_0_port, opcode_28_1_port, opcode_28_0_port, 
      opcode_29_1_port, opcode_29_0_port, opcode_30_1_port, opcode_30_0_port, 
      opcode_31_1_port, opcode_31_0_port, memory_0_7_port, memory_0_6_port, 
      memory_0_5_port, memory_0_4_port, memory_0_3_port, memory_0_2_port, 
      memory_0_1_port, memory_0_0_port, memory_1_7_port, memory_1_6_port, 
      memory_1_5_port, memory_1_4_port, memory_1_3_port, memory_1_2_port, 
      memory_1_1_port, memory_1_0_port, memory_2_7_port, memory_2_6_port, 
      memory_2_5_port, memory_2_4_port, memory_2_3_port, memory_2_2_port, 
      memory_2_1_port, memory_2_0_port, memory_3_7_port, memory_3_6_port, 
      memory_3_5_port, memory_3_4_port, memory_3_3_port, memory_3_2_port, 
      memory_3_1_port, memory_3_0_port, memory_4_7_port, memory_4_6_port, 
      memory_4_5_port, memory_4_4_port, memory_4_3_port, memory_4_2_port, 
      memory_4_1_port, memory_4_0_port, memory_5_7_port, memory_5_6_port, 
      memory_5_5_port, memory_5_4_port, memory_5_3_port, memory_5_2_port, 
      memory_5_1_port, memory_5_0_port, memory_6_7_port, memory_6_6_port, 
      memory_6_5_port, memory_6_4_port, memory_6_3_port, memory_6_2_port, 
      memory_6_1_port, memory_6_0_port, memory_7_7_port, memory_7_6_port, 
      memory_7_5_port, memory_7_4_port, memory_7_3_port, memory_7_2_port, 
      memory_7_1_port, memory_7_0_port, memory_8_7_port, memory_8_6_port, 
      memory_8_5_port, memory_8_4_port, memory_8_3_port, memory_8_2_port, 
      memory_8_1_port, memory_8_0_port, memory_9_7_port, memory_9_6_port, 
      memory_9_5_port, memory_9_4_port, memory_9_3_port, memory_9_2_port, 
      memory_9_1_port, memory_9_0_port, memory_10_7_port, memory_10_6_port, 
      memory_10_5_port, memory_10_4_port, memory_10_3_port, memory_10_2_port, 
      memory_10_1_port, memory_10_0_port, memory_11_7_port, memory_11_6_port, 
      memory_11_5_port, memory_11_4_port, memory_11_3_port, memory_11_2_port, 
      memory_11_1_port, memory_11_0_port, memory_12_7_port, memory_12_6_port, 
      memory_12_5_port, memory_12_4_port, memory_12_3_port, memory_12_2_port, 
      memory_12_1_port, memory_12_0_port, memory_13_7_port, memory_13_6_port, 
      memory_13_5_port, memory_13_4_port, memory_13_3_port, memory_13_2_port, 
      memory_13_1_port, memory_13_0_port, memory_14_7_port, memory_14_6_port, 
      memory_14_5_port, memory_14_4_port, memory_14_3_port, memory_14_2_port, 
      memory_14_1_port, memory_14_0_port, memory_15_7_port, memory_15_6_port, 
      memory_15_5_port, memory_15_4_port, memory_15_3_port, memory_15_2_port, 
      memory_15_1_port, memory_15_0_port, memory_16_7_port, memory_16_6_port, 
      memory_16_5_port, memory_16_4_port, memory_16_3_port, memory_16_2_port, 
      memory_16_1_port, memory_16_0_port, memory_17_7_port, memory_17_6_port, 
      memory_17_5_port, memory_17_4_port, memory_17_3_port, memory_17_2_port, 
      memory_17_1_port, memory_17_0_port, memory_18_7_port, memory_18_6_port, 
      memory_18_5_port, memory_18_4_port, memory_18_3_port, memory_18_2_port, 
      memory_18_1_port, memory_18_0_port, memory_19_7_port, memory_19_6_port, 
      memory_19_5_port, memory_19_4_port, memory_19_3_port, memory_19_2_port, 
      memory_19_1_port, memory_19_0_port, memory_20_7_port, memory_20_6_port, 
      memory_20_5_port, memory_20_4_port, memory_20_3_port, memory_20_2_port, 
      memory_20_1_port, memory_20_0_port, memory_21_7_port, memory_21_6_port, 
      memory_21_5_port, memory_21_4_port, memory_21_3_port, memory_21_2_port, 
      memory_21_1_port, memory_21_0_port, memory_22_7_port, memory_22_6_port, 
      memory_22_5_port, memory_22_4_port, memory_22_3_port, memory_22_2_port, 
      memory_22_1_port, memory_22_0_port, memory_23_7_port, memory_23_6_port, 
      memory_23_5_port, memory_23_4_port, memory_23_3_port, memory_23_2_port, 
      memory_23_1_port, memory_23_0_port, memory_24_7_port, memory_24_6_port, 
      memory_24_5_port, memory_24_4_port, memory_24_3_port, memory_24_2_port, 
      memory_24_1_port, memory_24_0_port, memory_25_7_port, memory_25_6_port, 
      memory_25_5_port, memory_25_4_port, memory_25_3_port, memory_25_2_port, 
      memory_25_1_port, memory_25_0_port, memory_26_7_port, memory_26_6_port, 
      memory_26_5_port, memory_26_4_port, memory_26_3_port, memory_26_2_port, 
      memory_26_1_port, memory_26_0_port, memory_27_7_port, memory_27_6_port, 
      memory_27_5_port, memory_27_4_port, memory_27_3_port, memory_27_2_port, 
      memory_27_1_port, memory_27_0_port, memory_28_7_port, memory_28_6_port, 
      memory_28_5_port, memory_28_4_port, memory_28_3_port, memory_28_2_port, 
      memory_28_1_port, memory_28_0_port, memory_29_7_port, memory_29_6_port, 
      memory_29_5_port, memory_29_4_port, memory_29_3_port, memory_29_2_port, 
      memory_29_1_port, memory_29_0_port, memory_30_7_port, memory_30_6_port, 
      memory_30_5_port, memory_30_4_port, memory_30_3_port, memory_30_2_port, 
      memory_30_1_port, memory_30_0_port, memory_31_7_port, memory_31_6_port, 
      memory_31_5_port, memory_31_4_port, memory_31_3_port, memory_31_2_port, 
      memory_31_1_port, memory_31_0_port, N48, N49, N50, N51, N189, N190, N191,
      N192, N193, N195, N333, N334, N335, N336, N337, N338, N339, N340, N341, 
      N342, N343, N344, N345, N346, N347, add_76_aco_carry_1_port, 
      add_76_aco_carry_2_port, add_76_aco_carry_3_port, add_76_aco_carry_4_port
      , sub_72_carry_1_port, sub_72_carry_2_port, sub_72_carry_3_port, 
      sub_72_carry_4_port, add_67_carry_2_port, add_67_carry_3_port, 
      add_67_carry_4_port, r83_carry_2_port, r83_carry_3_port, r83_carry_4_port
      , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32_port, n33_port, n34_port, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43_port, n44_port, n45_port, n46_port, n47, n48_port, n49_port, n50_port
      , n51_port, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189_port, n190_port, n191_port, n192_port, n193_port, n194, n195_port, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333_port, n334_port, n335_port, n336_port,
      n337_port, n338_port, n339_port, n340_port, n341_port, n342_port, 
      n343_port, n344_port, n345_port, n346_port, n347_port, n348, n349, n350, 
      n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
      n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, 
      n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, 
      n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, 
      n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, 
      n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, 
      n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, 
      n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
      n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, 
      n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, 
      n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
      n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
      n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
      n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, 
      n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, 
      n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, 
      n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n855, 
      n857, n859, n861, n863, n864, n865, n866, n867, n909, n910, n911, n912, 
      n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, 
      n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, 
      n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, 
      n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, 
      n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, 
      n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
      n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
      n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
      n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
      n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, 
      n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
      n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, 
      n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
      n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, 
      n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
      n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377 : 
      std_logic;

begin
   DATA <= ( DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, 
      DATA_2_port, DATA_1_port, DATA_0_port );
   OUT_OPCODE <= ( OUT_OPCODE_1_port, OUT_OPCODE_0_port );
   EMPTY <= EMPTY_port;
   FULL <= FULL_port;
   
   X_Logic1_port <= '1';
   state_reg : DFFSR port map( D => X_Logic1_port, CLK => CLK, R => n98, S => 
                           n1372, Q => state);
   FULL_reg : DFFPOSX1 port map( D => n1200, CLK => CLK, Q => FULL_port);
   memory_reg_0_7_inst : DFFPOSX1 port map( D => n1175, CLK => CLK, Q => 
                           memory_0_7_port);
   memory_reg_0_6_inst : DFFPOSX1 port map( D => n1174, CLK => CLK, Q => 
                           memory_0_6_port);
   memory_reg_0_5_inst : DFFPOSX1 port map( D => n1173, CLK => CLK, Q => 
                           memory_0_5_port);
   memory_reg_0_4_inst : DFFPOSX1 port map( D => n1172, CLK => CLK, Q => 
                           memory_0_4_port);
   memory_reg_0_3_inst : DFFPOSX1 port map( D => n1171, CLK => CLK, Q => 
                           memory_0_3_port);
   memory_reg_0_2_inst : DFFPOSX1 port map( D => n1170, CLK => CLK, Q => 
                           memory_0_2_port);
   memory_reg_0_1_inst : DFFPOSX1 port map( D => n1169, CLK => CLK, Q => 
                           memory_0_1_port);
   memory_reg_0_0_inst : DFFPOSX1 port map( D => n1168, CLK => CLK, Q => 
                           memory_0_0_port);
   memory_reg_1_7_inst : DFFPOSX1 port map( D => n1183, CLK => CLK, Q => 
                           memory_1_7_port);
   memory_reg_1_6_inst : DFFPOSX1 port map( D => n1182, CLK => CLK, Q => 
                           memory_1_6_port);
   memory_reg_1_5_inst : DFFPOSX1 port map( D => n1181, CLK => CLK, Q => 
                           memory_1_5_port);
   memory_reg_1_4_inst : DFFPOSX1 port map( D => n1180, CLK => CLK, Q => 
                           memory_1_4_port);
   memory_reg_1_3_inst : DFFPOSX1 port map( D => n1179, CLK => CLK, Q => 
                           memory_1_3_port);
   memory_reg_1_2_inst : DFFPOSX1 port map( D => n1178, CLK => CLK, Q => 
                           memory_1_2_port);
   memory_reg_1_1_inst : DFFPOSX1 port map( D => n1177, CLK => CLK, Q => 
                           memory_1_1_port);
   memory_reg_1_0_inst : DFFPOSX1 port map( D => n1176, CLK => CLK, Q => 
                           memory_1_0_port);
   memory_reg_2_7_inst : DFFPOSX1 port map( D => n1191, CLK => CLK, Q => 
                           memory_2_7_port);
   memory_reg_2_6_inst : DFFPOSX1 port map( D => n1190, CLK => CLK, Q => 
                           memory_2_6_port);
   memory_reg_2_5_inst : DFFPOSX1 port map( D => n1189, CLK => CLK, Q => 
                           memory_2_5_port);
   memory_reg_2_4_inst : DFFPOSX1 port map( D => n1188, CLK => CLK, Q => 
                           memory_2_4_port);
   memory_reg_2_3_inst : DFFPOSX1 port map( D => n1187, CLK => CLK, Q => 
                           memory_2_3_port);
   memory_reg_2_2_inst : DFFPOSX1 port map( D => n1186, CLK => CLK, Q => 
                           memory_2_2_port);
   memory_reg_2_1_inst : DFFPOSX1 port map( D => n1185, CLK => CLK, Q => 
                           memory_2_1_port);
   memory_reg_2_0_inst : DFFPOSX1 port map( D => n1184, CLK => CLK, Q => 
                           memory_2_0_port);
   memory_reg_3_7_inst : DFFPOSX1 port map( D => n1199, CLK => CLK, Q => 
                           memory_3_7_port);
   memory_reg_3_6_inst : DFFPOSX1 port map( D => n1198, CLK => CLK, Q => 
                           memory_3_6_port);
   memory_reg_3_5_inst : DFFPOSX1 port map( D => n1197, CLK => CLK, Q => 
                           memory_3_5_port);
   memory_reg_3_4_inst : DFFPOSX1 port map( D => n1196, CLK => CLK, Q => 
                           memory_3_4_port);
   memory_reg_3_3_inst : DFFPOSX1 port map( D => n1195, CLK => CLK, Q => 
                           memory_3_3_port);
   memory_reg_3_2_inst : DFFPOSX1 port map( D => n1194, CLK => CLK, Q => 
                           memory_3_2_port);
   memory_reg_3_1_inst : DFFPOSX1 port map( D => n1193, CLK => CLK, Q => 
                           memory_3_1_port);
   memory_reg_3_0_inst : DFFPOSX1 port map( D => n1192, CLK => CLK, Q => 
                           memory_3_0_port);
   memory_reg_4_7_inst : DFFPOSX1 port map( D => n1371, CLK => CLK, Q => 
                           memory_4_7_port);
   memory_reg_4_6_inst : DFFPOSX1 port map( D => n1370, CLK => CLK, Q => 
                           memory_4_6_port);
   memory_reg_4_5_inst : DFFPOSX1 port map( D => n1369, CLK => CLK, Q => 
                           memory_4_5_port);
   memory_reg_4_4_inst : DFFPOSX1 port map( D => n1368, CLK => CLK, Q => 
                           memory_4_4_port);
   memory_reg_4_3_inst : DFFPOSX1 port map( D => n1367, CLK => CLK, Q => 
                           memory_4_3_port);
   memory_reg_4_2_inst : DFFPOSX1 port map( D => n1366, CLK => CLK, Q => 
                           memory_4_2_port);
   memory_reg_4_1_inst : DFFPOSX1 port map( D => n1365, CLK => CLK, Q => 
                           memory_4_1_port);
   memory_reg_4_0_inst : DFFPOSX1 port map( D => n1364, CLK => CLK, Q => 
                           memory_4_0_port);
   memory_reg_5_7_inst : DFFPOSX1 port map( D => n1361, CLK => CLK, Q => 
                           memory_5_7_port);
   memory_reg_5_6_inst : DFFPOSX1 port map( D => n1360, CLK => CLK, Q => 
                           memory_5_6_port);
   memory_reg_5_5_inst : DFFPOSX1 port map( D => n1359, CLK => CLK, Q => 
                           memory_5_5_port);
   memory_reg_5_4_inst : DFFPOSX1 port map( D => n1358, CLK => CLK, Q => 
                           memory_5_4_port);
   memory_reg_5_3_inst : DFFPOSX1 port map( D => n1357, CLK => CLK, Q => 
                           memory_5_3_port);
   memory_reg_5_2_inst : DFFPOSX1 port map( D => n1356, CLK => CLK, Q => 
                           memory_5_2_port);
   memory_reg_5_1_inst : DFFPOSX1 port map( D => n1355, CLK => CLK, Q => 
                           memory_5_1_port);
   memory_reg_5_0_inst : DFFPOSX1 port map( D => n1354, CLK => CLK, Q => 
                           memory_5_0_port);
   memory_reg_6_7_inst : DFFPOSX1 port map( D => n1351, CLK => CLK, Q => 
                           memory_6_7_port);
   memory_reg_6_6_inst : DFFPOSX1 port map( D => n1350, CLK => CLK, Q => 
                           memory_6_6_port);
   memory_reg_6_5_inst : DFFPOSX1 port map( D => n1349, CLK => CLK, Q => 
                           memory_6_5_port);
   memory_reg_6_4_inst : DFFPOSX1 port map( D => n1348, CLK => CLK, Q => 
                           memory_6_4_port);
   memory_reg_6_3_inst : DFFPOSX1 port map( D => n1347, CLK => CLK, Q => 
                           memory_6_3_port);
   memory_reg_6_2_inst : DFFPOSX1 port map( D => n1346, CLK => CLK, Q => 
                           memory_6_2_port);
   memory_reg_6_1_inst : DFFPOSX1 port map( D => n1345, CLK => CLK, Q => 
                           memory_6_1_port);
   memory_reg_6_0_inst : DFFPOSX1 port map( D => n1344, CLK => CLK, Q => 
                           memory_6_0_port);
   memory_reg_7_7_inst : DFFPOSX1 port map( D => n1341, CLK => CLK, Q => 
                           memory_7_7_port);
   memory_reg_7_6_inst : DFFPOSX1 port map( D => n1340, CLK => CLK, Q => 
                           memory_7_6_port);
   memory_reg_7_5_inst : DFFPOSX1 port map( D => n1339, CLK => CLK, Q => 
                           memory_7_5_port);
   memory_reg_7_4_inst : DFFPOSX1 port map( D => n1338, CLK => CLK, Q => 
                           memory_7_4_port);
   memory_reg_7_3_inst : DFFPOSX1 port map( D => n1337, CLK => CLK, Q => 
                           memory_7_3_port);
   memory_reg_7_2_inst : DFFPOSX1 port map( D => n1336, CLK => CLK, Q => 
                           memory_7_2_port);
   memory_reg_7_1_inst : DFFPOSX1 port map( D => n1335, CLK => CLK, Q => 
                           memory_7_1_port);
   memory_reg_7_0_inst : DFFPOSX1 port map( D => n1334, CLK => CLK, Q => 
                           memory_7_0_port);
   memory_reg_8_7_inst : DFFPOSX1 port map( D => n1202, CLK => CLK, Q => 
                           memory_8_7_port);
   memory_reg_8_6_inst : DFFPOSX1 port map( D => n1203, CLK => CLK, Q => 
                           memory_8_6_port);
   memory_reg_8_5_inst : DFFPOSX1 port map( D => n1204, CLK => CLK, Q => 
                           memory_8_5_port);
   memory_reg_8_4_inst : DFFPOSX1 port map( D => n1205, CLK => CLK, Q => 
                           memory_8_4_port);
   memory_reg_8_3_inst : DFFPOSX1 port map( D => n1206, CLK => CLK, Q => 
                           memory_8_3_port);
   memory_reg_8_2_inst : DFFPOSX1 port map( D => n1207, CLK => CLK, Q => 
                           memory_8_2_port);
   memory_reg_8_1_inst : DFFPOSX1 port map( D => n1208, CLK => CLK, Q => 
                           memory_8_1_port);
   memory_reg_8_0_inst : DFFPOSX1 port map( D => n1209, CLK => CLK, Q => 
                           memory_8_0_port);
   memory_reg_9_7_inst : DFFPOSX1 port map( D => n1210, CLK => CLK, Q => 
                           memory_9_7_port);
   memory_reg_9_6_inst : DFFPOSX1 port map( D => n1211, CLK => CLK, Q => 
                           memory_9_6_port);
   memory_reg_9_5_inst : DFFPOSX1 port map( D => n1212, CLK => CLK, Q => 
                           memory_9_5_port);
   memory_reg_9_4_inst : DFFPOSX1 port map( D => n1213, CLK => CLK, Q => 
                           memory_9_4_port);
   memory_reg_9_3_inst : DFFPOSX1 port map( D => n1214, CLK => CLK, Q => 
                           memory_9_3_port);
   memory_reg_9_2_inst : DFFPOSX1 port map( D => n1215, CLK => CLK, Q => 
                           memory_9_2_port);
   memory_reg_9_1_inst : DFFPOSX1 port map( D => n1216, CLK => CLK, Q => 
                           memory_9_1_port);
   memory_reg_9_0_inst : DFFPOSX1 port map( D => n1217, CLK => CLK, Q => 
                           memory_9_0_port);
   memory_reg_10_7_inst : DFFPOSX1 port map( D => n1218, CLK => CLK, Q => 
                           memory_10_7_port);
   memory_reg_10_6_inst : DFFPOSX1 port map( D => n1219, CLK => CLK, Q => 
                           memory_10_6_port);
   memory_reg_10_5_inst : DFFPOSX1 port map( D => n1220, CLK => CLK, Q => 
                           memory_10_5_port);
   memory_reg_10_4_inst : DFFPOSX1 port map( D => n1221, CLK => CLK, Q => 
                           memory_10_4_port);
   memory_reg_10_3_inst : DFFPOSX1 port map( D => n1222, CLK => CLK, Q => 
                           memory_10_3_port);
   memory_reg_10_2_inst : DFFPOSX1 port map( D => n1223, CLK => CLK, Q => 
                           memory_10_2_port);
   memory_reg_10_1_inst : DFFPOSX1 port map( D => n1224, CLK => CLK, Q => 
                           memory_10_1_port);
   memory_reg_10_0_inst : DFFPOSX1 port map( D => n1225, CLK => CLK, Q => 
                           memory_10_0_port);
   memory_reg_11_7_inst : DFFPOSX1 port map( D => n1226, CLK => CLK, Q => 
                           memory_11_7_port);
   memory_reg_11_6_inst : DFFPOSX1 port map( D => n1227, CLK => CLK, Q => 
                           memory_11_6_port);
   memory_reg_11_5_inst : DFFPOSX1 port map( D => n1228, CLK => CLK, Q => 
                           memory_11_5_port);
   memory_reg_11_4_inst : DFFPOSX1 port map( D => n1229, CLK => CLK, Q => 
                           memory_11_4_port);
   memory_reg_11_3_inst : DFFPOSX1 port map( D => n1230, CLK => CLK, Q => 
                           memory_11_3_port);
   memory_reg_11_2_inst : DFFPOSX1 port map( D => n1231, CLK => CLK, Q => 
                           memory_11_2_port);
   memory_reg_11_1_inst : DFFPOSX1 port map( D => n1232, CLK => CLK, Q => 
                           memory_11_1_port);
   memory_reg_11_0_inst : DFFPOSX1 port map( D => n1233, CLK => CLK, Q => 
                           memory_11_0_port);
   memory_reg_12_7_inst : DFFPOSX1 port map( D => n1064, CLK => CLK, Q => 
                           memory_12_7_port);
   memory_reg_12_6_inst : DFFPOSX1 port map( D => n1065, CLK => CLK, Q => 
                           memory_12_6_port);
   memory_reg_12_5_inst : DFFPOSX1 port map( D => n1066, CLK => CLK, Q => 
                           memory_12_5_port);
   memory_reg_12_4_inst : DFFPOSX1 port map( D => n1067, CLK => CLK, Q => 
                           memory_12_4_port);
   memory_reg_12_3_inst : DFFPOSX1 port map( D => n1068, CLK => CLK, Q => 
                           memory_12_3_port);
   memory_reg_12_2_inst : DFFPOSX1 port map( D => n1069, CLK => CLK, Q => 
                           memory_12_2_port);
   memory_reg_12_1_inst : DFFPOSX1 port map( D => n1070, CLK => CLK, Q => 
                           memory_12_1_port);
   memory_reg_12_0_inst : DFFPOSX1 port map( D => n1071, CLK => CLK, Q => 
                           memory_12_0_port);
   memory_reg_13_7_inst : DFFPOSX1 port map( D => n1022, CLK => CLK, Q => 
                           memory_13_7_port);
   memory_reg_13_6_inst : DFFPOSX1 port map( D => n1023, CLK => CLK, Q => 
                           memory_13_6_port);
   memory_reg_13_5_inst : DFFPOSX1 port map( D => n1024, CLK => CLK, Q => 
                           memory_13_5_port);
   memory_reg_13_4_inst : DFFPOSX1 port map( D => n1025, CLK => CLK, Q => 
                           memory_13_4_port);
   memory_reg_13_3_inst : DFFPOSX1 port map( D => n1026, CLK => CLK, Q => 
                           memory_13_3_port);
   memory_reg_13_2_inst : DFFPOSX1 port map( D => n1027, CLK => CLK, Q => 
                           memory_13_2_port);
   memory_reg_13_1_inst : DFFPOSX1 port map( D => n1028, CLK => CLK, Q => 
                           memory_13_1_port);
   memory_reg_13_0_inst : DFFPOSX1 port map( D => n1029, CLK => CLK, Q => 
                           memory_13_0_port);
   memory_reg_14_7_inst : DFFPOSX1 port map( D => n1014, CLK => CLK, Q => 
                           memory_14_7_port);
   memory_reg_14_6_inst : DFFPOSX1 port map( D => n1015, CLK => CLK, Q => 
                           memory_14_6_port);
   memory_reg_14_5_inst : DFFPOSX1 port map( D => n1016, CLK => CLK, Q => 
                           memory_14_5_port);
   memory_reg_14_4_inst : DFFPOSX1 port map( D => n1017, CLK => CLK, Q => 
                           memory_14_4_port);
   memory_reg_14_3_inst : DFFPOSX1 port map( D => n1018, CLK => CLK, Q => 
                           memory_14_3_port);
   memory_reg_14_2_inst : DFFPOSX1 port map( D => n1019, CLK => CLK, Q => 
                           memory_14_2_port);
   memory_reg_14_1_inst : DFFPOSX1 port map( D => n1020, CLK => CLK, Q => 
                           memory_14_1_port);
   memory_reg_14_0_inst : DFFPOSX1 port map( D => n1021, CLK => CLK, Q => 
                           memory_14_0_port);
   memory_reg_15_7_inst : DFFPOSX1 port map( D => n1006, CLK => CLK, Q => 
                           memory_15_7_port);
   memory_reg_15_6_inst : DFFPOSX1 port map( D => n1007, CLK => CLK, Q => 
                           memory_15_6_port);
   memory_reg_15_5_inst : DFFPOSX1 port map( D => n1008, CLK => CLK, Q => 
                           memory_15_5_port);
   memory_reg_15_4_inst : DFFPOSX1 port map( D => n1009, CLK => CLK, Q => 
                           memory_15_4_port);
   memory_reg_15_3_inst : DFFPOSX1 port map( D => n1010, CLK => CLK, Q => 
                           memory_15_3_port);
   memory_reg_15_2_inst : DFFPOSX1 port map( D => n1011, CLK => CLK, Q => 
                           memory_15_2_port);
   memory_reg_15_1_inst : DFFPOSX1 port map( D => n1012, CLK => CLK, Q => 
                           memory_15_1_port);
   memory_reg_15_0_inst : DFFPOSX1 port map( D => n1013, CLK => CLK, Q => 
                           memory_15_0_port);
   memory_reg_16_7_inst : DFFPOSX1 port map( D => n1234, CLK => CLK, Q => 
                           memory_16_7_port);
   memory_reg_16_6_inst : DFFPOSX1 port map( D => n1235, CLK => CLK, Q => 
                           memory_16_6_port);
   memory_reg_16_5_inst : DFFPOSX1 port map( D => n1236, CLK => CLK, Q => 
                           memory_16_5_port);
   memory_reg_16_4_inst : DFFPOSX1 port map( D => n1237, CLK => CLK, Q => 
                           memory_16_4_port);
   memory_reg_16_3_inst : DFFPOSX1 port map( D => n1238, CLK => CLK, Q => 
                           memory_16_3_port);
   memory_reg_16_2_inst : DFFPOSX1 port map( D => n1239, CLK => CLK, Q => 
                           memory_16_2_port);
   memory_reg_16_1_inst : DFFPOSX1 port map( D => n1240, CLK => CLK, Q => 
                           memory_16_1_port);
   memory_reg_16_0_inst : DFFPOSX1 port map( D => n1241, CLK => CLK, Q => 
                           memory_16_0_port);
   memory_reg_17_7_inst : DFFPOSX1 port map( D => n1242, CLK => CLK, Q => 
                           memory_17_7_port);
   memory_reg_17_6_inst : DFFPOSX1 port map( D => n1243, CLK => CLK, Q => 
                           memory_17_6_port);
   memory_reg_17_5_inst : DFFPOSX1 port map( D => n1244, CLK => CLK, Q => 
                           memory_17_5_port);
   memory_reg_17_4_inst : DFFPOSX1 port map( D => n1245, CLK => CLK, Q => 
                           memory_17_4_port);
   memory_reg_17_3_inst : DFFPOSX1 port map( D => n1246, CLK => CLK, Q => 
                           memory_17_3_port);
   memory_reg_17_2_inst : DFFPOSX1 port map( D => n1247, CLK => CLK, Q => 
                           memory_17_2_port);
   memory_reg_17_1_inst : DFFPOSX1 port map( D => n1248, CLK => CLK, Q => 
                           memory_17_1_port);
   memory_reg_17_0_inst : DFFPOSX1 port map( D => n1249, CLK => CLK, Q => 
                           memory_17_0_port);
   memory_reg_18_7_inst : DFFPOSX1 port map( D => n1250, CLK => CLK, Q => 
                           memory_18_7_port);
   memory_reg_18_6_inst : DFFPOSX1 port map( D => n1251, CLK => CLK, Q => 
                           memory_18_6_port);
   memory_reg_18_5_inst : DFFPOSX1 port map( D => n1252, CLK => CLK, Q => 
                           memory_18_5_port);
   memory_reg_18_4_inst : DFFPOSX1 port map( D => n1253, CLK => CLK, Q => 
                           memory_18_4_port);
   memory_reg_18_3_inst : DFFPOSX1 port map( D => n1254, CLK => CLK, Q => 
                           memory_18_3_port);
   memory_reg_18_2_inst : DFFPOSX1 port map( D => n1255, CLK => CLK, Q => 
                           memory_18_2_port);
   memory_reg_18_1_inst : DFFPOSX1 port map( D => n1256, CLK => CLK, Q => 
                           memory_18_1_port);
   memory_reg_18_0_inst : DFFPOSX1 port map( D => n1257, CLK => CLK, Q => 
                           memory_18_0_port);
   memory_reg_19_7_inst : DFFPOSX1 port map( D => n1258, CLK => CLK, Q => 
                           memory_19_7_port);
   memory_reg_19_6_inst : DFFPOSX1 port map( D => n1259, CLK => CLK, Q => 
                           memory_19_6_port);
   memory_reg_19_5_inst : DFFPOSX1 port map( D => n1260, CLK => CLK, Q => 
                           memory_19_5_port);
   memory_reg_19_4_inst : DFFPOSX1 port map( D => n1261, CLK => CLK, Q => 
                           memory_19_4_port);
   memory_reg_19_3_inst : DFFPOSX1 port map( D => n1262, CLK => CLK, Q => 
                           memory_19_3_port);
   memory_reg_19_2_inst : DFFPOSX1 port map( D => n1263, CLK => CLK, Q => 
                           memory_19_2_port);
   memory_reg_19_1_inst : DFFPOSX1 port map( D => n1264, CLK => CLK, Q => 
                           memory_19_1_port);
   memory_reg_19_0_inst : DFFPOSX1 port map( D => n1265, CLK => CLK, Q => 
                           memory_19_0_port);
   memory_reg_20_7_inst : DFFPOSX1 port map( D => n998, CLK => CLK, Q => 
                           memory_20_7_port);
   memory_reg_20_6_inst : DFFPOSX1 port map( D => n999, CLK => CLK, Q => 
                           memory_20_6_port);
   memory_reg_20_5_inst : DFFPOSX1 port map( D => n1000, CLK => CLK, Q => 
                           memory_20_5_port);
   memory_reg_20_4_inst : DFFPOSX1 port map( D => n1001, CLK => CLK, Q => 
                           memory_20_4_port);
   memory_reg_20_3_inst : DFFPOSX1 port map( D => n1002, CLK => CLK, Q => 
                           memory_20_3_port);
   memory_reg_20_2_inst : DFFPOSX1 port map( D => n1003, CLK => CLK, Q => 
                           memory_20_2_port);
   memory_reg_20_1_inst : DFFPOSX1 port map( D => n1004, CLK => CLK, Q => 
                           memory_20_1_port);
   memory_reg_20_0_inst : DFFPOSX1 port map( D => n1005, CLK => CLK, Q => 
                           memory_20_0_port);
   memory_reg_21_7_inst : DFFPOSX1 port map( D => n990, CLK => CLK, Q => 
                           memory_21_7_port);
   memory_reg_21_6_inst : DFFPOSX1 port map( D => n991, CLK => CLK, Q => 
                           memory_21_6_port);
   memory_reg_21_5_inst : DFFPOSX1 port map( D => n992, CLK => CLK, Q => 
                           memory_21_5_port);
   memory_reg_21_4_inst : DFFPOSX1 port map( D => n993, CLK => CLK, Q => 
                           memory_21_4_port);
   memory_reg_21_3_inst : DFFPOSX1 port map( D => n994, CLK => CLK, Q => 
                           memory_21_3_port);
   memory_reg_21_2_inst : DFFPOSX1 port map( D => n995, CLK => CLK, Q => 
                           memory_21_2_port);
   memory_reg_21_1_inst : DFFPOSX1 port map( D => n996, CLK => CLK, Q => 
                           memory_21_1_port);
   memory_reg_21_0_inst : DFFPOSX1 port map( D => n997, CLK => CLK, Q => 
                           memory_21_0_port);
   memory_reg_22_7_inst : DFFPOSX1 port map( D => n982, CLK => CLK, Q => 
                           memory_22_7_port);
   memory_reg_22_6_inst : DFFPOSX1 port map( D => n983, CLK => CLK, Q => 
                           memory_22_6_port);
   memory_reg_22_5_inst : DFFPOSX1 port map( D => n984, CLK => CLK, Q => 
                           memory_22_5_port);
   memory_reg_22_4_inst : DFFPOSX1 port map( D => n985, CLK => CLK, Q => 
                           memory_22_4_port);
   memory_reg_22_3_inst : DFFPOSX1 port map( D => n986, CLK => CLK, Q => 
                           memory_22_3_port);
   memory_reg_22_2_inst : DFFPOSX1 port map( D => n987, CLK => CLK, Q => 
                           memory_22_2_port);
   memory_reg_22_1_inst : DFFPOSX1 port map( D => n988, CLK => CLK, Q => 
                           memory_22_1_port);
   memory_reg_22_0_inst : DFFPOSX1 port map( D => n989, CLK => CLK, Q => 
                           memory_22_0_port);
   memory_reg_23_7_inst : DFFPOSX1 port map( D => n974, CLK => CLK, Q => 
                           memory_23_7_port);
   memory_reg_23_6_inst : DFFPOSX1 port map( D => n975, CLK => CLK, Q => 
                           memory_23_6_port);
   memory_reg_23_5_inst : DFFPOSX1 port map( D => n976, CLK => CLK, Q => 
                           memory_23_5_port);
   memory_reg_23_4_inst : DFFPOSX1 port map( D => n977, CLK => CLK, Q => 
                           memory_23_4_port);
   memory_reg_23_3_inst : DFFPOSX1 port map( D => n978, CLK => CLK, Q => 
                           memory_23_3_port);
   memory_reg_23_2_inst : DFFPOSX1 port map( D => n979, CLK => CLK, Q => 
                           memory_23_2_port);
   memory_reg_23_1_inst : DFFPOSX1 port map( D => n980, CLK => CLK, Q => 
                           memory_23_1_port);
   memory_reg_23_0_inst : DFFPOSX1 port map( D => n981, CLK => CLK, Q => 
                           memory_23_0_port);
   memory_reg_24_7_inst : DFFPOSX1 port map( D => n966, CLK => CLK, Q => 
                           memory_24_7_port);
   memory_reg_24_6_inst : DFFPOSX1 port map( D => n967, CLK => CLK, Q => 
                           memory_24_6_port);
   memory_reg_24_5_inst : DFFPOSX1 port map( D => n968, CLK => CLK, Q => 
                           memory_24_5_port);
   memory_reg_24_4_inst : DFFPOSX1 port map( D => n969, CLK => CLK, Q => 
                           memory_24_4_port);
   memory_reg_24_3_inst : DFFPOSX1 port map( D => n970, CLK => CLK, Q => 
                           memory_24_3_port);
   memory_reg_24_2_inst : DFFPOSX1 port map( D => n971, CLK => CLK, Q => 
                           memory_24_2_port);
   memory_reg_24_1_inst : DFFPOSX1 port map( D => n972, CLK => CLK, Q => 
                           memory_24_1_port);
   memory_reg_24_0_inst : DFFPOSX1 port map( D => n973, CLK => CLK, Q => 
                           memory_24_0_port);
   memory_reg_25_7_inst : DFFPOSX1 port map( D => n958, CLK => CLK, Q => 
                           memory_25_7_port);
   memory_reg_25_6_inst : DFFPOSX1 port map( D => n959, CLK => CLK, Q => 
                           memory_25_6_port);
   memory_reg_25_5_inst : DFFPOSX1 port map( D => n960, CLK => CLK, Q => 
                           memory_25_5_port);
   memory_reg_25_4_inst : DFFPOSX1 port map( D => n961, CLK => CLK, Q => 
                           memory_25_4_port);
   memory_reg_25_3_inst : DFFPOSX1 port map( D => n962, CLK => CLK, Q => 
                           memory_25_3_port);
   memory_reg_25_2_inst : DFFPOSX1 port map( D => n963, CLK => CLK, Q => 
                           memory_25_2_port);
   memory_reg_25_1_inst : DFFPOSX1 port map( D => n964, CLK => CLK, Q => 
                           memory_25_1_port);
   memory_reg_25_0_inst : DFFPOSX1 port map( D => n965, CLK => CLK, Q => 
                           memory_25_0_port);
   memory_reg_26_7_inst : DFFPOSX1 port map( D => n950, CLK => CLK, Q => 
                           memory_26_7_port);
   memory_reg_26_6_inst : DFFPOSX1 port map( D => n951, CLK => CLK, Q => 
                           memory_26_6_port);
   memory_reg_26_5_inst : DFFPOSX1 port map( D => n952, CLK => CLK, Q => 
                           memory_26_5_port);
   memory_reg_26_4_inst : DFFPOSX1 port map( D => n953, CLK => CLK, Q => 
                           memory_26_4_port);
   memory_reg_26_3_inst : DFFPOSX1 port map( D => n954, CLK => CLK, Q => 
                           memory_26_3_port);
   memory_reg_26_2_inst : DFFPOSX1 port map( D => n955, CLK => CLK, Q => 
                           memory_26_2_port);
   memory_reg_26_1_inst : DFFPOSX1 port map( D => n956, CLK => CLK, Q => 
                           memory_26_1_port);
   memory_reg_26_0_inst : DFFPOSX1 port map( D => n957, CLK => CLK, Q => 
                           memory_26_0_port);
   memory_reg_27_7_inst : DFFPOSX1 port map( D => n942, CLK => CLK, Q => 
                           memory_27_7_port);
   memory_reg_27_6_inst : DFFPOSX1 port map( D => n943, CLK => CLK, Q => 
                           memory_27_6_port);
   memory_reg_27_5_inst : DFFPOSX1 port map( D => n944, CLK => CLK, Q => 
                           memory_27_5_port);
   memory_reg_27_4_inst : DFFPOSX1 port map( D => n945, CLK => CLK, Q => 
                           memory_27_4_port);
   memory_reg_27_3_inst : DFFPOSX1 port map( D => n946, CLK => CLK, Q => 
                           memory_27_3_port);
   memory_reg_27_2_inst : DFFPOSX1 port map( D => n947, CLK => CLK, Q => 
                           memory_27_2_port);
   memory_reg_27_1_inst : DFFPOSX1 port map( D => n948, CLK => CLK, Q => 
                           memory_27_1_port);
   memory_reg_27_0_inst : DFFPOSX1 port map( D => n949, CLK => CLK, Q => 
                           memory_27_0_port);
   memory_reg_28_7_inst : DFFPOSX1 port map( D => n1266, CLK => CLK, Q => 
                           memory_28_7_port);
   memory_reg_28_6_inst : DFFPOSX1 port map( D => n1267, CLK => CLK, Q => 
                           memory_28_6_port);
   memory_reg_28_5_inst : DFFPOSX1 port map( D => n1268, CLK => CLK, Q => 
                           memory_28_5_port);
   memory_reg_28_4_inst : DFFPOSX1 port map( D => n1269, CLK => CLK, Q => 
                           memory_28_4_port);
   memory_reg_28_3_inst : DFFPOSX1 port map( D => n1270, CLK => CLK, Q => 
                           memory_28_3_port);
   memory_reg_28_2_inst : DFFPOSX1 port map( D => n1271, CLK => CLK, Q => 
                           memory_28_2_port);
   memory_reg_28_1_inst : DFFPOSX1 port map( D => n1272, CLK => CLK, Q => 
                           memory_28_1_port);
   memory_reg_28_0_inst : DFFPOSX1 port map( D => n1273, CLK => CLK, Q => 
                           memory_28_0_port);
   memory_reg_29_7_inst : DFFPOSX1 port map( D => n1274, CLK => CLK, Q => 
                           memory_29_7_port);
   memory_reg_29_6_inst : DFFPOSX1 port map( D => n1275, CLK => CLK, Q => 
                           memory_29_6_port);
   memory_reg_29_5_inst : DFFPOSX1 port map( D => n1276, CLK => CLK, Q => 
                           memory_29_5_port);
   memory_reg_29_4_inst : DFFPOSX1 port map( D => n1277, CLK => CLK, Q => 
                           memory_29_4_port);
   memory_reg_29_3_inst : DFFPOSX1 port map( D => n1278, CLK => CLK, Q => 
                           memory_29_3_port);
   memory_reg_29_2_inst : DFFPOSX1 port map( D => n1279, CLK => CLK, Q => 
                           memory_29_2_port);
   memory_reg_29_1_inst : DFFPOSX1 port map( D => n1280, CLK => CLK, Q => 
                           memory_29_1_port);
   memory_reg_29_0_inst : DFFPOSX1 port map( D => n1281, CLK => CLK, Q => 
                           memory_29_0_port);
   memory_reg_30_7_inst : DFFPOSX1 port map( D => n1282, CLK => CLK, Q => 
                           memory_30_7_port);
   memory_reg_30_6_inst : DFFPOSX1 port map( D => n1283, CLK => CLK, Q => 
                           memory_30_6_port);
   memory_reg_30_5_inst : DFFPOSX1 port map( D => n1284, CLK => CLK, Q => 
                           memory_30_5_port);
   memory_reg_30_4_inst : DFFPOSX1 port map( D => n1285, CLK => CLK, Q => 
                           memory_30_4_port);
   memory_reg_30_3_inst : DFFPOSX1 port map( D => n1286, CLK => CLK, Q => 
                           memory_30_3_port);
   memory_reg_30_2_inst : DFFPOSX1 port map( D => n1287, CLK => CLK, Q => 
                           memory_30_2_port);
   memory_reg_30_1_inst : DFFPOSX1 port map( D => n1288, CLK => CLK, Q => 
                           memory_30_1_port);
   memory_reg_30_0_inst : DFFPOSX1 port map( D => n1289, CLK => CLK, Q => 
                           memory_30_0_port);
   memory_reg_31_7_inst : DFFPOSX1 port map( D => n1290, CLK => CLK, Q => 
                           memory_31_7_port);
   memory_reg_31_6_inst : DFFPOSX1 port map( D => n1291, CLK => CLK, Q => 
                           memory_31_6_port);
   memory_reg_31_5_inst : DFFPOSX1 port map( D => n1292, CLK => CLK, Q => 
                           memory_31_5_port);
   memory_reg_31_4_inst : DFFPOSX1 port map( D => n1293, CLK => CLK, Q => 
                           memory_31_4_port);
   memory_reg_31_3_inst : DFFPOSX1 port map( D => n1294, CLK => CLK, Q => 
                           memory_31_3_port);
   memory_reg_31_2_inst : DFFPOSX1 port map( D => n1295, CLK => CLK, Q => 
                           memory_31_2_port);
   memory_reg_31_1_inst : DFFPOSX1 port map( D => n1296, CLK => CLK, Q => 
                           memory_31_1_port);
   memory_reg_31_0_inst : DFFPOSX1 port map( D => n1297, CLK => CLK, Q => 
                           memory_31_0_port);
   opcode_reg_0_1_inst : DFFPOSX1 port map( D => n935, CLK => CLK, Q => 
                           opcode_0_1_port);
   opcode_reg_0_0_inst : DFFPOSX1 port map( D => n934, CLK => CLK, Q => 
                           opcode_0_0_port);
   opcode_reg_1_1_inst : DFFPOSX1 port map( D => n937, CLK => CLK, Q => 
                           opcode_1_1_port);
   opcode_reg_1_0_inst : DFFPOSX1 port map( D => n936, CLK => CLK, Q => 
                           opcode_1_0_port);
   opcode_reg_2_1_inst : DFFPOSX1 port map( D => n939, CLK => CLK, Q => 
                           opcode_2_1_port);
   opcode_reg_2_0_inst : DFFPOSX1 port map( D => n938, CLK => CLK, Q => 
                           opcode_2_0_port);
   opcode_reg_3_1_inst : DFFPOSX1 port map( D => n941, CLK => CLK, Q => 
                           opcode_3_1_port);
   opcode_reg_3_0_inst : DFFPOSX1 port map( D => n940, CLK => CLK, Q => 
                           opcode_3_0_port);
   opcode_reg_4_1_inst : DFFPOSX1 port map( D => n1363, CLK => CLK, Q => 
                           opcode_4_1_port);
   opcode_reg_4_0_inst : DFFPOSX1 port map( D => n1362, CLK => CLK, Q => 
                           opcode_4_0_port);
   opcode_reg_5_1_inst : DFFPOSX1 port map( D => n1353, CLK => CLK, Q => 
                           opcode_5_1_port);
   opcode_reg_5_0_inst : DFFPOSX1 port map( D => n1352, CLK => CLK, Q => 
                           opcode_5_0_port);
   opcode_reg_6_1_inst : DFFPOSX1 port map( D => n1343, CLK => CLK, Q => 
                           opcode_6_1_port);
   opcode_reg_6_0_inst : DFFPOSX1 port map( D => n1342, CLK => CLK, Q => 
                           opcode_6_0_port);
   opcode_reg_7_1_inst : DFFPOSX1 port map( D => n1333, CLK => CLK, Q => 
                           opcode_7_1_port);
   opcode_reg_7_0_inst : DFFPOSX1 port map( D => n1332, CLK => CLK, Q => 
                           opcode_7_0_port);
   opcode_reg_8_1_inst : DFFPOSX1 port map( D => n1298, CLK => CLK, Q => 
                           opcode_8_1_port);
   opcode_reg_8_0_inst : DFFPOSX1 port map( D => n1299, CLK => CLK, Q => 
                           opcode_8_0_port);
   opcode_reg_9_1_inst : DFFPOSX1 port map( D => n1300, CLK => CLK, Q => 
                           opcode_9_1_port);
   opcode_reg_9_0_inst : DFFPOSX1 port map( D => n1301, CLK => CLK, Q => 
                           opcode_9_0_port);
   opcode_reg_10_1_inst : DFFPOSX1 port map( D => n1302, CLK => CLK, Q => 
                           opcode_10_1_port);
   opcode_reg_10_0_inst : DFFPOSX1 port map( D => n1303, CLK => CLK, Q => 
                           opcode_10_0_port);
   opcode_reg_11_1_inst : DFFPOSX1 port map( D => n1304, CLK => CLK, Q => 
                           opcode_11_1_port);
   opcode_reg_11_0_inst : DFFPOSX1 port map( D => n1305, CLK => CLK, Q => 
                           opcode_11_0_port);
   opcode_reg_12_1_inst : DFFPOSX1 port map( D => n932, CLK => CLK, Q => 
                           opcode_12_1_port);
   opcode_reg_12_0_inst : DFFPOSX1 port map( D => n933, CLK => CLK, Q => 
                           opcode_12_0_port);
   opcode_reg_13_1_inst : DFFPOSX1 port map( D => n930, CLK => CLK, Q => 
                           opcode_13_1_port);
   opcode_reg_13_0_inst : DFFPOSX1 port map( D => n931, CLK => CLK, Q => 
                           opcode_13_0_port);
   opcode_reg_14_1_inst : DFFPOSX1 port map( D => n928, CLK => CLK, Q => 
                           opcode_14_1_port);
   opcode_reg_14_0_inst : DFFPOSX1 port map( D => n929, CLK => CLK, Q => 
                           opcode_14_0_port);
   opcode_reg_15_1_inst : DFFPOSX1 port map( D => n926, CLK => CLK, Q => 
                           opcode_15_1_port);
   opcode_reg_15_0_inst : DFFPOSX1 port map( D => n927, CLK => CLK, Q => 
                           opcode_15_0_port);
   opcode_reg_16_1_inst : DFFPOSX1 port map( D => n1306, CLK => CLK, Q => 
                           opcode_16_1_port);
   opcode_reg_16_0_inst : DFFPOSX1 port map( D => n1307, CLK => CLK, Q => 
                           opcode_16_0_port);
   opcode_reg_17_1_inst : DFFPOSX1 port map( D => n1308, CLK => CLK, Q => 
                           opcode_17_1_port);
   opcode_reg_17_0_inst : DFFPOSX1 port map( D => n1309, CLK => CLK, Q => 
                           opcode_17_0_port);
   opcode_reg_18_1_inst : DFFPOSX1 port map( D => n1310, CLK => CLK, Q => 
                           opcode_18_1_port);
   opcode_reg_18_0_inst : DFFPOSX1 port map( D => n1311, CLK => CLK, Q => 
                           opcode_18_0_port);
   opcode_reg_19_1_inst : DFFPOSX1 port map( D => n1312, CLK => CLK, Q => 
                           opcode_19_1_port);
   opcode_reg_19_0_inst : DFFPOSX1 port map( D => n1313, CLK => CLK, Q => 
                           opcode_19_0_port);
   opcode_reg_20_1_inst : DFFPOSX1 port map( D => n924, CLK => CLK, Q => 
                           opcode_20_1_port);
   opcode_reg_20_0_inst : DFFPOSX1 port map( D => n925, CLK => CLK, Q => 
                           opcode_20_0_port);
   opcode_reg_21_1_inst : DFFPOSX1 port map( D => n922, CLK => CLK, Q => 
                           opcode_21_1_port);
   opcode_reg_21_0_inst : DFFPOSX1 port map( D => n923, CLK => CLK, Q => 
                           opcode_21_0_port);
   opcode_reg_22_1_inst : DFFPOSX1 port map( D => n920, CLK => CLK, Q => 
                           opcode_22_1_port);
   opcode_reg_22_0_inst : DFFPOSX1 port map( D => n921, CLK => CLK, Q => 
                           opcode_22_0_port);
   opcode_reg_23_1_inst : DFFPOSX1 port map( D => n918, CLK => CLK, Q => 
                           opcode_23_1_port);
   opcode_reg_23_0_inst : DFFPOSX1 port map( D => n919, CLK => CLK, Q => 
                           opcode_23_0_port);
   opcode_reg_24_1_inst : DFFPOSX1 port map( D => n916, CLK => CLK, Q => 
                           opcode_24_1_port);
   opcode_reg_24_0_inst : DFFPOSX1 port map( D => n917, CLK => CLK, Q => 
                           opcode_24_0_port);
   opcode_reg_25_1_inst : DFFPOSX1 port map( D => n914, CLK => CLK, Q => 
                           opcode_25_1_port);
   opcode_reg_25_0_inst : DFFPOSX1 port map( D => n915, CLK => CLK, Q => 
                           opcode_25_0_port);
   opcode_reg_26_1_inst : DFFPOSX1 port map( D => n912, CLK => CLK, Q => 
                           opcode_26_1_port);
   opcode_reg_26_0_inst : DFFPOSX1 port map( D => n913, CLK => CLK, Q => 
                           opcode_26_0_port);
   opcode_reg_27_1_inst : DFFPOSX1 port map( D => n910, CLK => CLK, Q => 
                           opcode_27_1_port);
   opcode_reg_27_0_inst : DFFPOSX1 port map( D => n911, CLK => CLK, Q => 
                           opcode_27_0_port);
   opcode_reg_28_1_inst : DFFPOSX1 port map( D => n1314, CLK => CLK, Q => 
                           opcode_28_1_port);
   opcode_reg_28_0_inst : DFFPOSX1 port map( D => n1315, CLK => CLK, Q => 
                           opcode_28_0_port);
   opcode_reg_29_1_inst : DFFPOSX1 port map( D => n1316, CLK => CLK, Q => 
                           opcode_29_1_port);
   opcode_reg_29_0_inst : DFFPOSX1 port map( D => n1317, CLK => CLK, Q => 
                           opcode_29_0_port);
   opcode_reg_30_1_inst : DFFPOSX1 port map( D => n1318, CLK => CLK, Q => 
                           opcode_30_1_port);
   opcode_reg_30_0_inst : DFFPOSX1 port map( D => n1319, CLK => CLK, Q => 
                           opcode_30_0_port);
   opcode_reg_31_1_inst : DFFPOSX1 port map( D => n1320, CLK => CLK, Q => 
                           opcode_31_1_port);
   opcode_reg_31_0_inst : DFFPOSX1 port map( D => n1321, CLK => CLK, Q => 
                           opcode_31_0_port);
   DATA_reg_7_inst : DFFPOSX1 port map( D => n1322, CLK => CLK, Q => 
                           DATA_7_port);
   DATA_reg_6_inst : DFFPOSX1 port map( D => n1323, CLK => CLK, Q => 
                           DATA_6_port);
   DATA_reg_5_inst : DFFPOSX1 port map( D => n1324, CLK => CLK, Q => 
                           DATA_5_port);
   DATA_reg_4_inst : DFFPOSX1 port map( D => n1325, CLK => CLK, Q => 
                           DATA_4_port);
   DATA_reg_3_inst : DFFPOSX1 port map( D => n1326, CLK => CLK, Q => 
                           DATA_3_port);
   DATA_reg_2_inst : DFFPOSX1 port map( D => n1327, CLK => CLK, Q => 
                           DATA_2_port);
   DATA_reg_1_inst : DFFPOSX1 port map( D => n1328, CLK => CLK, Q => 
                           DATA_1_port);
   DATA_reg_0_inst : DFFPOSX1 port map( D => n1329, CLK => CLK, Q => 
                           DATA_0_port);
   OUT_OPCODE_reg_1_inst : DFFPOSX1 port map( D => n1330, CLK => CLK, Q => 
                           OUT_OPCODE_1_port);
   OUT_OPCODE_reg_0_inst : DFFPOSX1 port map( D => n1331, CLK => CLK, Q => 
                           OUT_OPCODE_0_port);
   EMPTY_reg : DFFPOSX1 port map( D => n1201, CLK => CLK, Q => EMPTY_port);
   n1372 <= '1';
   sub_72_U2_1 : FAX1 port map( A => n78, B => n517, C => sub_72_carry_1_port, 
                           YC => sub_72_carry_2_port, YS => N190);
   sub_72_U2_2 : FAX1 port map( A => n76, B => n855, C => sub_72_carry_2_port, 
                           YC => sub_72_carry_3_port, YS => N191);
   sub_72_U2_3 : FAX1 port map( A => n83, B => n824, C => sub_72_carry_3_port, 
                           YC => sub_72_carry_4_port, YS => N192);
   sub_72_U2_4 : FAX1 port map( A => writeptr_4_port, B => n845, C => 
                           sub_72_carry_4_port, YC => n103, YS => N193);
   add_67_U1_1_1 : HAX1 port map( A => n79, B => n81, YC => add_67_carry_2_port
                           , YS => N48);
   add_67_U1_1_2 : HAX1 port map( A => n76, B => add_67_carry_2_port, YC => 
                           add_67_carry_3_port, YS => N49);
   add_67_U1_1_3 : HAX1 port map( A => n83, B => add_67_carry_3_port, YC => 
                           add_67_carry_4_port, YS => N50);
   r83_U1_1_1 : HAX1 port map( A => n78, B => writeptr_0_port, YC => 
                           r83_carry_2_port, YS => N32);
   r83_U1_1_2 : HAX1 port map( A => writeptr_2_port, B => r83_carry_2_port, YC 
                           => r83_carry_3_port, YS => N33);
   r83_U1_1_3 : HAX1 port map( A => writeptr_3_port, B => r83_carry_3_port, YC 
                           => r83_carry_4_port, YS => N34);
   BYTE_COUNT_reg_0_inst : DFFSR port map( D => N338, CLK => CLK, R => n98, S 
                           => n42, Q => BYTE_COUNT(0));
   BYTE_COUNT_reg_1_inst : DFFSR port map( D => N339, CLK => CLK, R => n98, S 
                           => n41, Q => BYTE_COUNT(1));
   BYTE_COUNT_reg_2_inst : DFFSR port map( D => N340, CLK => CLK, R => n98, S 
                           => n40, Q => BYTE_COUNT(2));
   readptr_reg_0_inst : DFFSR port map( D => N343, CLK => CLK, R => n98, S => 
                           n39, Q => readptr_0_port);
   readptr_reg_1_inst : DFFSR port map( D => N344, CLK => CLK, R => n98, S => 
                           n38, Q => readptr_1_port);
   BYTE_COUNT_reg_3_inst : DFFSR port map( D => N341, CLK => CLK, R => n98, S 
                           => n37, Q => BYTE_COUNT(3));
   readptr_reg_2_inst : DFFSR port map( D => N345, CLK => CLK, R => n98, S => 
                           n36, Q => readptr_2_port);
   BYTE_COUNT_reg_4_inst : DFFSR port map( D => N342, CLK => CLK, R => n98, S 
                           => n35, Q => BYTE_COUNT(4));
   readptr_reg_3_inst : DFFSR port map( D => N346, CLK => CLK, R => n98, S => 
                           n34_port, Q => readptr_3_port);
   writeptr_reg_4_inst : DFFSR port map( D => n1373, CLK => CLK, R => n98, S =>
                           n33_port, Q => writeptr_4_port);
   writeptr_reg_3_inst : DFFSR port map( D => n1374, CLK => CLK, R => n98, S =>
                           n32_port, Q => writeptr_3_port);
   writeptr_reg_2_inst : DFFSR port map( D => n1377, CLK => CLK, R => n98, S =>
                           n31, Q => writeptr_2_port);
   writeptr_reg_1_inst : DFFSR port map( D => n1376, CLK => CLK, R => n98, S =>
                           n30, Q => writeptr_1_port);
   writeptr_reg_0_inst : DFFSR port map( D => n1375, CLK => CLK, R => n98, S =>
                           n29, Q => writeptr_0_port);
   readptr_reg_4_inst : DFFSR port map( D => N347, CLK => CLK, R => n98, S => 
                           n28, Q => readptr_4_port);
   U3 : INVX4 port map( A => n55, Y => n124);
   U4 : OR2X1 port map( A => n152, B => n43_port, Y => n55);
   U5 : INVX4 port map( A => n50_port, Y => n119);
   U6 : OR2X1 port map( A => n147, B => n43_port, Y => n50_port);
   U7 : INVX4 port map( A => n56, Y => n114);
   U8 : OR2X1 port map( A => n193_port, B => n43_port, Y => n56);
   U9 : INVX4 port map( A => n49_port, Y => n435);
   U10 : OR2X1 port map( A => n244, B => n43_port, Y => n49_port);
   U11 : INVX4 port map( A => n57, Y => n461);
   U12 : OR2X1 port map( A => n156, B => n43_port, Y => n57);
   U13 : BUFX2 port map( A => n218, Y => n1);
   U14 : INVX2 port map( A => n77, Y => n78);
   U15 : INVX2 port map( A => n503, Y => n109);
   U16 : BUFX2 port map( A => n452, Y => n74);
   U17 : INVX2 port map( A => n23, Y => n73);
   U18 : INVX2 port map( A => n6, Y => n58);
   U19 : INVX2 port map( A => n11, Y => n59);
   U20 : INVX2 port map( A => n12, Y => n60);
   U21 : INVX2 port map( A => n14, Y => n72);
   U22 : INVX2 port map( A => n3, Y => n71);
   U23 : INVX2 port map( A => n4, Y => n70);
   U24 : INVX2 port map( A => n13, Y => n69);
   U25 : INVX2 port map( A => n24, Y => n65);
   U26 : INVX2 port map( A => n10, Y => n66);
   U27 : INVX2 port map( A => n15, Y => n67);
   U28 : INVX2 port map( A => n25, Y => n68);
   U29 : INVX2 port map( A => n7, Y => n64);
   U30 : INVX2 port map( A => n9, Y => n63);
   U31 : INVX2 port map( A => n26, Y => n62);
   U32 : INVX2 port map( A => n8, Y => n61);
   U33 : AND2X2 port map( A => n483, B => n361, Y => n2);
   U34 : OR2X2 port map( A => n1, B => n193_port, Y => n3);
   U35 : OR2X2 port map( A => n1, B => n147, Y => n4);
   U36 : AND2X2 port map( A => n496, B => n82, Y => n5);
   U37 : OR2X2 port map( A => n43_port, B => n184, Y => n6);
   U38 : OR2X2 port map( A => n44_port, B => n184, Y => n7);
   U39 : OR2X2 port map( A => n45_port, B => n152, Y => n8);
   U40 : OR2X2 port map( A => n44_port, B => n193_port, Y => n9);
   U41 : OR2X2 port map( A => n46_port, B => n161, Y => n10);
   U42 : OR2X2 port map( A => n1, B => n235, Y => n11);
   U43 : OR2X2 port map( A => n1, B => n244, Y => n12);
   U44 : OR2X2 port map( A => n1, B => n152, Y => n13);
   U45 : OR2X2 port map( A => n1, B => n184, Y => n14);
   U46 : OR2X2 port map( A => n46_port, B => n235, Y => n15);
   U47 : NAND2X1 port map( A => n253, B => n128, Y => n16);
   U48 : NAND2X1 port map( A => n253, B => n138, Y => n17);
   U49 : NAND2X1 port map( A => n253, B => n143, Y => n18);
   U50 : NAND2X1 port map( A => n253, B => n123, Y => n19);
   U51 : NAND2X1 port map( A => n253, B => n108, Y => n20);
   U52 : NAND2X1 port map( A => n253, B => n133, Y => n21);
   U53 : NAND2X1 port map( A => n253, B => n113, Y => n22);
   U54 : OR2X2 port map( A => n43_port, B => n235, Y => n23);
   U55 : OR2X2 port map( A => n45_port, B => n156, Y => n24);
   U56 : OR2X2 port map( A => n44_port, B => n244, Y => n25);
   U57 : OR2X2 port map( A => n45_port, B => n147, Y => n26);
   U58 : AND2X2 port map( A => n496, B => n83, Y => n27);
   U59 : INVX2 port map( A => n106, Y => n89);
   n28 <= '1';
   n29 <= '1';
   n30 <= '1';
   n31 <= '1';
   n32_port <= '1';
   n33_port <= '1';
   n34_port <= '1';
   n35 <= '1';
   n36 <= '1';
   n37 <= '1';
   n38 <= '1';
   n39 <= '1';
   n40 <= '1';
   n41 <= '1';
   n42 <= '1';
   U75 : BUFX2 port map( A => n183, Y => n43_port);
   U76 : NAND2X1 port map( A => n47, B => n27, Y => n183);
   U77 : NAND2X1 port map( A => n47, B => n5, Y => n218);
   U78 : OR2X2 port map( A => n156, B => n1, Y => n48_port);
   U79 : INVX2 port map( A => n148, Y => n139);
   U80 : INVX2 port map( A => n510, Y => n361);
   U81 : INVX2 port map( A => n511, Y => n165);
   U82 : BUFX2 port map( A => n286, Y => n44_port);
   U83 : BUFX2 port map( A => n286, Y => n45_port);
   U84 : BUFX2 port map( A => n286, Y => n46_port);
   U85 : NOR2X1 port map( A => n510, B => n483, Y => n47);
   U86 : INVX2 port map( A => writeptr_2_port, Y => n75);
   U87 : INVX2 port map( A => n89, Y => n88);
   U88 : INVX4 port map( A => n48_port, Y => n129);
   U89 : INVX4 port map( A => n54, Y => n134);
   U90 : XNOR2X1 port map( A => readptr_0_port, B => n81, Y => n519);
   U91 : INVX2 port map( A => RST, Y => n98);
   U92 : INVX2 port map( A => n82, Y => n83);
   U93 : INVX2 port map( A => n75, Y => n76);
   U94 : INVX2 port map( A => RCV_DATA(7), Y => n90);
   U95 : INVX2 port map( A => RCV_DATA(1), Y => n96);
   U96 : INVX2 port map( A => RCV_DATA(3), Y => n94);
   U97 : INVX2 port map( A => RCV_DATA(5), Y => n92);
   U98 : INVX2 port map( A => RCV_DATA(0), Y => n97);
   U99 : INVX2 port map( A => RCV_DATA(2), Y => n95);
   U100 : INVX2 port map( A => RCV_DATA(4), Y => n93);
   U101 : INVX2 port map( A => RCV_DATA(6), Y => n91);
   U102 : XNOR2X1 port map( A => readptr_4_port, B => n51_port, Y => n516);
   U103 : XNOR2X1 port map( A => r83_carry_4_port, B => writeptr_4_port, Y => 
                           n51_port);
   U104 : INVX2 port map( A => writeptr_3_port, Y => n82);
   U105 : BUFX2 port map( A => state, Y => n84);
   U106 : INVX1 port map( A => n80, Y => n81);
   U107 : INVX2 port map( A => writeptr_0_port, Y => n80);
   U108 : INVX1 port map( A => n47, Y => n52);
   U109 : INVX2 port map( A => n52, Y => n53);
   U110 : INVX1 port map( A => n77, Y => n79);
   U111 : INVX1 port map( A => writeptr_1_port, Y => n77);
   U112 : OR2X2 port map( A => n161, B => n1, Y => n54);
   U113 : INVX1 port map( A => RCV_OPCODE(0), Y => n106);
   U114 : AND2X2 port map( A => RCV_OPCODE(1), B => n89, Y => n483);
   U115 : INVX1 port map( A => RCV_OPCODE(1), Y => n87);
   U116 : INVX1 port map( A => RCV_OPCODE(1), Y => n86);
   U117 : INVX1 port map( A => RCV_OPCODE(1), Y => n85);
   U118 : AND2X2 port map( A => n478, B => n47, Y => n253);
   U119 : AND2X2 port map( A => n253, B => n118, Y => n394);
   U120 : AND2X2 port map( A => n818, B => n820, Y => n537);
   U121 : AND2X2 port map( A => n816, B => n820, Y => n536);
   U122 : AND2X2 port map( A => n818, B => n821, Y => n539);
   U123 : AND2X2 port map( A => n816, B => n821, Y => n538);
   U124 : AND2X2 port map( A => n832, B => n820, Y => n550);
   U125 : AND2X2 port map( A => n820, B => n831, Y => n549);
   U126 : AND2X2 port map( A => n821, B => n832, Y => n552);
   U127 : AND2X2 port map( A => n821, B => n831, Y => n551);
   U128 : AND2X2 port map( A => n843, B => n821, Y => n565);
   U129 : AND2X2 port map( A => n842, B => n821, Y => n564);
   U130 : AND2X2 port map( A => n843, B => n820, Y => n567);
   U131 : AND2X2 port map( A => n842, B => n820, Y => n566);
   U132 : AND2X2 port map( A => n853, B => n820, Y => n578);
   U133 : AND2X2 port map( A => n852, B => n820, Y => n577);
   U134 : AND2X2 port map( A => n853, B => n821, Y => n580);
   U135 : AND2X2 port map( A => n852, B => n821, Y => n579);
   U136 : OR2X1 port map( A => n823, B => n81, Y => sub_72_carry_1_port);
   U137 : XNOR2X1 port map( A => writeptr_0_port, B => n823, Y => N189);
   U138 : XOR2X1 port map( A => readptr_4_port, B => add_76_aco_carry_4_port, Y
                           => N337);
   U139 : AND2X1 port map( A => readptr_3_port, B => add_76_aco_carry_3_port, Y
                           => add_76_aco_carry_4_port);
   U140 : XOR2X1 port map( A => add_76_aco_carry_3_port, B => readptr_3_port, Y
                           => N336);
   U141 : AND2X1 port map( A => readptr_2_port, B => add_76_aco_carry_2_port, Y
                           => add_76_aco_carry_3_port);
   U142 : XOR2X1 port map( A => add_76_aco_carry_2_port, B => readptr_2_port, Y
                           => N335);
   U143 : AND2X1 port map( A => readptr_1_port, B => add_76_aco_carry_1_port, Y
                           => add_76_aco_carry_2_port);
   U144 : XOR2X1 port map( A => add_76_aco_carry_1_port, B => readptr_1_port, Y
                           => N334);
   U145 : AND2X1 port map( A => readptr_0_port, B => N195, Y => 
                           add_76_aco_carry_1_port);
   U146 : XOR2X1 port map( A => N195, B => readptr_0_port, Y => N333);
   U147 : NOR2X1 port map( A => n79, B => n81, Y => n100);
   U148 : AOI21X1 port map( A => n81, B => n79, C => n100, Y => n99);
   U149 : NAND2X1 port map( A => n100, B => n75, Y => n101);
   U150 : OAI21X1 port map( A => n100, B => n75, C => n101, Y => N44);
   U151 : XNOR2X1 port map( A => n83, B => n101, Y => N45);
   U152 : NOR2X1 port map( A => n83, B => n101, Y => n102);
   U153 : XOR2X1 port map( A => writeptr_4_port, B => n102, Y => N46);
   U154 : INVX2 port map( A => n99, Y => N43);
   U155 : XOR2X1 port map( A => add_67_carry_4_port, B => writeptr_4_port, Y =>
                           N51);
   U156 : MUX2X1 port map( B => n86, A => n104, S => n105, Y => n910);
   U157 : MUX2X1 port map( B => n88, A => n107, S => n105, Y => n911);
   U158 : AOI21X1 port map( A => n108, B => n109, C => n58, Y => n105);
   U159 : MUX2X1 port map( B => n85, A => n110, S => n111, Y => n912);
   U160 : MUX2X1 port map( B => n88, A => n112, S => n111, Y => n913);
   U161 : AOI21X1 port map( A => n109, B => n113, C => n114, Y => n111);
   U162 : MUX2X1 port map( B => n85, A => n115, S => n116, Y => n914);
   U163 : MUX2X1 port map( B => n88, A => n117, S => n116, Y => n915);
   U164 : AOI21X1 port map( A => n109, B => n118, C => n119, Y => n116);
   U165 : MUX2X1 port map( B => n85, A => n120, S => n121, Y => n916);
   U166 : MUX2X1 port map( B => n88, A => n122, S => n121, Y => n917);
   U167 : AOI21X1 port map( A => n109, B => n123, C => n124, Y => n121);
   U168 : MUX2X1 port map( B => n85, A => n125, S => n126, Y => n918);
   U169 : INVX1 port map( A => opcode_23_1_port, Y => n125);
   U170 : MUX2X1 port map( B => n88, A => n127, S => n126, Y => n919);
   U171 : AOI21X1 port map( A => n109, B => n128, C => n129, Y => n126);
   U172 : INVX1 port map( A => opcode_23_0_port, Y => n127);
   U173 : MUX2X1 port map( B => n85, A => n130, S => n131, Y => n920);
   U174 : INVX1 port map( A => opcode_22_1_port, Y => n130);
   U175 : MUX2X1 port map( B => n88, A => n132, S => n131, Y => n921);
   U176 : AOI21X1 port map( A => n109, B => n133, C => n134, Y => n131);
   U177 : INVX1 port map( A => opcode_22_0_port, Y => n132);
   U178 : MUX2X1 port map( B => n85, A => n135, S => n136, Y => n922);
   U179 : INVX1 port map( A => opcode_21_1_port, Y => n135);
   U180 : MUX2X1 port map( B => n88, A => n137, S => n136, Y => n923);
   U181 : AOI21X1 port map( A => n138, B => n139, C => n59, Y => n136);
   U182 : INVX1 port map( A => opcode_21_0_port, Y => n137);
   U183 : MUX2X1 port map( B => n85, A => n140, S => n141, Y => n924);
   U184 : INVX1 port map( A => opcode_20_1_port, Y => n140);
   U185 : MUX2X1 port map( B => n88, A => n142, S => n141, Y => n925);
   U186 : AOI21X1 port map( A => n143, B => n139, C => n60, Y => n141);
   U187 : INVX1 port map( A => opcode_20_0_port, Y => n142);
   U188 : INVX1 port map( A => n144, Y => n926);
   U189 : MUX2X1 port map( B => opcode_15_1_port, A => RCV_OPCODE(1), S => n145
                           , Y => n144);
   U190 : INVX1 port map( A => n146, Y => n927);
   U191 : MUX2X1 port map( B => opcode_15_0_port, A => RCV_OPCODE(0), S => n145
                           , Y => n146);
   U192 : OAI21X1 port map( A => n147, B => n148, C => n17, Y => n145);
   U193 : INVX1 port map( A => n149, Y => n928);
   U194 : MUX2X1 port map( B => opcode_14_1_port, A => RCV_OPCODE(1), S => n150
                           , Y => n149);
   U195 : INVX1 port map( A => n151, Y => n929);
   U196 : MUX2X1 port map( B => opcode_14_0_port, A => RCV_OPCODE(0), S => n150
                           , Y => n151);
   U197 : OAI21X1 port map( A => n152, B => n148, C => n18, Y => n150);
   U198 : MUX2X1 port map( B => n153, A => n87, S => n154, Y => n930);
   U199 : INVX1 port map( A => opcode_13_1_port, Y => n153);
   U200 : MUX2X1 port map( B => n155, A => n88, S => n154, Y => n931);
   U201 : OAI21X1 port map( A => n156, B => n157, C => n20, Y => n154);
   U202 : INVX1 port map( A => opcode_13_0_port, Y => n155);
   U203 : MUX2X1 port map( B => n158, A => n87, S => n159, Y => n932);
   U204 : INVX1 port map( A => opcode_12_1_port, Y => n158);
   U205 : MUX2X1 port map( B => n160, A => n88, S => n159, Y => n933);
   U206 : OAI21X1 port map( A => n161, B => n157, C => n22, Y => n159);
   U207 : INVX1 port map( A => opcode_12_0_port, Y => n160);
   U208 : MUX2X1 port map( B => n88, A => n162, S => n163, Y => n934);
   U209 : MUX2X1 port map( B => n85, A => n164, S => n163, Y => n935);
   U210 : AOI21X1 port map( A => n123, B => n165, C => n61, Y => n163);
   U211 : MUX2X1 port map( B => n88, A => n166, S => n167, Y => n936);
   U212 : MUX2X1 port map( B => n85, A => n168, S => n167, Y => n937);
   U213 : AOI21X1 port map( A => n118, B => n165, C => n62, Y => n167);
   U214 : MUX2X1 port map( B => n88, A => n169, S => n170, Y => n938);
   U215 : MUX2X1 port map( B => n85, A => n171, S => n170, Y => n939);
   U216 : AOI21X1 port map( A => n113, B => n165, C => n63, Y => n170);
   U217 : MUX2X1 port map( B => n88, A => n172, S => n173, Y => n940);
   U218 : MUX2X1 port map( B => n85, A => n174, S => n173, Y => n941);
   U219 : AOI21X1 port map( A => n108, B => n165, C => n64, Y => n173);
   U220 : MUX2X1 port map( B => n175, A => n90, S => n58, Y => n942);
   U221 : MUX2X1 port map( B => n176, A => n91, S => n58, Y => n943);
   U222 : MUX2X1 port map( B => n177, A => n92, S => n58, Y => n944);
   U223 : MUX2X1 port map( B => n178, A => n93, S => n58, Y => n945);
   U224 : MUX2X1 port map( B => n179, A => n94, S => n58, Y => n946);
   U225 : MUX2X1 port map( B => n180, A => n95, S => n58, Y => n947);
   U226 : MUX2X1 port map( B => n181, A => n96, S => n58, Y => n948);
   U227 : MUX2X1 port map( B => n182, A => n97, S => n58, Y => n949);
   U228 : MUX2X1 port map( B => n185, A => n90, S => n114, Y => n950);
   U229 : MUX2X1 port map( B => n186, A => n91, S => n114, Y => n951);
   U230 : MUX2X1 port map( B => n187, A => n92, S => n114, Y => n952);
   U231 : MUX2X1 port map( B => n188, A => n93, S => n114, Y => n953);
   U232 : MUX2X1 port map( B => n189_port, A => n94, S => n114, Y => n954);
   U233 : MUX2X1 port map( B => n190_port, A => n95, S => n114, Y => n955);
   U234 : MUX2X1 port map( B => n191_port, A => n96, S => n114, Y => n956);
   U235 : MUX2X1 port map( B => n192_port, A => n97, S => n114, Y => n957);
   U236 : MUX2X1 port map( B => n194, A => n90, S => n119, Y => n958);
   U237 : MUX2X1 port map( B => n195_port, A => n91, S => n119, Y => n959);
   U238 : MUX2X1 port map( B => n196, A => n92, S => n119, Y => n960);
   U239 : MUX2X1 port map( B => n197, A => n93, S => n119, Y => n961);
   U240 : MUX2X1 port map( B => n198, A => n94, S => n119, Y => n962);
   U241 : MUX2X1 port map( B => n199, A => n95, S => n119, Y => n963);
   U242 : MUX2X1 port map( B => n200, A => n96, S => n119, Y => n964);
   U243 : MUX2X1 port map( B => n201, A => n97, S => n119, Y => n965);
   U244 : MUX2X1 port map( B => n202, A => n90, S => n124, Y => n966);
   U245 : MUX2X1 port map( B => n203, A => n91, S => n124, Y => n967);
   U246 : MUX2X1 port map( B => n204, A => n92, S => n124, Y => n968);
   U247 : MUX2X1 port map( B => n205, A => n93, S => n124, Y => n969);
   U248 : MUX2X1 port map( B => n206, A => n94, S => n124, Y => n970);
   U249 : MUX2X1 port map( B => n207, A => n95, S => n124, Y => n971);
   U250 : MUX2X1 port map( B => n208, A => n96, S => n124, Y => n972);
   U251 : MUX2X1 port map( B => n209, A => n97, S => n124, Y => n973);
   U252 : MUX2X1 port map( B => n210, A => n90, S => n129, Y => n974);
   U253 : INVX1 port map( A => memory_23_7_port, Y => n210);
   U254 : MUX2X1 port map( B => n211, A => n91, S => n129, Y => n975);
   U255 : INVX1 port map( A => memory_23_6_port, Y => n211);
   U256 : MUX2X1 port map( B => n212, A => n92, S => n129, Y => n976);
   U257 : INVX1 port map( A => memory_23_5_port, Y => n212);
   U258 : MUX2X1 port map( B => n213, A => n93, S => n129, Y => n977);
   U259 : INVX1 port map( A => memory_23_4_port, Y => n213);
   U260 : MUX2X1 port map( B => n214, A => n94, S => n129, Y => n978);
   U261 : INVX1 port map( A => memory_23_3_port, Y => n214);
   U262 : MUX2X1 port map( B => n215, A => n95, S => n129, Y => n979);
   U263 : INVX1 port map( A => memory_23_2_port, Y => n215);
   U264 : MUX2X1 port map( B => n216, A => n96, S => n129, Y => n980);
   U265 : INVX1 port map( A => memory_23_1_port, Y => n216);
   U266 : MUX2X1 port map( B => n217, A => n97, S => n129, Y => n981);
   U267 : INVX1 port map( A => memory_23_0_port, Y => n217);
   U268 : MUX2X1 port map( B => n219, A => n90, S => n134, Y => n982);
   U269 : INVX1 port map( A => memory_22_7_port, Y => n219);
   U270 : MUX2X1 port map( B => n220, A => n91, S => n134, Y => n983);
   U271 : INVX1 port map( A => memory_22_6_port, Y => n220);
   U272 : MUX2X1 port map( B => n221, A => n92, S => n134, Y => n984);
   U273 : INVX1 port map( A => memory_22_5_port, Y => n221);
   U274 : MUX2X1 port map( B => n222, A => n93, S => n134, Y => n985);
   U275 : INVX1 port map( A => memory_22_4_port, Y => n222);
   U276 : MUX2X1 port map( B => n223, A => n94, S => n134, Y => n986);
   U277 : INVX1 port map( A => memory_22_3_port, Y => n223);
   U278 : MUX2X1 port map( B => n224, A => n95, S => n134, Y => n987);
   U279 : INVX1 port map( A => memory_22_2_port, Y => n224);
   U280 : MUX2X1 port map( B => n225, A => n96, S => n134, Y => n988);
   U281 : INVX1 port map( A => memory_22_1_port, Y => n225);
   U282 : MUX2X1 port map( B => n226, A => n97, S => n134, Y => n989);
   U283 : INVX1 port map( A => memory_22_0_port, Y => n226);
   U284 : MUX2X1 port map( B => n227, A => n90, S => n59, Y => n990);
   U285 : INVX1 port map( A => memory_21_7_port, Y => n227);
   U286 : MUX2X1 port map( B => n228, A => n91, S => n59, Y => n991);
   U287 : INVX1 port map( A => memory_21_6_port, Y => n228);
   U288 : MUX2X1 port map( B => n229, A => n92, S => n59, Y => n992);
   U289 : INVX1 port map( A => memory_21_5_port, Y => n229);
   U290 : MUX2X1 port map( B => n230, A => n93, S => n59, Y => n993);
   U291 : INVX1 port map( A => memory_21_4_port, Y => n230);
   U292 : MUX2X1 port map( B => n231, A => n94, S => n59, Y => n994);
   U293 : INVX1 port map( A => memory_21_3_port, Y => n231);
   U294 : MUX2X1 port map( B => n232, A => n95, S => n59, Y => n995);
   U295 : INVX1 port map( A => memory_21_2_port, Y => n232);
   U296 : MUX2X1 port map( B => n233, A => n96, S => n59, Y => n996);
   U297 : INVX1 port map( A => memory_21_1_port, Y => n233);
   U298 : MUX2X1 port map( B => n234, A => n97, S => n59, Y => n997);
   U299 : INVX1 port map( A => memory_21_0_port, Y => n234);
   U300 : MUX2X1 port map( B => n236, A => n90, S => n60, Y => n998);
   U301 : INVX1 port map( A => memory_20_7_port, Y => n236);
   U302 : MUX2X1 port map( B => n237, A => n91, S => n60, Y => n999);
   U303 : INVX1 port map( A => memory_20_6_port, Y => n237);
   U304 : MUX2X1 port map( B => n238, A => n92, S => n60, Y => n1000);
   U305 : INVX1 port map( A => memory_20_5_port, Y => n238);
   U306 : MUX2X1 port map( B => n239, A => n93, S => n60, Y => n1001);
   U307 : INVX1 port map( A => memory_20_4_port, Y => n239);
   U308 : MUX2X1 port map( B => n240, A => n94, S => n60, Y => n1002);
   U309 : INVX1 port map( A => memory_20_3_port, Y => n240);
   U310 : MUX2X1 port map( B => n241, A => n95, S => n60, Y => n1003);
   U311 : INVX1 port map( A => memory_20_2_port, Y => n241);
   U312 : MUX2X1 port map( B => n242, A => n96, S => n60, Y => n1004);
   U313 : INVX1 port map( A => memory_20_1_port, Y => n242);
   U314 : MUX2X1 port map( B => n243, A => n97, S => n60, Y => n1005);
   U315 : INVX1 port map( A => memory_20_0_port, Y => n243);
   U316 : MUX2X1 port map( B => n90, A => n245, S => n17, Y => n1006);
   U317 : INVX1 port map( A => memory_15_7_port, Y => n245);
   U318 : MUX2X1 port map( B => n91, A => n246, S => n17, Y => n1007);
   U319 : INVX1 port map( A => memory_15_6_port, Y => n246);
   U320 : MUX2X1 port map( B => n92, A => n247, S => n17, Y => n1008);
   U321 : INVX1 port map( A => memory_15_5_port, Y => n247);
   U322 : MUX2X1 port map( B => n93, A => n248, S => n17, Y => n1009);
   U323 : INVX1 port map( A => memory_15_4_port, Y => n248);
   U324 : MUX2X1 port map( B => n94, A => n249, S => n17, Y => n1010);
   U325 : INVX1 port map( A => memory_15_3_port, Y => n249);
   U326 : MUX2X1 port map( B => n95, A => n250, S => n17, Y => n1011);
   U327 : INVX1 port map( A => memory_15_2_port, Y => n250);
   U328 : MUX2X1 port map( B => n96, A => n251, S => n17, Y => n1012);
   U329 : INVX1 port map( A => memory_15_1_port, Y => n251);
   U330 : MUX2X1 port map( B => n97, A => n252, S => n17, Y => n1013);
   U331 : INVX1 port map( A => memory_15_0_port, Y => n252);
   U332 : MUX2X1 port map( B => n90, A => n254, S => n18, Y => n1014);
   U333 : INVX1 port map( A => memory_14_7_port, Y => n254);
   U334 : MUX2X1 port map( B => n91, A => n255, S => n18, Y => n1015);
   U335 : INVX1 port map( A => memory_14_6_port, Y => n255);
   U336 : MUX2X1 port map( B => n92, A => n256, S => n18, Y => n1016);
   U337 : INVX1 port map( A => memory_14_5_port, Y => n256);
   U338 : MUX2X1 port map( B => n93, A => n257, S => n18, Y => n1017);
   U339 : INVX1 port map( A => memory_14_4_port, Y => n257);
   U340 : MUX2X1 port map( B => n94, A => n258, S => n18, Y => n1018);
   U341 : INVX1 port map( A => memory_14_3_port, Y => n258);
   U342 : MUX2X1 port map( B => n95, A => n259, S => n18, Y => n1019);
   U343 : INVX1 port map( A => memory_14_2_port, Y => n259);
   U344 : MUX2X1 port map( B => n96, A => n260, S => n18, Y => n1020);
   U345 : INVX1 port map( A => memory_14_1_port, Y => n260);
   U346 : MUX2X1 port map( B => n97, A => n261, S => n18, Y => n1021);
   U347 : INVX1 port map( A => memory_14_0_port, Y => n261);
   U348 : MUX2X1 port map( B => n90, A => n262, S => n20, Y => n1022);
   U349 : INVX1 port map( A => memory_13_7_port, Y => n262);
   U350 : MUX2X1 port map( B => n91, A => n263, S => n20, Y => n1023);
   U351 : INVX1 port map( A => memory_13_6_port, Y => n263);
   U352 : MUX2X1 port map( B => n92, A => n264, S => n20, Y => n1024);
   U353 : INVX1 port map( A => memory_13_5_port, Y => n264);
   U354 : MUX2X1 port map( B => n93, A => n265, S => n20, Y => n1025);
   U355 : INVX1 port map( A => memory_13_4_port, Y => n265);
   U356 : MUX2X1 port map( B => n94, A => n266, S => n20, Y => n1026);
   U357 : INVX1 port map( A => memory_13_3_port, Y => n266);
   U358 : MUX2X1 port map( B => n95, A => n267, S => n20, Y => n1027);
   U359 : INVX1 port map( A => memory_13_2_port, Y => n267);
   U360 : MUX2X1 port map( B => n96, A => n268, S => n20, Y => n1028);
   U361 : INVX1 port map( A => memory_13_1_port, Y => n268);
   U362 : MUX2X1 port map( B => n97, A => n269, S => n20, Y => n1029);
   U363 : INVX1 port map( A => memory_13_0_port, Y => n269);
   U364 : MUX2X1 port map( B => n90, A => n270, S => n22, Y => n1064);
   U365 : INVX1 port map( A => memory_12_7_port, Y => n270);
   U366 : MUX2X1 port map( B => n91, A => n271, S => n22, Y => n1065);
   U367 : INVX1 port map( A => memory_12_6_port, Y => n271);
   U368 : MUX2X1 port map( B => n92, A => n272, S => n22, Y => n1066);
   U369 : INVX1 port map( A => memory_12_5_port, Y => n272);
   U370 : MUX2X1 port map( B => n93, A => n273, S => n22, Y => n1067);
   U371 : INVX1 port map( A => memory_12_4_port, Y => n273);
   U372 : MUX2X1 port map( B => n94, A => n274, S => n22, Y => n1068);
   U373 : INVX1 port map( A => memory_12_3_port, Y => n274);
   U374 : MUX2X1 port map( B => n95, A => n275, S => n22, Y => n1069);
   U375 : INVX1 port map( A => memory_12_2_port, Y => n275);
   U376 : MUX2X1 port map( B => n96, A => n276, S => n22, Y => n1070);
   U377 : INVX1 port map( A => memory_12_1_port, Y => n276);
   U378 : MUX2X1 port map( B => n97, A => n277, S => n22, Y => n1071);
   U379 : INVX1 port map( A => memory_12_0_port, Y => n277);
   U380 : MUX2X1 port map( B => n278, A => n97, S => n61, Y => n1168);
   U381 : MUX2X1 port map( B => n279, A => n96, S => n61, Y => n1169);
   U382 : MUX2X1 port map( B => n280, A => n95, S => n61, Y => n1170);
   U383 : MUX2X1 port map( B => n281, A => n94, S => n61, Y => n1171);
   U384 : MUX2X1 port map( B => n282, A => n93, S => n61, Y => n1172);
   U385 : MUX2X1 port map( B => n283, A => n92, S => n61, Y => n1173);
   U386 : MUX2X1 port map( B => n284, A => n91, S => n61, Y => n1174);
   U387 : MUX2X1 port map( B => n285, A => n90, S => n61, Y => n1175);
   U388 : MUX2X1 port map( B => n287, A => n97, S => n62, Y => n1176);
   U389 : MUX2X1 port map( B => n288, A => n96, S => n62, Y => n1177);
   U390 : MUX2X1 port map( B => n289, A => n95, S => n62, Y => n1178);
   U391 : MUX2X1 port map( B => n290, A => n94, S => n62, Y => n1179);
   U392 : MUX2X1 port map( B => n291, A => n93, S => n62, Y => n1180);
   U393 : MUX2X1 port map( B => n292, A => n92, S => n62, Y => n1181);
   U394 : MUX2X1 port map( B => n293, A => n91, S => n62, Y => n1182);
   U395 : MUX2X1 port map( B => n294, A => n90, S => n62, Y => n1183);
   U396 : MUX2X1 port map( B => n295, A => n97, S => n63, Y => n1184);
   U397 : MUX2X1 port map( B => n296, A => n96, S => n63, Y => n1185);
   U398 : MUX2X1 port map( B => n297, A => n95, S => n63, Y => n1186);
   U399 : MUX2X1 port map( B => n298, A => n94, S => n63, Y => n1187);
   U400 : MUX2X1 port map( B => n299, A => n93, S => n63, Y => n1188);
   U401 : MUX2X1 port map( B => n300, A => n92, S => n63, Y => n1189);
   U402 : MUX2X1 port map( B => n301, A => n91, S => n63, Y => n1190);
   U403 : MUX2X1 port map( B => n302, A => n90, S => n63, Y => n1191);
   U404 : MUX2X1 port map( B => n303, A => n97, S => n64, Y => n1192);
   U405 : MUX2X1 port map( B => n304, A => n96, S => n64, Y => n1193);
   U406 : MUX2X1 port map( B => n305, A => n95, S => n64, Y => n1194);
   U407 : MUX2X1 port map( B => n306, A => n94, S => n64, Y => n1195);
   U408 : MUX2X1 port map( B => n307, A => n93, S => n64, Y => n1196);
   U409 : MUX2X1 port map( B => n308, A => n92, S => n64, Y => n1197);
   U410 : MUX2X1 port map( B => n309, A => n91, S => n64, Y => n1198);
   U411 : MUX2X1 port map( B => n310, A => n90, S => n64, Y => n1199);
   U412 : MUX2X1 port map( B => n311, A => n312, S => RST, Y => n1200);
   U413 : INVX1 port map( A => FULL_port, Y => n312);
   U414 : MUX2X1 port map( B => n313, A => n314, S => RST, Y => n1201);
   U415 : INVX1 port map( A => EMPTY_port, Y => n314);
   U416 : MUX2X1 port map( B => n88, A => n315, S => n316, Y => n1332);
   U417 : INVX1 port map( A => opcode_7_0_port, Y => n315);
   U418 : MUX2X1 port map( B => n85, A => n317, S => n316, Y => n1333);
   U419 : AOI21X1 port map( A => n128, B => n318, C => n65, Y => n316);
   U420 : INVX1 port map( A => opcode_7_1_port, Y => n317);
   U421 : MUX2X1 port map( B => n319, A => n97, S => n65, Y => n1334);
   U422 : INVX1 port map( A => memory_7_0_port, Y => n319);
   U423 : MUX2X1 port map( B => n320, A => n96, S => n65, Y => n1335);
   U424 : INVX1 port map( A => memory_7_1_port, Y => n320);
   U425 : MUX2X1 port map( B => n321, A => n95, S => n65, Y => n1336);
   U426 : INVX1 port map( A => memory_7_2_port, Y => n321);
   U427 : MUX2X1 port map( B => n322, A => n94, S => n65, Y => n1337);
   U428 : INVX1 port map( A => memory_7_3_port, Y => n322);
   U429 : MUX2X1 port map( B => n323, A => n93, S => n65, Y => n1338);
   U430 : INVX1 port map( A => memory_7_4_port, Y => n323);
   U431 : MUX2X1 port map( B => n324, A => n92, S => n65, Y => n1339);
   U432 : INVX1 port map( A => memory_7_5_port, Y => n324);
   U433 : MUX2X1 port map( B => n325, A => n91, S => n65, Y => n1340);
   U434 : INVX1 port map( A => memory_7_6_port, Y => n325);
   U435 : MUX2X1 port map( B => n326, A => n90, S => n65, Y => n1341);
   U436 : INVX1 port map( A => memory_7_7_port, Y => n326);
   U437 : MUX2X1 port map( B => n88, A => n327, S => n328, Y => n1342);
   U438 : INVX1 port map( A => opcode_6_0_port, Y => n327);
   U439 : MUX2X1 port map( B => n86, A => n329, S => n328, Y => n1343);
   U440 : AOI21X1 port map( A => n133, B => n318, C => n66, Y => n328);
   U441 : INVX1 port map( A => n157, Y => n318);
   U442 : INVX1 port map( A => opcode_6_1_port, Y => n329);
   U443 : MUX2X1 port map( B => n330, A => n97, S => n66, Y => n1344);
   U444 : INVX1 port map( A => memory_6_0_port, Y => n330);
   U445 : MUX2X1 port map( B => n331, A => n96, S => n66, Y => n1345);
   U446 : INVX1 port map( A => memory_6_1_port, Y => n331);
   U447 : MUX2X1 port map( B => n332, A => n95, S => n66, Y => n1346);
   U448 : INVX1 port map( A => memory_6_2_port, Y => n332);
   U449 : MUX2X1 port map( B => n333_port, A => n94, S => n66, Y => n1347);
   U450 : INVX1 port map( A => memory_6_3_port, Y => n333_port);
   U451 : MUX2X1 port map( B => n334_port, A => n93, S => n66, Y => n1348);
   U452 : INVX1 port map( A => memory_6_4_port, Y => n334_port);
   U453 : MUX2X1 port map( B => n335_port, A => n92, S => n66, Y => n1349);
   U454 : INVX1 port map( A => memory_6_5_port, Y => n335_port);
   U455 : MUX2X1 port map( B => n336_port, A => n91, S => n66, Y => n1350);
   U456 : INVX1 port map( A => memory_6_6_port, Y => n336_port);
   U457 : MUX2X1 port map( B => n337_port, A => n90, S => n66, Y => n1351);
   U458 : INVX1 port map( A => memory_6_7_port, Y => n337_port);
   U459 : MUX2X1 port map( B => n106, A => n338_port, S => n339_port, Y => 
                           n1352);
   U460 : INVX1 port map( A => opcode_5_0_port, Y => n338_port);
   U461 : MUX2X1 port map( B => n86, A => n340_port, S => n339_port, Y => n1353
                           );
   U462 : AOI21X1 port map( A => n138, B => n165, C => n67, Y => n339_port);
   U463 : INVX1 port map( A => opcode_5_1_port, Y => n340_port);
   U464 : MUX2X1 port map( B => n341_port, A => n97, S => n67, Y => n1354);
   U465 : INVX1 port map( A => memory_5_0_port, Y => n341_port);
   U466 : MUX2X1 port map( B => n342_port, A => n96, S => n67, Y => n1355);
   U467 : INVX1 port map( A => memory_5_1_port, Y => n342_port);
   U468 : MUX2X1 port map( B => n343_port, A => n95, S => n67, Y => n1356);
   U469 : INVX1 port map( A => memory_5_2_port, Y => n343_port);
   U470 : MUX2X1 port map( B => n344_port, A => n94, S => n67, Y => n1357);
   U471 : INVX1 port map( A => memory_5_3_port, Y => n344_port);
   U472 : MUX2X1 port map( B => n345_port, A => n93, S => n67, Y => n1358);
   U473 : INVX1 port map( A => memory_5_4_port, Y => n345_port);
   U474 : MUX2X1 port map( B => n346_port, A => n92, S => n67, Y => n1359);
   U475 : INVX1 port map( A => memory_5_5_port, Y => n346_port);
   U476 : MUX2X1 port map( B => n347_port, A => n91, S => n67, Y => n1360);
   U477 : INVX1 port map( A => memory_5_6_port, Y => n347_port);
   U478 : MUX2X1 port map( B => n348, A => n90, S => n67, Y => n1361);
   U479 : INVX1 port map( A => memory_5_7_port, Y => n348);
   U480 : MUX2X1 port map( B => n88, A => n349, S => n350, Y => n1362);
   U481 : INVX1 port map( A => opcode_4_0_port, Y => n349);
   U482 : MUX2X1 port map( B => n86, A => n351, S => n350, Y => n1363);
   U483 : AOI21X1 port map( A => n143, B => n165, C => n68, Y => n350);
   U484 : INVX1 port map( A => opcode_4_1_port, Y => n351);
   U485 : MUX2X1 port map( B => n352, A => n97, S => n68, Y => n1364);
   U486 : INVX1 port map( A => memory_4_0_port, Y => n352);
   U487 : MUX2X1 port map( B => n353, A => n96, S => n68, Y => n1365);
   U488 : INVX1 port map( A => memory_4_1_port, Y => n353);
   U489 : MUX2X1 port map( B => n354, A => n95, S => n68, Y => n1366);
   U490 : INVX1 port map( A => memory_4_2_port, Y => n354);
   U491 : MUX2X1 port map( B => n355, A => n94, S => n68, Y => n1367);
   U492 : INVX1 port map( A => memory_4_3_port, Y => n355);
   U493 : MUX2X1 port map( B => n356, A => n93, S => n68, Y => n1368);
   U494 : INVX1 port map( A => memory_4_4_port, Y => n356);
   U495 : MUX2X1 port map( B => n357, A => n92, S => n68, Y => n1369);
   U496 : INVX1 port map( A => memory_4_5_port, Y => n357);
   U497 : MUX2X1 port map( B => n358, A => n91, S => n68, Y => n1370);
   U498 : INVX1 port map( A => memory_4_6_port, Y => n358);
   U499 : MUX2X1 port map( B => n359, A => n90, S => n68, Y => n1371);
   U500 : NAND3X1 port map( A => n47, B => n82, C => n360, Y => n286);
   U501 : INVX1 port map( A => memory_4_7_port, Y => n359);
   U502 : OAI21X1 port map( A => n361, B => n362, C => n363, Y => n1373);
   U503 : AOI22X1 port map( A => N51, B => n53, C => N46, D => n2, Y => n363);
   U504 : OAI21X1 port map( A => n361, B => n82, C => n364, Y => n1374);
   U505 : AOI22X1 port map( A => N50, B => n53, C => N45, D => n2, Y => n364);
   U506 : OAI21X1 port map( A => n361, B => n80, C => n365, Y => n1375);
   U507 : AOI22X1 port map( A => n80, B => n53, C => n80, D => n2, Y => n365);
   U508 : OAI21X1 port map( A => n361, B => n366, C => n367, Y => n1376);
   U509 : AOI22X1 port map( A => N48, B => n53, C => N43, D => n2, Y => n367);
   U510 : OAI21X1 port map( A => n361, B => n75, C => n368, Y => n1377);
   U511 : AOI22X1 port map( A => N49, B => n53, C => N44, D => n2, Y => n368);
   U512 : MUX2X1 port map( B => n90, A => n369, S => n21, Y => n1202);
   U513 : MUX2X1 port map( B => n91, A => n370, S => n21, Y => n1203);
   U514 : MUX2X1 port map( B => n92, A => n371, S => n21, Y => n1204);
   U515 : MUX2X1 port map( B => n93, A => n372, S => n21, Y => n1205);
   U516 : MUX2X1 port map( B => n94, A => n373, S => n21, Y => n1206);
   U517 : MUX2X1 port map( B => n95, A => n374, S => n21, Y => n1207);
   U518 : MUX2X1 port map( B => n96, A => n375, S => n21, Y => n1208);
   U519 : MUX2X1 port map( B => n97, A => n376, S => n21, Y => n1209);
   U520 : MUX2X1 port map( B => n90, A => n377, S => n16, Y => n1210);
   U521 : MUX2X1 port map( B => n91, A => n378, S => n16, Y => n1211);
   U522 : MUX2X1 port map( B => n92, A => n379, S => n16, Y => n1212);
   U523 : MUX2X1 port map( B => n93, A => n380, S => n16, Y => n1213);
   U524 : MUX2X1 port map( B => n94, A => n381, S => n16, Y => n1214);
   U525 : MUX2X1 port map( B => n95, A => n382, S => n16, Y => n1215);
   U526 : MUX2X1 port map( B => n96, A => n383, S => n16, Y => n1216);
   U527 : MUX2X1 port map( B => n97, A => n384, S => n16, Y => n1217);
   U528 : MUX2X1 port map( B => n90, A => n385, S => n19, Y => n1218);
   U529 : MUX2X1 port map( B => n91, A => n386, S => n19, Y => n1219);
   U530 : MUX2X1 port map( B => n92, A => n387, S => n19, Y => n1220);
   U531 : MUX2X1 port map( B => n93, A => n388, S => n19, Y => n1221);
   U532 : MUX2X1 port map( B => n94, A => n389, S => n19, Y => n1222);
   U533 : MUX2X1 port map( B => n95, A => n390, S => n19, Y => n1223);
   U534 : MUX2X1 port map( B => n96, A => n391, S => n19, Y => n1224);
   U535 : MUX2X1 port map( B => n97, A => n392, S => n19, Y => n1225);
   U536 : MUX2X1 port map( B => n393, A => n90, S => n394, Y => n1226);
   U537 : MUX2X1 port map( B => n395, A => n91, S => n394, Y => n1227);
   U538 : MUX2X1 port map( B => n396, A => n92, S => n394, Y => n1228);
   U539 : MUX2X1 port map( B => n397, A => n93, S => n394, Y => n1229);
   U540 : MUX2X1 port map( B => n398, A => n94, S => n394, Y => n1230);
   U541 : MUX2X1 port map( B => n399, A => n95, S => n394, Y => n1231);
   U542 : MUX2X1 port map( B => n400, A => n96, S => n394, Y => n1232);
   U543 : MUX2X1 port map( B => n401, A => n97, S => n394, Y => n1233);
   U544 : MUX2X1 port map( B => n402, A => n90, S => n69, Y => n1234);
   U545 : MUX2X1 port map( B => n403, A => n91, S => n69, Y => n1235);
   U546 : MUX2X1 port map( B => n404, A => n92, S => n69, Y => n1236);
   U547 : MUX2X1 port map( B => n405, A => n93, S => n69, Y => n1237);
   U548 : MUX2X1 port map( B => n406, A => n94, S => n69, Y => n1238);
   U549 : MUX2X1 port map( B => n407, A => n95, S => n69, Y => n1239);
   U550 : MUX2X1 port map( B => n408, A => n96, S => n69, Y => n1240);
   U551 : MUX2X1 port map( B => n409, A => n97, S => n69, Y => n1241);
   U552 : MUX2X1 port map( B => n410, A => n90, S => n70, Y => n1242);
   U553 : MUX2X1 port map( B => n411, A => n91, S => n70, Y => n1243);
   U554 : MUX2X1 port map( B => n412, A => n92, S => n70, Y => n1244);
   U555 : MUX2X1 port map( B => n413, A => n93, S => n70, Y => n1245);
   U556 : MUX2X1 port map( B => n414, A => n94, S => n70, Y => n1246);
   U557 : MUX2X1 port map( B => n415, A => n95, S => n70, Y => n1247);
   U558 : MUX2X1 port map( B => n416, A => n96, S => n70, Y => n1248);
   U559 : MUX2X1 port map( B => n417, A => n97, S => n70, Y => n1249);
   U560 : MUX2X1 port map( B => n418, A => n90, S => n71, Y => n1250);
   U561 : MUX2X1 port map( B => n419, A => n91, S => n71, Y => n1251);
   U562 : MUX2X1 port map( B => n420, A => n92, S => n71, Y => n1252);
   U563 : MUX2X1 port map( B => n421, A => n93, S => n71, Y => n1253);
   U564 : MUX2X1 port map( B => n422, A => n94, S => n71, Y => n1254);
   U565 : MUX2X1 port map( B => n423, A => n95, S => n71, Y => n1255);
   U566 : MUX2X1 port map( B => n424, A => n96, S => n71, Y => n1256);
   U567 : MUX2X1 port map( B => n425, A => n97, S => n71, Y => n1257);
   U568 : MUX2X1 port map( B => n426, A => n90, S => n72, Y => n1258);
   U569 : MUX2X1 port map( B => n427, A => n91, S => n72, Y => n1259);
   U570 : MUX2X1 port map( B => n428, A => n92, S => n72, Y => n1260);
   U571 : MUX2X1 port map( B => n429, A => n93, S => n72, Y => n1261);
   U572 : MUX2X1 port map( B => n430, A => n94, S => n72, Y => n1262);
   U573 : MUX2X1 port map( B => n431, A => n95, S => n72, Y => n1263);
   U574 : MUX2X1 port map( B => n432, A => n96, S => n72, Y => n1264);
   U575 : MUX2X1 port map( B => n433, A => n97, S => n72, Y => n1265);
   U576 : INVX1 port map( A => n434, Y => n1266);
   U577 : MUX2X1 port map( B => memory_28_7_port, A => RCV_DATA(7), S => n435, 
                           Y => n434);
   U578 : INVX1 port map( A => n436, Y => n1267);
   U579 : MUX2X1 port map( B => memory_28_6_port, A => RCV_DATA(6), S => n435, 
                           Y => n436);
   U580 : INVX1 port map( A => n437, Y => n1268);
   U581 : MUX2X1 port map( B => memory_28_5_port, A => RCV_DATA(5), S => n435, 
                           Y => n437);
   U582 : INVX1 port map( A => n438, Y => n1269);
   U583 : MUX2X1 port map( B => memory_28_4_port, A => RCV_DATA(4), S => n435, 
                           Y => n438);
   U584 : INVX1 port map( A => n439, Y => n1270);
   U585 : MUX2X1 port map( B => memory_28_3_port, A => RCV_DATA(3), S => n435, 
                           Y => n439);
   U586 : INVX1 port map( A => n440, Y => n1271);
   U587 : MUX2X1 port map( B => memory_28_2_port, A => RCV_DATA(2), S => n435, 
                           Y => n440);
   U588 : INVX1 port map( A => n441, Y => n1272);
   U589 : MUX2X1 port map( B => memory_28_1_port, A => RCV_DATA(1), S => n435, 
                           Y => n441);
   U590 : INVX1 port map( A => n442, Y => n1273);
   U591 : MUX2X1 port map( B => memory_28_0_port, A => RCV_DATA(0), S => n435, 
                           Y => n442);
   U592 : INVX1 port map( A => n443, Y => n1274);
   U593 : MUX2X1 port map( B => memory_29_7_port, A => RCV_DATA(7), S => n73, Y
                           => n443);
   U594 : INVX1 port map( A => n444, Y => n1275);
   U595 : MUX2X1 port map( B => memory_29_6_port, A => RCV_DATA(6), S => n73, Y
                           => n444);
   U596 : INVX1 port map( A => n445, Y => n1276);
   U597 : MUX2X1 port map( B => memory_29_5_port, A => RCV_DATA(5), S => n73, Y
                           => n445);
   U598 : INVX1 port map( A => n446, Y => n1277);
   U599 : MUX2X1 port map( B => memory_29_4_port, A => RCV_DATA(4), S => n73, Y
                           => n446);
   U600 : INVX1 port map( A => n447, Y => n1278);
   U601 : MUX2X1 port map( B => memory_29_3_port, A => RCV_DATA(3), S => n73, Y
                           => n447);
   U602 : INVX1 port map( A => n448, Y => n1279);
   U603 : MUX2X1 port map( B => memory_29_2_port, A => RCV_DATA(2), S => n73, Y
                           => n448);
   U604 : INVX1 port map( A => n449, Y => n1280);
   U605 : MUX2X1 port map( B => memory_29_1_port, A => RCV_DATA(1), S => n73, Y
                           => n449);
   U606 : INVX1 port map( A => n450, Y => n1281);
   U607 : MUX2X1 port map( B => memory_29_0_port, A => RCV_DATA(0), S => n73, Y
                           => n450);
   U608 : INVX1 port map( A => n451, Y => n1282);
   U609 : MUX2X1 port map( B => memory_30_7_port, A => RCV_DATA(7), S => n74, Y
                           => n451);
   U610 : INVX1 port map( A => n453, Y => n1283);
   U611 : MUX2X1 port map( B => memory_30_6_port, A => RCV_DATA(6), S => n74, Y
                           => n453);
   U612 : INVX1 port map( A => n454, Y => n1284);
   U613 : MUX2X1 port map( B => memory_30_5_port, A => RCV_DATA(5), S => n74, Y
                           => n454);
   U614 : INVX1 port map( A => n455, Y => n1285);
   U615 : MUX2X1 port map( B => memory_30_4_port, A => RCV_DATA(4), S => n74, Y
                           => n455);
   U616 : INVX1 port map( A => n456, Y => n1286);
   U617 : MUX2X1 port map( B => memory_30_3_port, A => RCV_DATA(3), S => n74, Y
                           => n456);
   U618 : INVX1 port map( A => n457, Y => n1287);
   U619 : MUX2X1 port map( B => memory_30_2_port, A => RCV_DATA(2), S => n74, Y
                           => n457);
   U620 : INVX1 port map( A => n458, Y => n1288);
   U621 : MUX2X1 port map( B => memory_30_1_port, A => RCV_DATA(1), S => n74, Y
                           => n458);
   U622 : INVX1 port map( A => n459, Y => n1289);
   U623 : MUX2X1 port map( B => memory_30_0_port, A => RCV_DATA(0), S => n74, Y
                           => n459);
   U624 : INVX1 port map( A => n460, Y => n1290);
   U625 : MUX2X1 port map( B => memory_31_7_port, A => RCV_DATA(7), S => n461, 
                           Y => n460);
   U626 : INVX1 port map( A => n462, Y => n1291);
   U627 : MUX2X1 port map( B => memory_31_6_port, A => RCV_DATA(6), S => n461, 
                           Y => n462);
   U628 : INVX1 port map( A => n463, Y => n1292);
   U629 : MUX2X1 port map( B => memory_31_5_port, A => RCV_DATA(5), S => n461, 
                           Y => n463);
   U630 : INVX1 port map( A => n464, Y => n1293);
   U631 : MUX2X1 port map( B => memory_31_4_port, A => RCV_DATA(4), S => n461, 
                           Y => n464);
   U632 : INVX1 port map( A => n465, Y => n1294);
   U633 : MUX2X1 port map( B => memory_31_3_port, A => RCV_DATA(3), S => n461, 
                           Y => n465);
   U634 : INVX1 port map( A => n466, Y => n1295);
   U635 : MUX2X1 port map( B => memory_31_2_port, A => RCV_DATA(2), S => n461, 
                           Y => n466);
   U636 : INVX1 port map( A => n467, Y => n1296);
   U637 : MUX2X1 port map( B => memory_31_1_port, A => RCV_DATA(1), S => n461, 
                           Y => n467);
   U638 : INVX1 port map( A => n468, Y => n1297);
   U639 : MUX2X1 port map( B => memory_31_0_port, A => RCV_DATA(0), S => n461, 
                           Y => n468);
   U640 : MUX2X1 port map( B => n469, A => n87, S => n470, Y => n1298);
   U641 : MUX2X1 port map( B => n471, A => n88, S => n470, Y => n1299);
   U642 : OAI21X1 port map( A => n193_port, B => n157, C => n21, Y => n470);
   U643 : MUX2X1 port map( B => n472, A => n87, S => n473, Y => n1300);
   U644 : MUX2X1 port map( B => n474, A => n88, S => n473, Y => n1301);
   U645 : OAI21X1 port map( A => n184, B => n157, C => n16, Y => n473);
   U646 : MUX2X1 port map( B => n475, A => n87, S => n476, Y => n1302);
   U647 : MUX2X1 port map( B => n477, A => n88, S => n476, Y => n1303);
   U648 : OAI21X1 port map( A => n244, B => n157, C => n19, Y => n476);
   U649 : NAND2X1 port map( A => n478, B => n2, Y => n157);
   U650 : MUX2X1 port map( B => n86, A => n479, S => n480, Y => n1304);
   U651 : MUX2X1 port map( B => n88, A => n481, S => n480, Y => n1305);
   U652 : NAND3X1 port map( A => n478, B => n361, C => n482, Y => n480);
   U653 : MUX2X1 port map( B => n184, A => n235, S => n483, Y => n482);
   U654 : AND2X1 port map( A => n360, B => n83, Y => n478);
   U655 : MUX2X1 port map( B => n86, A => n484, S => n485, Y => n1306);
   U656 : MUX2X1 port map( B => n88, A => n486, S => n485, Y => n1307);
   U657 : AOI21X1 port map( A => n123, B => n139, C => n69, Y => n485);
   U658 : INVX1 port map( A => n193_port, Y => n123);
   U659 : MUX2X1 port map( B => n86, A => n487, S => n488, Y => n1308);
   U660 : MUX2X1 port map( B => n88, A => n489, S => n488, Y => n1309);
   U661 : AOI21X1 port map( A => n118, B => n139, C => n70, Y => n488);
   U662 : INVX1 port map( A => n184, Y => n118);
   U663 : MUX2X1 port map( B => n86, A => n490, S => n491, Y => n1310);
   U664 : MUX2X1 port map( B => n88, A => n492, S => n491, Y => n1311);
   U665 : AOI21X1 port map( A => n113, B => n139, C => n71, Y => n491);
   U666 : NAND3X1 port map( A => n80, B => n75, C => n79, Y => n193_port);
   U667 : INVX1 port map( A => n244, Y => n113);
   U668 : MUX2X1 port map( B => n86, A => n493, S => n494, Y => n1312);
   U669 : MUX2X1 port map( B => n88, A => n495, S => n494, Y => n1313);
   U670 : AOI21X1 port map( A => n108, B => n139, C => n72, Y => n494);
   U671 : NAND3X1 port map( A => n81, B => n75, C => n79, Y => n184);
   U672 : NAND3X1 port map( A => n496, B => n82, C => n2, Y => n148);
   U673 : INVX1 port map( A => n235, Y => n108);
   U674 : MUX2X1 port map( B => n86, A => n497, S => n498, Y => n1314);
   U675 : INVX1 port map( A => opcode_28_1_port, Y => n497);
   U676 : MUX2X1 port map( B => n88, A => n499, S => n498, Y => n1315);
   U677 : AOI21X1 port map( A => n109, B => n143, C => n435, Y => n498);
   U678 : NAND3X1 port map( A => n80, B => n366, C => n76, Y => n244);
   U679 : INVX1 port map( A => n161, Y => n143);
   U680 : INVX1 port map( A => opcode_28_0_port, Y => n499);
   U681 : MUX2X1 port map( B => n86, A => n500, S => n501, Y => n1316);
   U682 : INVX1 port map( A => opcode_29_1_port, Y => n500);
   U683 : MUX2X1 port map( B => n88, A => n502, S => n501, Y => n1317);
   U684 : AOI21X1 port map( A => n109, B => n138, C => n73, Y => n501);
   U685 : NAND3X1 port map( A => n81, B => n366, C => n76, Y => n235);
   U686 : INVX1 port map( A => n156, Y => n138);
   U687 : NAND3X1 port map( A => n2, B => n496, C => n83, Y => n503);
   U688 : INVX1 port map( A => opcode_29_0_port, Y => n502);
   U689 : MUX2X1 port map( B => n86, A => n504, S => n505, Y => n1318);
   U690 : INVX1 port map( A => opcode_30_1_port, Y => n504);
   U691 : MUX2X1 port map( B => n88, A => n506, S => n505, Y => n1319);
   U692 : AOI21X1 port map( A => n133, B => n165, C => n74, Y => n505);
   U693 : NOR2X1 port map( A => n161, B => n43_port, Y => n452);
   U694 : NAND3X1 port map( A => n76, B => n80, C => n79, Y => n161);
   U695 : INVX1 port map( A => n152, Y => n133);
   U696 : NAND3X1 port map( A => n366, B => n75, C => n80, Y => n152);
   U697 : INVX1 port map( A => opcode_30_0_port, Y => n506);
   U698 : MUX2X1 port map( B => n87, A => n507, S => n508, Y => n1320);
   U699 : INVX1 port map( A => opcode_31_1_port, Y => n507);
   U700 : MUX2X1 port map( B => n106, A => n509, S => n508, Y => n1321);
   U701 : AOI21X1 port map( A => n128, B => n165, C => n461, Y => n508);
   U702 : NOR2X1 port map( A => n362, B => RST, Y => n496);
   U703 : INVX1 port map( A => writeptr_4_port, Y => n362);
   U704 : NAND3X1 port map( A => n76, B => n81, C => n79, Y => n156);
   U705 : NAND3X1 port map( A => n2, B => n82, C => n360, Y => n511);
   U706 : NOR2X1 port map( A => writeptr_4_port, B => RST, Y => n360);
   U707 : NAND2X1 port map( A => W_ENABLE, B => n311, Y => n510);
   U708 : NAND3X1 port map( A => n512, B => n513, C => n514, Y => n311);
   U709 : NOR2X1 port map( A => n515, B => n516, Y => n514);
   U710 : XOR2X1 port map( A => readptr_3_port, B => N34, Y => n515);
   U711 : XOR2X1 port map( A => n517, B => N32, Y => n513);
   U712 : NOR2X1 port map( A => n518, B => n519, Y => n512);
   U713 : XOR2X1 port map( A => readptr_2_port, B => N33, Y => n518);
   U714 : INVX1 port map( A => n147, Y => n128);
   U715 : NAND3X1 port map( A => n366, B => n75, C => n81, Y => n147);
   U716 : INVX1 port map( A => n79, Y => n366);
   U717 : INVX1 port map( A => opcode_31_0_port, Y => n509);
   U718 : INVX1 port map( A => n520, Y => n1322);
   U719 : MUX2X1 port map( B => n521, A => DATA_7_port, S => n522, Y => n520);
   U720 : NAND2X1 port map( A => n523, B => n524, Y => n521);
   U721 : NOR2X1 port map( A => n525, B => n526, Y => n524);
   U722 : NAND3X1 port map( A => n527, B => n528, C => n529, Y => n526);
   U723 : NOR2X1 port map( A => n530, B => n531, Y => n529);
   U724 : OAI22X1 port map( A => n402, B => n532, C => n410, D => n533, Y => 
                           n531);
   U725 : INVX1 port map( A => memory_17_7_port, Y => n410);
   U726 : INVX1 port map( A => memory_16_7_port, Y => n402);
   U727 : OAI22X1 port map( A => n418, B => n534, C => n426, D => n535, Y => 
                           n530);
   U728 : INVX1 port map( A => memory_19_7_port, Y => n426);
   U729 : INVX1 port map( A => memory_18_7_port, Y => n418);
   U730 : AOI22X1 port map( A => n536, B => memory_23_7_port, C => n537, D => 
                           memory_22_7_port, Y => n528);
   U731 : AOI22X1 port map( A => n538, B => memory_21_7_port, C => n539, D => 
                           memory_20_7_port, Y => n527);
   U732 : NAND3X1 port map( A => n540, B => n541, C => n542, Y => n525);
   U733 : NOR2X1 port map( A => n543, B => n544, Y => n542);
   U734 : OAI22X1 port map( A => n202, B => n545, C => n194, D => n546, Y => 
                           n544);
   U735 : INVX1 port map( A => memory_25_7_port, Y => n194);
   U736 : INVX1 port map( A => memory_24_7_port, Y => n202);
   U737 : OAI22X1 port map( A => n185, B => n547, C => n175, D => n548, Y => 
                           n543);
   U738 : INVX1 port map( A => memory_27_7_port, Y => n175);
   U739 : INVX1 port map( A => memory_26_7_port, Y => n185);
   U740 : AOI22X1 port map( A => n549, B => memory_31_7_port, C => n550, D => 
                           memory_30_7_port, Y => n541);
   U741 : AOI22X1 port map( A => n551, B => memory_29_7_port, C => n552, D => 
                           memory_28_7_port, Y => n540);
   U742 : NOR2X1 port map( A => n553, B => n554, Y => n523);
   U743 : NAND3X1 port map( A => n555, B => n556, C => n557, Y => n554);
   U744 : NOR2X1 port map( A => n558, B => n559, Y => n557);
   U745 : OAI22X1 port map( A => n310, B => n560, C => n302, D => n561, Y => 
                           n559);
   U746 : INVX1 port map( A => memory_2_7_port, Y => n302);
   U747 : INVX1 port map( A => memory_3_7_port, Y => n310);
   U748 : OAI22X1 port map( A => n294, B => n562, C => n285, D => n563, Y => 
                           n558);
   U749 : INVX1 port map( A => memory_0_7_port, Y => n285);
   U750 : INVX1 port map( A => memory_1_7_port, Y => n294);
   U751 : AOI22X1 port map( A => n564, B => memory_4_7_port, C => n565, D => 
                           memory_5_7_port, Y => n556);
   U752 : AOI22X1 port map( A => n566, B => memory_6_7_port, C => n567, D => 
                           memory_7_7_port, Y => n555);
   U753 : NAND3X1 port map( A => n568, B => n569, C => n570, Y => n553);
   U754 : NOR2X1 port map( A => n571, B => n572, Y => n570);
   U755 : OAI22X1 port map( A => n369, B => n573, C => n377, D => n574, Y => 
                           n572);
   U756 : INVX1 port map( A => memory_9_7_port, Y => n377);
   U757 : INVX1 port map( A => memory_8_7_port, Y => n369);
   U758 : OAI22X1 port map( A => n385, B => n575, C => n393, D => n576, Y => 
                           n571);
   U759 : INVX1 port map( A => memory_11_7_port, Y => n393);
   U760 : INVX1 port map( A => memory_10_7_port, Y => n385);
   U761 : AOI22X1 port map( A => n577, B => memory_15_7_port, C => n578, D => 
                           memory_14_7_port, Y => n569);
   U762 : AOI22X1 port map( A => n579, B => memory_13_7_port, C => n580, D => 
                           memory_12_7_port, Y => n568);
   U763 : INVX1 port map( A => n581, Y => n1323);
   U764 : MUX2X1 port map( B => n582, A => DATA_6_port, S => n522, Y => n581);
   U765 : NAND2X1 port map( A => n583, B => n584, Y => n582);
   U766 : NOR2X1 port map( A => n585, B => n586, Y => n584);
   U767 : NAND3X1 port map( A => n587, B => n588, C => n589, Y => n586);
   U768 : NOR2X1 port map( A => n590, B => n591, Y => n589);
   U769 : OAI22X1 port map( A => n403, B => n532, C => n411, D => n533, Y => 
                           n591);
   U770 : INVX1 port map( A => memory_17_6_port, Y => n411);
   U771 : INVX1 port map( A => memory_16_6_port, Y => n403);
   U772 : OAI22X1 port map( A => n419, B => n534, C => n427, D => n535, Y => 
                           n590);
   U773 : INVX1 port map( A => memory_19_6_port, Y => n427);
   U774 : INVX1 port map( A => memory_18_6_port, Y => n419);
   U775 : AOI22X1 port map( A => n536, B => memory_23_6_port, C => n537, D => 
                           memory_22_6_port, Y => n588);
   U776 : AOI22X1 port map( A => n538, B => memory_21_6_port, C => n539, D => 
                           memory_20_6_port, Y => n587);
   U777 : NAND3X1 port map( A => n592, B => n593, C => n594, Y => n585);
   U778 : NOR2X1 port map( A => n595, B => n596, Y => n594);
   U779 : OAI22X1 port map( A => n203, B => n545, C => n195_port, D => n546, Y 
                           => n596);
   U780 : INVX1 port map( A => memory_25_6_port, Y => n195_port);
   U781 : INVX1 port map( A => memory_24_6_port, Y => n203);
   U782 : OAI22X1 port map( A => n186, B => n547, C => n176, D => n548, Y => 
                           n595);
   U783 : INVX1 port map( A => memory_27_6_port, Y => n176);
   U784 : INVX1 port map( A => memory_26_6_port, Y => n186);
   U785 : AOI22X1 port map( A => n549, B => memory_31_6_port, C => n550, D => 
                           memory_30_6_port, Y => n593);
   U786 : AOI22X1 port map( A => n551, B => memory_29_6_port, C => n552, D => 
                           memory_28_6_port, Y => n592);
   U787 : NOR2X1 port map( A => n597, B => n598, Y => n583);
   U788 : NAND3X1 port map( A => n599, B => n600, C => n601, Y => n598);
   U789 : NOR2X1 port map( A => n602, B => n603, Y => n601);
   U790 : OAI22X1 port map( A => n309, B => n560, C => n301, D => n561, Y => 
                           n603);
   U791 : INVX1 port map( A => memory_2_6_port, Y => n301);
   U792 : INVX1 port map( A => memory_3_6_port, Y => n309);
   U793 : OAI22X1 port map( A => n293, B => n562, C => n284, D => n563, Y => 
                           n602);
   U794 : INVX1 port map( A => memory_0_6_port, Y => n284);
   U795 : INVX1 port map( A => memory_1_6_port, Y => n293);
   U796 : AOI22X1 port map( A => n564, B => memory_4_6_port, C => n565, D => 
                           memory_5_6_port, Y => n600);
   U797 : AOI22X1 port map( A => n566, B => memory_6_6_port, C => n567, D => 
                           memory_7_6_port, Y => n599);
   U798 : NAND3X1 port map( A => n604, B => n605, C => n606, Y => n597);
   U799 : NOR2X1 port map( A => n607, B => n608, Y => n606);
   U800 : OAI22X1 port map( A => n370, B => n573, C => n378, D => n574, Y => 
                           n608);
   U801 : INVX1 port map( A => memory_9_6_port, Y => n378);
   U802 : INVX1 port map( A => memory_8_6_port, Y => n370);
   U803 : OAI22X1 port map( A => n386, B => n575, C => n395, D => n576, Y => 
                           n607);
   U804 : INVX1 port map( A => memory_11_6_port, Y => n395);
   U805 : INVX1 port map( A => memory_10_6_port, Y => n386);
   U806 : AOI22X1 port map( A => n577, B => memory_15_6_port, C => n578, D => 
                           memory_14_6_port, Y => n605);
   U807 : AOI22X1 port map( A => n579, B => memory_13_6_port, C => n580, D => 
                           memory_12_6_port, Y => n604);
   U808 : INVX1 port map( A => n609, Y => n1324);
   U809 : MUX2X1 port map( B => n610, A => DATA_5_port, S => n522, Y => n609);
   U810 : NAND2X1 port map( A => n611, B => n612, Y => n610);
   U811 : NOR2X1 port map( A => n613, B => n614, Y => n612);
   U812 : NAND3X1 port map( A => n615, B => n616, C => n617, Y => n614);
   U813 : NOR2X1 port map( A => n618, B => n619, Y => n617);
   U814 : OAI22X1 port map( A => n404, B => n532, C => n412, D => n533, Y => 
                           n619);
   U815 : INVX1 port map( A => memory_17_5_port, Y => n412);
   U816 : INVX1 port map( A => memory_16_5_port, Y => n404);
   U817 : OAI22X1 port map( A => n420, B => n534, C => n428, D => n535, Y => 
                           n618);
   U818 : INVX1 port map( A => memory_19_5_port, Y => n428);
   U819 : INVX1 port map( A => memory_18_5_port, Y => n420);
   U820 : AOI22X1 port map( A => n536, B => memory_23_5_port, C => n537, D => 
                           memory_22_5_port, Y => n616);
   U821 : AOI22X1 port map( A => n538, B => memory_21_5_port, C => n539, D => 
                           memory_20_5_port, Y => n615);
   U822 : NAND3X1 port map( A => n620, B => n621, C => n622, Y => n613);
   U823 : NOR2X1 port map( A => n623, B => n624, Y => n622);
   U824 : OAI22X1 port map( A => n204, B => n545, C => n196, D => n546, Y => 
                           n624);
   U825 : INVX1 port map( A => memory_25_5_port, Y => n196);
   U826 : INVX1 port map( A => memory_24_5_port, Y => n204);
   U827 : OAI22X1 port map( A => n187, B => n547, C => n177, D => n548, Y => 
                           n623);
   U828 : INVX1 port map( A => memory_27_5_port, Y => n177);
   U829 : INVX1 port map( A => memory_26_5_port, Y => n187);
   U830 : AOI22X1 port map( A => n549, B => memory_31_5_port, C => n550, D => 
                           memory_30_5_port, Y => n621);
   U831 : AOI22X1 port map( A => n551, B => memory_29_5_port, C => n552, D => 
                           memory_28_5_port, Y => n620);
   U832 : NOR2X1 port map( A => n625, B => n626, Y => n611);
   U833 : NAND3X1 port map( A => n627, B => n628, C => n629, Y => n626);
   U834 : NOR2X1 port map( A => n630, B => n631, Y => n629);
   U835 : OAI22X1 port map( A => n308, B => n560, C => n300, D => n561, Y => 
                           n631);
   U836 : INVX1 port map( A => memory_2_5_port, Y => n300);
   U837 : INVX1 port map( A => memory_3_5_port, Y => n308);
   U838 : OAI22X1 port map( A => n292, B => n562, C => n283, D => n563, Y => 
                           n630);
   U839 : INVX1 port map( A => memory_0_5_port, Y => n283);
   U840 : INVX1 port map( A => memory_1_5_port, Y => n292);
   U841 : AOI22X1 port map( A => n564, B => memory_4_5_port, C => n565, D => 
                           memory_5_5_port, Y => n628);
   U842 : AOI22X1 port map( A => n566, B => memory_6_5_port, C => n567, D => 
                           memory_7_5_port, Y => n627);
   U843 : NAND3X1 port map( A => n632, B => n633, C => n634, Y => n625);
   U844 : NOR2X1 port map( A => n635, B => n636, Y => n634);
   U845 : OAI22X1 port map( A => n371, B => n573, C => n379, D => n574, Y => 
                           n636);
   U846 : INVX1 port map( A => memory_9_5_port, Y => n379);
   U847 : INVX1 port map( A => memory_8_5_port, Y => n371);
   U848 : OAI22X1 port map( A => n387, B => n575, C => n396, D => n576, Y => 
                           n635);
   U849 : INVX1 port map( A => memory_11_5_port, Y => n396);
   U850 : INVX1 port map( A => memory_10_5_port, Y => n387);
   U851 : AOI22X1 port map( A => n577, B => memory_15_5_port, C => n578, D => 
                           memory_14_5_port, Y => n633);
   U852 : AOI22X1 port map( A => n579, B => memory_13_5_port, C => n580, D => 
                           memory_12_5_port, Y => n632);
   U853 : INVX1 port map( A => n637, Y => n1325);
   U854 : MUX2X1 port map( B => n638, A => DATA_4_port, S => n522, Y => n637);
   U855 : NAND2X1 port map( A => n639, B => n640, Y => n638);
   U856 : NOR2X1 port map( A => n641, B => n642, Y => n640);
   U857 : NAND3X1 port map( A => n643, B => n644, C => n645, Y => n642);
   U858 : NOR2X1 port map( A => n646, B => n647, Y => n645);
   U859 : OAI22X1 port map( A => n405, B => n532, C => n413, D => n533, Y => 
                           n647);
   U860 : INVX1 port map( A => memory_17_4_port, Y => n413);
   U861 : INVX1 port map( A => memory_16_4_port, Y => n405);
   U862 : OAI22X1 port map( A => n421, B => n534, C => n429, D => n535, Y => 
                           n646);
   U863 : INVX1 port map( A => memory_19_4_port, Y => n429);
   U864 : INVX1 port map( A => memory_18_4_port, Y => n421);
   U865 : AOI22X1 port map( A => n536, B => memory_23_4_port, C => n537, D => 
                           memory_22_4_port, Y => n644);
   U866 : AOI22X1 port map( A => n538, B => memory_21_4_port, C => n539, D => 
                           memory_20_4_port, Y => n643);
   U867 : NAND3X1 port map( A => n648, B => n649, C => n650, Y => n641);
   U868 : NOR2X1 port map( A => n651, B => n652, Y => n650);
   U869 : OAI22X1 port map( A => n205, B => n545, C => n197, D => n546, Y => 
                           n652);
   U870 : INVX1 port map( A => memory_25_4_port, Y => n197);
   U871 : INVX1 port map( A => memory_24_4_port, Y => n205);
   U872 : OAI22X1 port map( A => n188, B => n547, C => n178, D => n548, Y => 
                           n651);
   U873 : INVX1 port map( A => memory_27_4_port, Y => n178);
   U874 : INVX1 port map( A => memory_26_4_port, Y => n188);
   U875 : AOI22X1 port map( A => n549, B => memory_31_4_port, C => n550, D => 
                           memory_30_4_port, Y => n649);
   U876 : AOI22X1 port map( A => n551, B => memory_29_4_port, C => n552, D => 
                           memory_28_4_port, Y => n648);
   U877 : NOR2X1 port map( A => n653, B => n654, Y => n639);
   U878 : NAND3X1 port map( A => n655, B => n656, C => n657, Y => n654);
   U879 : NOR2X1 port map( A => n658, B => n659, Y => n657);
   U880 : OAI22X1 port map( A => n307, B => n560, C => n299, D => n561, Y => 
                           n659);
   U881 : INVX1 port map( A => memory_2_4_port, Y => n299);
   U882 : INVX1 port map( A => memory_3_4_port, Y => n307);
   U883 : OAI22X1 port map( A => n291, B => n562, C => n282, D => n563, Y => 
                           n658);
   U884 : INVX1 port map( A => memory_0_4_port, Y => n282);
   U885 : INVX1 port map( A => memory_1_4_port, Y => n291);
   U886 : AOI22X1 port map( A => n564, B => memory_4_4_port, C => n565, D => 
                           memory_5_4_port, Y => n656);
   U887 : AOI22X1 port map( A => n566, B => memory_6_4_port, C => n567, D => 
                           memory_7_4_port, Y => n655);
   U888 : NAND3X1 port map( A => n660, B => n661, C => n662, Y => n653);
   U889 : NOR2X1 port map( A => n663, B => n664, Y => n662);
   U890 : OAI22X1 port map( A => n372, B => n573, C => n380, D => n574, Y => 
                           n664);
   U891 : INVX1 port map( A => memory_9_4_port, Y => n380);
   U892 : INVX1 port map( A => memory_8_4_port, Y => n372);
   U893 : OAI22X1 port map( A => n388, B => n575, C => n397, D => n576, Y => 
                           n663);
   U894 : INVX1 port map( A => memory_11_4_port, Y => n397);
   U895 : INVX1 port map( A => memory_10_4_port, Y => n388);
   U896 : AOI22X1 port map( A => n577, B => memory_15_4_port, C => n578, D => 
                           memory_14_4_port, Y => n661);
   U897 : AOI22X1 port map( A => n579, B => memory_13_4_port, C => n580, D => 
                           memory_12_4_port, Y => n660);
   U898 : INVX1 port map( A => n665, Y => n1326);
   U899 : MUX2X1 port map( B => n666, A => DATA_3_port, S => n522, Y => n665);
   U900 : NAND2X1 port map( A => n667, B => n668, Y => n666);
   U901 : NOR2X1 port map( A => n669, B => n670, Y => n668);
   U902 : NAND3X1 port map( A => n671, B => n672, C => n673, Y => n670);
   U903 : NOR2X1 port map( A => n674, B => n675, Y => n673);
   U904 : OAI22X1 port map( A => n406, B => n532, C => n414, D => n533, Y => 
                           n675);
   U905 : INVX1 port map( A => memory_17_3_port, Y => n414);
   U906 : INVX1 port map( A => memory_16_3_port, Y => n406);
   U907 : OAI22X1 port map( A => n422, B => n534, C => n430, D => n535, Y => 
                           n674);
   U908 : INVX1 port map( A => memory_19_3_port, Y => n430);
   U909 : INVX1 port map( A => memory_18_3_port, Y => n422);
   U910 : AOI22X1 port map( A => n536, B => memory_23_3_port, C => n537, D => 
                           memory_22_3_port, Y => n672);
   U911 : AOI22X1 port map( A => n538, B => memory_21_3_port, C => n539, D => 
                           memory_20_3_port, Y => n671);
   U912 : NAND3X1 port map( A => n676, B => n677, C => n678, Y => n669);
   U913 : NOR2X1 port map( A => n679, B => n680, Y => n678);
   U914 : OAI22X1 port map( A => n206, B => n545, C => n198, D => n546, Y => 
                           n680);
   U915 : INVX1 port map( A => memory_25_3_port, Y => n198);
   U916 : INVX1 port map( A => memory_24_3_port, Y => n206);
   U917 : OAI22X1 port map( A => n189_port, B => n547, C => n179, D => n548, Y 
                           => n679);
   U918 : INVX1 port map( A => memory_27_3_port, Y => n179);
   U919 : INVX1 port map( A => memory_26_3_port, Y => n189_port);
   U920 : AOI22X1 port map( A => n549, B => memory_31_3_port, C => n550, D => 
                           memory_30_3_port, Y => n677);
   U921 : AOI22X1 port map( A => n551, B => memory_29_3_port, C => n552, D => 
                           memory_28_3_port, Y => n676);
   U922 : NOR2X1 port map( A => n681, B => n682, Y => n667);
   U923 : NAND3X1 port map( A => n683, B => n684, C => n685, Y => n682);
   U924 : NOR2X1 port map( A => n686, B => n687, Y => n685);
   U925 : OAI22X1 port map( A => n306, B => n560, C => n298, D => n561, Y => 
                           n687);
   U926 : INVX1 port map( A => memory_2_3_port, Y => n298);
   U927 : INVX1 port map( A => memory_3_3_port, Y => n306);
   U928 : OAI22X1 port map( A => n290, B => n562, C => n281, D => n563, Y => 
                           n686);
   U929 : INVX1 port map( A => memory_0_3_port, Y => n281);
   U930 : INVX1 port map( A => memory_1_3_port, Y => n290);
   U931 : AOI22X1 port map( A => n564, B => memory_4_3_port, C => n565, D => 
                           memory_5_3_port, Y => n684);
   U932 : AOI22X1 port map( A => n566, B => memory_6_3_port, C => n567, D => 
                           memory_7_3_port, Y => n683);
   U933 : NAND3X1 port map( A => n688, B => n689, C => n690, Y => n681);
   U934 : NOR2X1 port map( A => n691, B => n692, Y => n690);
   U935 : OAI22X1 port map( A => n373, B => n573, C => n381, D => n574, Y => 
                           n692);
   U936 : INVX1 port map( A => memory_9_3_port, Y => n381);
   U937 : INVX1 port map( A => memory_8_3_port, Y => n373);
   U938 : OAI22X1 port map( A => n389, B => n575, C => n398, D => n576, Y => 
                           n691);
   U939 : INVX1 port map( A => memory_11_3_port, Y => n398);
   U940 : INVX1 port map( A => memory_10_3_port, Y => n389);
   U941 : AOI22X1 port map( A => n577, B => memory_15_3_port, C => n578, D => 
                           memory_14_3_port, Y => n689);
   U942 : AOI22X1 port map( A => n579, B => memory_13_3_port, C => n580, D => 
                           memory_12_3_port, Y => n688);
   U943 : INVX1 port map( A => n693, Y => n1327);
   U944 : MUX2X1 port map( B => n694, A => DATA_2_port, S => n522, Y => n693);
   U945 : NAND2X1 port map( A => n695, B => n696, Y => n694);
   U946 : NOR2X1 port map( A => n697, B => n698, Y => n696);
   U947 : NAND3X1 port map( A => n699, B => n700, C => n701, Y => n698);
   U948 : NOR2X1 port map( A => n702, B => n703, Y => n701);
   U949 : OAI22X1 port map( A => n407, B => n532, C => n415, D => n533, Y => 
                           n703);
   U950 : INVX1 port map( A => memory_17_2_port, Y => n415);
   U951 : INVX1 port map( A => memory_16_2_port, Y => n407);
   U952 : OAI22X1 port map( A => n423, B => n534, C => n431, D => n535, Y => 
                           n702);
   U953 : INVX1 port map( A => memory_19_2_port, Y => n431);
   U954 : INVX1 port map( A => memory_18_2_port, Y => n423);
   U955 : AOI22X1 port map( A => n536, B => memory_23_2_port, C => n537, D => 
                           memory_22_2_port, Y => n700);
   U956 : AOI22X1 port map( A => n538, B => memory_21_2_port, C => n539, D => 
                           memory_20_2_port, Y => n699);
   U957 : NAND3X1 port map( A => n704, B => n705, C => n706, Y => n697);
   U958 : NOR2X1 port map( A => n707, B => n708, Y => n706);
   U959 : OAI22X1 port map( A => n207, B => n545, C => n199, D => n546, Y => 
                           n708);
   U960 : INVX1 port map( A => memory_25_2_port, Y => n199);
   U961 : INVX1 port map( A => memory_24_2_port, Y => n207);
   U962 : OAI22X1 port map( A => n190_port, B => n547, C => n180, D => n548, Y 
                           => n707);
   U963 : INVX1 port map( A => memory_27_2_port, Y => n180);
   U964 : INVX1 port map( A => memory_26_2_port, Y => n190_port);
   U965 : AOI22X1 port map( A => n549, B => memory_31_2_port, C => n550, D => 
                           memory_30_2_port, Y => n705);
   U966 : AOI22X1 port map( A => n551, B => memory_29_2_port, C => n552, D => 
                           memory_28_2_port, Y => n704);
   U967 : NOR2X1 port map( A => n709, B => n710, Y => n695);
   U968 : NAND3X1 port map( A => n711, B => n712, C => n713, Y => n710);
   U969 : NOR2X1 port map( A => n714, B => n715, Y => n713);
   U970 : OAI22X1 port map( A => n305, B => n560, C => n297, D => n561, Y => 
                           n715);
   U971 : INVX1 port map( A => memory_2_2_port, Y => n297);
   U972 : INVX1 port map( A => memory_3_2_port, Y => n305);
   U973 : OAI22X1 port map( A => n289, B => n562, C => n280, D => n563, Y => 
                           n714);
   U974 : INVX1 port map( A => memory_0_2_port, Y => n280);
   U975 : INVX1 port map( A => memory_1_2_port, Y => n289);
   U976 : AOI22X1 port map( A => n564, B => memory_4_2_port, C => n565, D => 
                           memory_5_2_port, Y => n712);
   U977 : AOI22X1 port map( A => n566, B => memory_6_2_port, C => n567, D => 
                           memory_7_2_port, Y => n711);
   U978 : NAND3X1 port map( A => n716, B => n717, C => n718, Y => n709);
   U979 : NOR2X1 port map( A => n719, B => n720, Y => n718);
   U980 : OAI22X1 port map( A => n374, B => n573, C => n382, D => n574, Y => 
                           n720);
   U981 : INVX1 port map( A => memory_9_2_port, Y => n382);
   U982 : INVX1 port map( A => memory_8_2_port, Y => n374);
   U983 : OAI22X1 port map( A => n390, B => n575, C => n399, D => n576, Y => 
                           n719);
   U984 : INVX1 port map( A => memory_11_2_port, Y => n399);
   U985 : INVX1 port map( A => memory_10_2_port, Y => n390);
   U986 : AOI22X1 port map( A => n577, B => memory_15_2_port, C => n578, D => 
                           memory_14_2_port, Y => n717);
   U987 : AOI22X1 port map( A => n579, B => memory_13_2_port, C => n580, D => 
                           memory_12_2_port, Y => n716);
   U988 : INVX1 port map( A => n721, Y => n1328);
   U989 : MUX2X1 port map( B => n722, A => DATA_1_port, S => n522, Y => n721);
   U990 : NAND2X1 port map( A => n723, B => n724, Y => n722);
   U991 : NOR2X1 port map( A => n725, B => n726, Y => n724);
   U992 : NAND3X1 port map( A => n727, B => n728, C => n729, Y => n726);
   U993 : NOR2X1 port map( A => n730, B => n731, Y => n729);
   U994 : OAI22X1 port map( A => n408, B => n532, C => n416, D => n533, Y => 
                           n731);
   U995 : INVX1 port map( A => memory_17_1_port, Y => n416);
   U996 : INVX1 port map( A => memory_16_1_port, Y => n408);
   U997 : OAI22X1 port map( A => n424, B => n534, C => n432, D => n535, Y => 
                           n730);
   U998 : INVX1 port map( A => memory_19_1_port, Y => n432);
   U999 : INVX1 port map( A => memory_18_1_port, Y => n424);
   U1000 : AOI22X1 port map( A => n536, B => memory_23_1_port, C => n537, D => 
                           memory_22_1_port, Y => n728);
   U1001 : AOI22X1 port map( A => n538, B => memory_21_1_port, C => n539, D => 
                           memory_20_1_port, Y => n727);
   U1002 : NAND3X1 port map( A => n732, B => n733, C => n734, Y => n725);
   U1003 : NOR2X1 port map( A => n735, B => n736, Y => n734);
   U1004 : OAI22X1 port map( A => n208, B => n545, C => n200, D => n546, Y => 
                           n736);
   U1005 : INVX1 port map( A => memory_25_1_port, Y => n200);
   U1006 : INVX1 port map( A => memory_24_1_port, Y => n208);
   U1007 : OAI22X1 port map( A => n191_port, B => n547, C => n181, D => n548, Y
                           => n735);
   U1008 : INVX1 port map( A => memory_27_1_port, Y => n181);
   U1009 : INVX1 port map( A => memory_26_1_port, Y => n191_port);
   U1010 : AOI22X1 port map( A => n549, B => memory_31_1_port, C => n550, D => 
                           memory_30_1_port, Y => n733);
   U1011 : AOI22X1 port map( A => n551, B => memory_29_1_port, C => n552, D => 
                           memory_28_1_port, Y => n732);
   U1012 : NOR2X1 port map( A => n737, B => n738, Y => n723);
   U1013 : NAND3X1 port map( A => n739, B => n740, C => n741, Y => n738);
   U1014 : NOR2X1 port map( A => n742, B => n743, Y => n741);
   U1015 : OAI22X1 port map( A => n304, B => n560, C => n296, D => n561, Y => 
                           n743);
   U1016 : INVX1 port map( A => memory_2_1_port, Y => n296);
   U1017 : INVX1 port map( A => memory_3_1_port, Y => n304);
   U1018 : OAI22X1 port map( A => n288, B => n562, C => n279, D => n563, Y => 
                           n742);
   U1019 : INVX1 port map( A => memory_0_1_port, Y => n279);
   U1020 : INVX1 port map( A => memory_1_1_port, Y => n288);
   U1021 : AOI22X1 port map( A => n564, B => memory_4_1_port, C => n565, D => 
                           memory_5_1_port, Y => n740);
   U1022 : AOI22X1 port map( A => n566, B => memory_6_1_port, C => n567, D => 
                           memory_7_1_port, Y => n739);
   U1023 : NAND3X1 port map( A => n744, B => n745, C => n746, Y => n737);
   U1024 : NOR2X1 port map( A => n747, B => n748, Y => n746);
   U1025 : OAI22X1 port map( A => n375, B => n573, C => n383, D => n574, Y => 
                           n748);
   U1026 : INVX1 port map( A => memory_9_1_port, Y => n383);
   U1027 : INVX1 port map( A => memory_8_1_port, Y => n375);
   U1028 : OAI22X1 port map( A => n391, B => n575, C => n400, D => n576, Y => 
                           n747);
   U1029 : INVX1 port map( A => memory_11_1_port, Y => n400);
   U1030 : INVX1 port map( A => memory_10_1_port, Y => n391);
   U1031 : AOI22X1 port map( A => n577, B => memory_15_1_port, C => n578, D => 
                           memory_14_1_port, Y => n745);
   U1032 : AOI22X1 port map( A => n579, B => memory_13_1_port, C => n580, D => 
                           memory_12_1_port, Y => n744);
   U1033 : INVX1 port map( A => n749, Y => n1329);
   U1034 : MUX2X1 port map( B => n750, A => DATA_0_port, S => n522, Y => n749);
   U1035 : NAND2X1 port map( A => n751, B => n752, Y => n750);
   U1036 : NOR2X1 port map( A => n753, B => n754, Y => n752);
   U1037 : NAND3X1 port map( A => n755, B => n756, C => n757, Y => n754);
   U1038 : NOR2X1 port map( A => n758, B => n759, Y => n757);
   U1039 : OAI22X1 port map( A => n409, B => n532, C => n417, D => n533, Y => 
                           n759);
   U1040 : INVX1 port map( A => memory_17_0_port, Y => n417);
   U1041 : INVX1 port map( A => memory_16_0_port, Y => n409);
   U1042 : OAI22X1 port map( A => n425, B => n534, C => n433, D => n535, Y => 
                           n758);
   U1043 : INVX1 port map( A => memory_19_0_port, Y => n433);
   U1044 : INVX1 port map( A => memory_18_0_port, Y => n425);
   U1045 : AOI22X1 port map( A => n536, B => memory_23_0_port, C => n537, D => 
                           memory_22_0_port, Y => n756);
   U1046 : AOI22X1 port map( A => n538, B => memory_21_0_port, C => n539, D => 
                           memory_20_0_port, Y => n755);
   U1047 : NAND3X1 port map( A => n760, B => n761, C => n762, Y => n753);
   U1048 : NOR2X1 port map( A => n763, B => n764, Y => n762);
   U1049 : OAI22X1 port map( A => n209, B => n545, C => n201, D => n546, Y => 
                           n764);
   U1050 : INVX1 port map( A => memory_25_0_port, Y => n201);
   U1051 : INVX1 port map( A => memory_24_0_port, Y => n209);
   U1052 : OAI22X1 port map( A => n192_port, B => n547, C => n182, D => n548, Y
                           => n763);
   U1053 : INVX1 port map( A => memory_27_0_port, Y => n182);
   U1054 : INVX1 port map( A => memory_26_0_port, Y => n192_port);
   U1055 : AOI22X1 port map( A => n549, B => memory_31_0_port, C => n550, D => 
                           memory_30_0_port, Y => n761);
   U1056 : AOI22X1 port map( A => n551, B => memory_29_0_port, C => n552, D => 
                           memory_28_0_port, Y => n760);
   U1057 : NOR2X1 port map( A => n765, B => n766, Y => n751);
   U1058 : NAND3X1 port map( A => n767, B => n768, C => n769, Y => n766);
   U1059 : NOR2X1 port map( A => n770, B => n771, Y => n769);
   U1060 : OAI22X1 port map( A => n303, B => n560, C => n295, D => n561, Y => 
                           n771);
   U1061 : INVX1 port map( A => memory_2_0_port, Y => n295);
   U1062 : INVX1 port map( A => memory_3_0_port, Y => n303);
   U1063 : OAI22X1 port map( A => n287, B => n562, C => n278, D => n563, Y => 
                           n770);
   U1064 : INVX1 port map( A => memory_0_0_port, Y => n278);
   U1065 : INVX1 port map( A => memory_1_0_port, Y => n287);
   U1066 : AOI22X1 port map( A => n564, B => memory_4_0_port, C => n565, D => 
                           memory_5_0_port, Y => n768);
   U1067 : AOI22X1 port map( A => n566, B => memory_6_0_port, C => n567, D => 
                           memory_7_0_port, Y => n767);
   U1068 : NAND3X1 port map( A => n772, B => n773, C => n774, Y => n765);
   U1069 : NOR2X1 port map( A => n775, B => n776, Y => n774);
   U1070 : OAI22X1 port map( A => n376, B => n573, C => n384, D => n574, Y => 
                           n776);
   U1071 : INVX1 port map( A => memory_9_0_port, Y => n384);
   U1072 : INVX1 port map( A => memory_8_0_port, Y => n376);
   U1073 : OAI22X1 port map( A => n392, B => n575, C => n401, D => n576, Y => 
                           n775);
   U1074 : INVX1 port map( A => memory_11_0_port, Y => n401);
   U1075 : INVX1 port map( A => memory_10_0_port, Y => n392);
   U1076 : AOI22X1 port map( A => n577, B => memory_15_0_port, C => n578, D => 
                           memory_14_0_port, Y => n773);
   U1077 : AOI22X1 port map( A => n579, B => memory_13_0_port, C => n580, D => 
                           memory_12_0_port, Y => n772);
   U1078 : INVX1 port map( A => n777, Y => n1330);
   U1079 : MUX2X1 port map( B => n778, A => OUT_OPCODE_1_port, S => n522, Y => 
                           n777);
   U1080 : NAND2X1 port map( A => n779, B => n780, Y => n778);
   U1081 : NOR2X1 port map( A => n781, B => n782, Y => n780);
   U1082 : NAND3X1 port map( A => n783, B => n784, C => n785, Y => n782);
   U1083 : NOR2X1 port map( A => n786, B => n787, Y => n785);
   U1084 : OAI22X1 port map( A => n484, B => n532, C => n487, D => n533, Y => 
                           n787);
   U1085 : INVX1 port map( A => opcode_17_1_port, Y => n487);
   U1086 : INVX1 port map( A => opcode_16_1_port, Y => n484);
   U1087 : OAI22X1 port map( A => n490, B => n534, C => n493, D => n535, Y => 
                           n786);
   U1088 : INVX1 port map( A => opcode_19_1_port, Y => n493);
   U1089 : INVX1 port map( A => opcode_18_1_port, Y => n490);
   U1090 : AOI22X1 port map( A => n536, B => opcode_23_1_port, C => n537, D => 
                           opcode_22_1_port, Y => n784);
   U1091 : AOI22X1 port map( A => n538, B => opcode_21_1_port, C => n539, D => 
                           opcode_20_1_port, Y => n783);
   U1092 : NAND3X1 port map( A => n788, B => n789, C => n790, Y => n781);
   U1093 : NOR2X1 port map( A => n791, B => n792, Y => n790);
   U1094 : OAI22X1 port map( A => n120, B => n545, C => n115, D => n546, Y => 
                           n792);
   U1095 : INVX1 port map( A => opcode_25_1_port, Y => n115);
   U1096 : INVX1 port map( A => opcode_24_1_port, Y => n120);
   U1097 : OAI22X1 port map( A => n110, B => n547, C => n104, D => n548, Y => 
                           n791);
   U1098 : INVX1 port map( A => opcode_27_1_port, Y => n104);
   U1099 : INVX1 port map( A => opcode_26_1_port, Y => n110);
   U1100 : AOI22X1 port map( A => n549, B => opcode_31_1_port, C => n550, D => 
                           opcode_30_1_port, Y => n789);
   U1101 : AOI22X1 port map( A => n551, B => opcode_29_1_port, C => n552, D => 
                           opcode_28_1_port, Y => n788);
   U1102 : NOR2X1 port map( A => n793, B => n794, Y => n779);
   U1103 : NAND3X1 port map( A => n795, B => n796, C => n797, Y => n794);
   U1104 : NOR2X1 port map( A => n798, B => n799, Y => n797);
   U1105 : OAI22X1 port map( A => n174, B => n560, C => n171, D => n561, Y => 
                           n799);
   U1106 : INVX1 port map( A => opcode_2_1_port, Y => n171);
   U1107 : INVX1 port map( A => opcode_3_1_port, Y => n174);
   U1108 : OAI22X1 port map( A => n168, B => n562, C => n164, D => n563, Y => 
                           n798);
   U1109 : INVX1 port map( A => opcode_0_1_port, Y => n164);
   U1110 : INVX1 port map( A => opcode_1_1_port, Y => n168);
   U1111 : AOI22X1 port map( A => n564, B => opcode_4_1_port, C => n565, D => 
                           opcode_5_1_port, Y => n796);
   U1112 : AOI22X1 port map( A => n566, B => opcode_6_1_port, C => n567, D => 
                           opcode_7_1_port, Y => n795);
   U1113 : NAND3X1 port map( A => n800, B => n801, C => n802, Y => n793);
   U1114 : NOR2X1 port map( A => n803, B => n804, Y => n802);
   U1115 : OAI22X1 port map( A => n469, B => n573, C => n472, D => n574, Y => 
                           n804);
   U1116 : INVX1 port map( A => opcode_9_1_port, Y => n472);
   U1117 : INVX1 port map( A => opcode_8_1_port, Y => n469);
   U1118 : OAI22X1 port map( A => n475, B => n575, C => n479, D => n576, Y => 
                           n803);
   U1119 : INVX1 port map( A => opcode_11_1_port, Y => n479);
   U1120 : INVX1 port map( A => opcode_10_1_port, Y => n475);
   U1121 : AOI22X1 port map( A => n577, B => opcode_15_1_port, C => n578, D => 
                           opcode_14_1_port, Y => n801);
   U1122 : AOI22X1 port map( A => n579, B => opcode_13_1_port, C => n580, D => 
                           opcode_12_1_port, Y => n800);
   U1123 : INVX1 port map( A => n805, Y => n1331);
   U1124 : MUX2X1 port map( B => n806, A => OUT_OPCODE_0_port, S => n522, Y => 
                           n805);
   U1125 : NAND3X1 port map( A => N195, B => n98, C => n84, Y => n522);
   U1126 : NAND2X1 port map( A => n807, B => n808, Y => n806);
   U1127 : NOR2X1 port map( A => n809, B => n810, Y => n808);
   U1128 : NAND3X1 port map( A => n811, B => n812, C => n813, Y => n810);
   U1129 : NOR2X1 port map( A => n814, B => n815, Y => n813);
   U1130 : OAI22X1 port map( A => n486, B => n532, C => n489, D => n533, Y => 
                           n815);
   U1131 : NAND2X1 port map( A => n816, B => n817, Y => n533);
   U1132 : INVX1 port map( A => opcode_17_0_port, Y => n489);
   U1133 : NAND2X1 port map( A => n818, B => n817, Y => n532);
   U1134 : INVX1 port map( A => opcode_16_0_port, Y => n486);
   U1135 : OAI22X1 port map( A => n492, B => n534, C => n495, D => n535, Y => 
                           n814);
   U1136 : NAND2X1 port map( A => n816, B => n819, Y => n535);
   U1137 : INVX1 port map( A => opcode_19_0_port, Y => n495);
   U1138 : NAND2X1 port map( A => n818, B => n819, Y => n534);
   U1139 : INVX1 port map( A => opcode_18_0_port, Y => n492);
   U1140 : AOI22X1 port map( A => n536, B => opcode_23_0_port, C => n537, D => 
                           opcode_22_0_port, Y => n812);
   U1141 : AOI22X1 port map( A => n538, B => opcode_21_0_port, C => n539, D => 
                           opcode_20_0_port, Y => n811);
   U1142 : INVX1 port map( A => n822, Y => n818);
   U1143 : NAND3X1 port map( A => n823, B => n824, C => readptr_4_port, Y => 
                           n822);
   U1144 : INVX1 port map( A => n825, Y => n816);
   U1145 : NAND3X1 port map( A => readptr_0_port, B => n824, C => 
                           readptr_4_port, Y => n825);
   U1146 : NAND3X1 port map( A => n826, B => n827, C => n828, Y => n809);
   U1147 : NOR2X1 port map( A => n829, B => n830, Y => n828);
   U1148 : OAI22X1 port map( A => n122, B => n545, C => n117, D => n546, Y => 
                           n830);
   U1149 : NAND2X1 port map( A => n817, B => n831, Y => n546);
   U1150 : INVX1 port map( A => opcode_25_0_port, Y => n117);
   U1151 : NAND2X1 port map( A => n817, B => n832, Y => n545);
   U1152 : INVX1 port map( A => opcode_24_0_port, Y => n122);
   U1153 : OAI22X1 port map( A => n112, B => n547, C => n107, D => n548, Y => 
                           n829);
   U1154 : NAND2X1 port map( A => n819, B => n831, Y => n548);
   U1155 : INVX1 port map( A => opcode_27_0_port, Y => n107);
   U1156 : NAND2X1 port map( A => n819, B => n832, Y => n547);
   U1157 : INVX1 port map( A => opcode_26_0_port, Y => n112);
   U1158 : AOI22X1 port map( A => n549, B => opcode_31_0_port, C => n550, D => 
                           opcode_30_0_port, Y => n827);
   U1159 : AOI22X1 port map( A => n551, B => opcode_29_0_port, C => n552, D => 
                           opcode_28_0_port, Y => n826);
   U1160 : INVX1 port map( A => n833, Y => n832);
   U1161 : NAND3X1 port map( A => readptr_3_port, B => n823, C => 
                           readptr_4_port, Y => n833);
   U1162 : INVX1 port map( A => n834, Y => n831);
   U1163 : NAND3X1 port map( A => readptr_3_port, B => readptr_0_port, C => 
                           readptr_4_port, Y => n834);
   U1164 : NOR2X1 port map( A => n835, B => n836, Y => n807);
   U1165 : NAND3X1 port map( A => n837, B => n838, C => n839, Y => n836);
   U1166 : NOR2X1 port map( A => n840, B => n841, Y => n839);
   U1167 : OAI22X1 port map( A => n172, B => n560, C => n169, D => n561, Y => 
                           n841);
   U1168 : NAND2X1 port map( A => n842, B => n819, Y => n561);
   U1169 : INVX1 port map( A => opcode_2_0_port, Y => n169);
   U1170 : NAND2X1 port map( A => n843, B => n819, Y => n560);
   U1171 : INVX1 port map( A => opcode_3_0_port, Y => n172);
   U1172 : OAI22X1 port map( A => n166, B => n562, C => n162, D => n563, Y => 
                           n840);
   U1173 : NAND2X1 port map( A => n842, B => n817, Y => n563);
   U1174 : INVX1 port map( A => opcode_0_0_port, Y => n162);
   U1175 : NAND2X1 port map( A => n843, B => n817, Y => n562);
   U1176 : INVX1 port map( A => opcode_1_0_port, Y => n166);
   U1177 : AOI22X1 port map( A => n564, B => opcode_4_0_port, C => n565, D => 
                           opcode_5_0_port, Y => n838);
   U1178 : AOI22X1 port map( A => n566, B => opcode_6_0_port, C => n567, D => 
                           opcode_7_0_port, Y => n837);
   U1179 : INVX1 port map( A => n844, Y => n843);
   U1180 : NAND3X1 port map( A => n824, B => n845, C => readptr_0_port, Y => 
                           n844);
   U1181 : INVX1 port map( A => n846, Y => n842);
   U1182 : NAND3X1 port map( A => n824, B => n845, C => n823, Y => n846);
   U1183 : INVX1 port map( A => readptr_3_port, Y => n824);
   U1184 : NAND3X1 port map( A => n847, B => n848, C => n849, Y => n835);
   U1185 : NOR2X1 port map( A => n850, B => n851, Y => n849);
   U1186 : OAI22X1 port map( A => n471, B => n573, C => n474, D => n574, Y => 
                           n851);
   U1187 : NAND2X1 port map( A => n852, B => n817, Y => n574);
   U1188 : INVX1 port map( A => opcode_9_0_port, Y => n474);
   U1189 : NAND2X1 port map( A => n853, B => n817, Y => n573);
   U1190 : NOR2X1 port map( A => readptr_1_port, B => readptr_2_port, Y => n817
                           );
   U1191 : INVX1 port map( A => opcode_8_0_port, Y => n471);
   U1192 : OAI22X1 port map( A => n477, B => n575, C => n481, D => n576, Y => 
                           n850);
   U1193 : NAND2X1 port map( A => n852, B => n819, Y => n576);
   U1194 : INVX1 port map( A => opcode_11_0_port, Y => n481);
   U1195 : NAND2X1 port map( A => n853, B => n819, Y => n575);
   U1196 : NOR2X1 port map( A => n517, B => readptr_2_port, Y => n819);
   U1197 : INVX1 port map( A => opcode_10_0_port, Y => n477);
   U1198 : AOI22X1 port map( A => n577, B => opcode_15_0_port, C => n578, D => 
                           opcode_14_0_port, Y => n848);
   U1199 : NOR2X1 port map( A => n517, B => n855, Y => n820);
   U1200 : AOI22X1 port map( A => n579, B => opcode_13_0_port, C => n580, D => 
                           opcode_12_0_port, Y => n847);
   U1201 : INVX1 port map( A => n857, Y => n853);
   U1202 : NAND3X1 port map( A => n823, B => n845, C => readptr_3_port, Y => 
                           n857);
   U1203 : INVX1 port map( A => readptr_0_port, Y => n823);
   U1204 : NOR2X1 port map( A => n855, B => readptr_1_port, Y => n821);
   U1205 : INVX1 port map( A => readptr_2_port, Y => n855);
   U1207 : INVX1 port map( A => n859, Y => n852);
   U1208 : NAND3X1 port map( A => readptr_0_port, B => n845, C => 
                           readptr_3_port, Y => n859);
   U1209 : INVX1 port map( A => readptr_4_port, Y => n845);
   U1210 : AND2X1 port map( A => N337, B => n84, Y => N347);
   U1211 : AND2X1 port map( A => N336, B => n84, Y => N346);
   U1212 : AND2X1 port map( A => N335, B => n84, Y => N345);
   U1213 : AND2X1 port map( A => N334, B => n84, Y => N344);
   U1214 : AND2X1 port map( A => N333, B => n84, Y => N343);
   U1215 : AND2X1 port map( A => N193, B => n84, Y => N342);
   U1216 : AND2X1 port map( A => N192, B => n84, Y => N341);
   U1217 : AND2X1 port map( A => N191, B => n84, Y => N340);
   U1218 : AND2X1 port map( A => N190, B => n84, Y => N339);
   U1219 : AND2X1 port map( A => N189, B => n84, Y => N338);
   U1220 : AND2X1 port map( A => R_ENABLE, B => n313, Y => N195);
   U1221 : NAND3X1 port map( A => n861, B => n863, C => n864, Y => n313);
   U1222 : NOR2X1 port map( A => n865, B => n866, Y => n864);
   U1223 : XOR2X1 port map( A => writeptr_4_port, B => readptr_4_port, Y => 
                           n866);
   U1224 : XOR2X1 port map( A => n83, B => readptr_3_port, Y => n865);
   U1225 : XOR2X1 port map( A => n517, B => n78, Y => n863);
   U1226 : INVX1 port map( A => readptr_1_port, Y => n517);
   U1227 : NOR2X1 port map( A => n867, B => n909, Y => n861);
   U1228 : XOR2X1 port map( A => n81, B => readptr_0_port, Y => n909);
   U1229 : XOR2X1 port map( A => n76, B => readptr_2_port, Y => n867);

end SYN_BRFIFO;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RBUFFER_0 is

   port( CLK, RST, NEXT_BYTE : in std_logic;  DATA : in std_logic_vector (7 
         downto 0);  OPCODE : in std_logic_vector (1 downto 0);  BYTE_COUNT : 
         in std_logic_vector (4 downto 0);  EOP : in std_logic;  B_READY, 
         R_ENABLE : out std_logic;  PRGA_IN : out std_logic_vector (7 downto 0)
         ;  PRGA_OPCODE : out std_logic_vector (1 downto 0));

end RBUFFER_0;

architecture SYN_brbuffer of RBUFFER_0 is

   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal B_READY_port, R_ENABLE_port, PRGA_IN_7_port, PRGA_IN_6_port, 
      PRGA_IN_5_port, PRGA_IN_4_port, PRGA_IN_3_port, PRGA_IN_2_port, 
      PRGA_IN_1_port, PRGA_IN_0_port, PRGA_OPCODE_1_port, PRGA_OPCODE_0_port, 
      state_2_port, state_1_port, state_0_port, nextState_2_port, 
      nextState_1_port, nextState_0_port, tempData_7_port, tempData_6_port, 
      tempData_5_port, tempData_4_port, tempData_3_port, tempData_2_port, 
      tempData_1_port, tempData_0_port, tempOpcode_1_port, tempOpcode_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103 : std_logic;

begin
   B_READY <= B_READY_port;
   R_ENABLE <= R_ENABLE_port;
   PRGA_IN <= ( PRGA_IN_7_port, PRGA_IN_6_port, PRGA_IN_5_port, PRGA_IN_4_port,
      PRGA_IN_3_port, PRGA_IN_2_port, PRGA_IN_1_port, PRGA_IN_0_port );
   PRGA_OPCODE <= ( PRGA_OPCODE_1_port, PRGA_OPCODE_0_port );
   
   B_READY_reg : DFFPOSX1 port map( D => n92, CLK => CLK, Q => B_READY_port);
   tempData_reg_7_inst : DFFPOSX1 port map( D => n71, CLK => CLK, Q => 
                           tempData_7_port);
   tempData_reg_6_inst : DFFPOSX1 port map( D => n72, CLK => CLK, Q => 
                           tempData_6_port);
   tempData_reg_5_inst : DFFPOSX1 port map( D => n73, CLK => CLK, Q => 
                           tempData_5_port);
   tempData_reg_4_inst : DFFPOSX1 port map( D => n74, CLK => CLK, Q => 
                           tempData_4_port);
   tempData_reg_3_inst : DFFPOSX1 port map( D => n75, CLK => CLK, Q => 
                           tempData_3_port);
   tempData_reg_2_inst : DFFPOSX1 port map( D => n86, CLK => CLK, Q => 
                           tempData_2_port);
   tempData_reg_1_inst : DFFPOSX1 port map( D => n88, CLK => CLK, Q => 
                           tempData_1_port);
   tempData_reg_0_inst : DFFPOSX1 port map( D => n89, CLK => CLK, Q => 
                           tempData_0_port);
   tempOpcode_reg_1_inst : DFFPOSX1 port map( D => n90, CLK => CLK, Q => 
                           tempOpcode_1_port);
   PRGA_OPCODE_reg_1_inst : DFFPOSX1 port map( D => n93, CLK => CLK, Q => 
                           PRGA_OPCODE_1_port);
   tempOpcode_reg_0_inst : DFFPOSX1 port map( D => n91, CLK => CLK, Q => 
                           tempOpcode_0_port);
   PRGA_OPCODE_reg_0_inst : DFFPOSX1 port map( D => n94, CLK => CLK, Q => 
                           PRGA_OPCODE_0_port);
   R_ENABLE_reg : DFFPOSX1 port map( D => n95, CLK => CLK, Q => R_ENABLE_port);
   PRGA_IN_reg_7_inst : DFFPOSX1 port map( D => n96, CLK => CLK, Q => 
                           PRGA_IN_7_port);
   PRGA_IN_reg_6_inst : DFFPOSX1 port map( D => n97, CLK => CLK, Q => 
                           PRGA_IN_6_port);
   PRGA_IN_reg_5_inst : DFFPOSX1 port map( D => n98, CLK => CLK, Q => 
                           PRGA_IN_5_port);
   PRGA_IN_reg_4_inst : DFFPOSX1 port map( D => n99, CLK => CLK, Q => 
                           PRGA_IN_4_port);
   PRGA_IN_reg_3_inst : DFFPOSX1 port map( D => n100, CLK => CLK, Q => 
                           PRGA_IN_3_port);
   PRGA_IN_reg_2_inst : DFFPOSX1 port map( D => n101, CLK => CLK, Q => 
                           PRGA_IN_2_port);
   PRGA_IN_reg_1_inst : DFFPOSX1 port map( D => n102, CLK => CLK, Q => 
                           PRGA_IN_1_port);
   PRGA_IN_reg_0_inst : DFFPOSX1 port map( D => n103, CLK => CLK, Q => 
                           PRGA_IN_0_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n4, S => n3, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n4, S => n2, Q => state_2_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n4, S => n1, Q => state_0_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   U6 : INVX2 port map( A => n44, Y => n31);
   U7 : INVX2 port map( A => RST, Y => n4);
   U8 : OR2X2 port map( A => n42, B => RST, Y => n32);
   U9 : AND2X2 port map( A => n42, B => n4, Y => n47);
   U10 : OAI21X1 port map( A => n5, B => n6, C => n7, Y => nextState_2_port);
   U11 : MUX2X1 port map( B => n8, A => n9, S => state_0_port, Y => n7);
   U12 : NOR2X1 port map( A => state_2_port, B => n10, Y => n9);
   U13 : AND2X1 port map( A => state_2_port, B => n11, Y => n8);
   U14 : OAI21X1 port map( A => NEXT_BYTE, B => n12, C => state_1_port, Y => 
                           n11);
   U15 : AND2X1 port map( A => n13, B => NEXT_BYTE, Y => n5);
   U16 : OAI21X1 port map( A => state_2_port, B => n14, C => n15, Y => 
                           nextState_1_port);
   U17 : OAI21X1 port map( A => n16, B => n17, C => n18, Y => n15);
   U18 : INVX1 port map( A => n6, Y => n17);
   U19 : OAI21X1 port map( A => state_2_port, B => n19, C => n20, Y => 
                           nextState_0_port);
   U20 : AOI22X1 port map( A => n21, B => n22, C => NEXT_BYTE, D => n23, Y => 
                           n20);
   U21 : OAI21X1 port map( A => n13, B => n6, C => n24, Y => n23);
   U22 : INVX1 port map( A => n16, Y => n24);
   U23 : NOR2X1 port map( A => n19, B => n12, Y => n16);
   U24 : NOR2X1 port map( A => n25, B => BYTE_COUNT(4), Y => n12);
   U25 : NAND3X1 port map( A => state_0_port, B => n10, C => state_2_port, Y =>
                           n6);
   U26 : AND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n13);
   U27 : OAI21X1 port map( A => n26, B => n18, C => n27, Y => n22);
   U28 : INVX1 port map( A => NEXT_BYTE, Y => n18);
   U29 : AOI21X1 port map( A => EOP, B => n25, C => BYTE_COUNT(4), Y => n26);
   U30 : NAND2X1 port map( A => n28, B => n29, Y => n25);
   U31 : NOR2X1 port map( A => BYTE_COUNT(3), B => BYTE_COUNT(2), Y => n29);
   U32 : NOR2X1 port map( A => BYTE_COUNT(1), B => BYTE_COUNT(0), Y => n28);
   U33 : NOR2X1 port map( A => state_1_port, B => state_0_port, Y => n21);
   U34 : INVX1 port map( A => n30, Y => n71);
   U35 : AOI22X1 port map( A => n31, B => DATA(7), C => n32, D => 
                           tempData_7_port, Y => n30);
   U36 : INVX1 port map( A => n33, Y => n72);
   U37 : AOI22X1 port map( A => n31, B => DATA(6), C => n32, D => 
                           tempData_6_port, Y => n33);
   U38 : INVX1 port map( A => n34, Y => n73);
   U39 : AOI22X1 port map( A => n31, B => DATA(5), C => n32, D => 
                           tempData_5_port, Y => n34);
   U40 : INVX1 port map( A => n35, Y => n74);
   U41 : AOI22X1 port map( A => n31, B => DATA(4), C => n32, D => 
                           tempData_4_port, Y => n35);
   U42 : INVX1 port map( A => n36, Y => n75);
   U43 : AOI22X1 port map( A => n31, B => DATA(3), C => n32, D => 
                           tempData_3_port, Y => n36);
   U44 : INVX1 port map( A => n37, Y => n86);
   U45 : AOI22X1 port map( A => n31, B => DATA(2), C => n32, D => 
                           tempData_2_port, Y => n37);
   U46 : INVX1 port map( A => n38, Y => n88);
   U47 : AOI22X1 port map( A => n31, B => DATA(1), C => n32, D => 
                           tempData_1_port, Y => n38);
   U48 : INVX1 port map( A => n39, Y => n89);
   U49 : AOI22X1 port map( A => n31, B => DATA(0), C => n32, D => 
                           tempData_0_port, Y => n39);
   U50 : INVX1 port map( A => n40, Y => n90);
   U51 : AOI22X1 port map( A => OPCODE(1), B => n31, C => n32, D => 
                           tempOpcode_1_port, Y => n40);
   U52 : INVX1 port map( A => n41, Y => n91);
   U53 : AOI22X1 port map( A => OPCODE(0), B => n31, C => n32, D => 
                           tempOpcode_0_port, Y => n41);
   U54 : OAI21X1 port map( A => n4, B => n43, C => n44, Y => n92);
   U55 : INVX1 port map( A => B_READY_port, Y => n43);
   U56 : OAI21X1 port map( A => n4, B => n45, C => n46, Y => n93);
   U57 : AOI22X1 port map( A => n31, B => OPCODE(1), C => n47, D => 
                           tempOpcode_1_port, Y => n46);
   U58 : INVX1 port map( A => PRGA_OPCODE_1_port, Y => n45);
   U59 : OAI21X1 port map( A => n4, B => n48, C => n49, Y => n94);
   U60 : AOI22X1 port map( A => n31, B => OPCODE(0), C => n47, D => 
                           tempOpcode_0_port, Y => n49);
   U61 : INVX1 port map( A => PRGA_OPCODE_0_port, Y => n48);
   U62 : MUX2X1 port map( B => n50, A => n51, S => RST, Y => n95);
   U63 : INVX1 port map( A => R_ENABLE_port, Y => n51);
   U64 : NAND3X1 port map( A => n10, B => n27, C => state_0_port, Y => n50);
   U65 : OAI21X1 port map( A => n4, B => n52, C => n53, Y => n96);
   U66 : AOI22X1 port map( A => DATA(7), B => n31, C => n47, D => 
                           tempData_7_port, Y => n53);
   U67 : INVX1 port map( A => PRGA_IN_7_port, Y => n52);
   U68 : OAI21X1 port map( A => n4, B => n54, C => n55, Y => n97);
   U69 : AOI22X1 port map( A => DATA(6), B => n31, C => n47, D => 
                           tempData_6_port, Y => n55);
   U70 : INVX1 port map( A => PRGA_IN_6_port, Y => n54);
   U71 : OAI21X1 port map( A => n4, B => n56, C => n57, Y => n98);
   U72 : AOI22X1 port map( A => DATA(5), B => n31, C => n47, D => 
                           tempData_5_port, Y => n57);
   U73 : INVX1 port map( A => PRGA_IN_5_port, Y => n56);
   U74 : OAI21X1 port map( A => n4, B => n58, C => n59, Y => n99);
   U75 : AOI22X1 port map( A => DATA(4), B => n31, C => n47, D => 
                           tempData_4_port, Y => n59);
   U76 : INVX1 port map( A => PRGA_IN_4_port, Y => n58);
   U77 : OAI21X1 port map( A => n4, B => n60, C => n61, Y => n100);
   U78 : AOI22X1 port map( A => DATA(3), B => n31, C => n47, D => 
                           tempData_3_port, Y => n61);
   U79 : INVX1 port map( A => PRGA_IN_3_port, Y => n60);
   U80 : OAI21X1 port map( A => n4, B => n62, C => n63, Y => n101);
   U81 : AOI22X1 port map( A => DATA(2), B => n31, C => n47, D => 
                           tempData_2_port, Y => n63);
   U82 : INVX1 port map( A => PRGA_IN_2_port, Y => n62);
   U83 : OAI21X1 port map( A => n4, B => n64, C => n65, Y => n102);
   U84 : AOI22X1 port map( A => DATA(1), B => n31, C => n47, D => 
                           tempData_1_port, Y => n65);
   U85 : INVX1 port map( A => PRGA_IN_1_port, Y => n64);
   U86 : OAI21X1 port map( A => n4, B => n66, C => n67, Y => n103);
   U87 : AOI22X1 port map( A => DATA(0), B => n31, C => n47, D => 
                           tempData_0_port, Y => n67);
   U88 : NAND2X1 port map( A => n14, B => state_2_port, Y => n42);
   U89 : INVX1 port map( A => n68, Y => n14);
   U90 : OAI21X1 port map( A => state_1_port, B => n69, C => n19, Y => n68);
   U91 : NAND2X1 port map( A => state_1_port, B => n69, Y => n19);
   U92 : NAND3X1 port map( A => n69, B => n10, C => n70, Y => n44);
   U93 : NOR2X1 port map( A => RST, B => n27, Y => n70);
   U94 : INVX1 port map( A => state_2_port, Y => n27);
   U95 : INVX1 port map( A => state_1_port, Y => n10);
   U96 : INVX1 port map( A => state_0_port, Y => n69);
   U97 : INVX1 port map( A => PRGA_IN_0_port, Y => n66);

end SYN_brbuffer;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_block_0 is

   port( CLK, RST, SERIAL_IN : in std_logic;  KEY_ERROR, PROG_ERROR : out 
         std_logic;  PLAINKEY : out std_logic_vector (63 downto 0);  RBUF_FULL,
         PARITY_ERROR : out std_logic);

end uart_rcv_block_0;

architecture SYN_struct1 of uart_rcv_block_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component uart_timer_0
      port( CLK, RST, TIMER_TRIG : in std_logic;  STOP_RCVING, SHIFT_STROBE : 
            out std_logic);
   end component;
   
   component keyreg_0
      port( CLK, RST, SBE, OE, RBUF_FULL : in std_logic;  RCV_DATA : in 
            std_logic_vector (7 downto 0);  PLAINKEY : out std_logic_vector (63
            downto 0);  KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR : out 
            std_logic);
   end component;
   
   component uart_sr_10bit_0
      port( CLK, RST, SHIFT_STROBE, SERIAL_IN : in std_logic;  LOAD_DATA : out 
            std_logic_vector (7 downto 0);  STOP_DATA : out std_logic_vector (1
            downto 0));
   end component;
   
   component uart_sb_check_0
      port( RST, CLK, SBC_CLR, SBC_EN : in std_logic;  STOP_DATA : in 
            std_logic_vector (1 downto 0);  SB_DETECT, SBE : out std_logic);
   end component;
   
   component uart_rcv_buf_full_0
      port( CLK, RST, CLR_RBUF, SET_RBUF_FULL : in std_logic;  RBUF_FULL : out 
            std_logic);
   end component;
   
   component uart_rcv_buf_0
      port( CLK, RST, LOAD_RBUF : in std_logic;  LOAD_DATA : in 
            std_logic_vector (7 downto 0);  RCV_DATA : out std_logic_vector (7 
            downto 0));
   end component;
   
   component uart_rcu_0
      port( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT : in std_logic;  
            RBUF_LOAD, TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR : 
            out std_logic);
   end component;
   
   component uart_error_0
      port( RST, CLK, RBUF_FULL, CHK_ERROR : in std_logic;  OE : out std_logic
            );
   end component;
   
   component uart_edge_detector_0
      port( CLK, RST, SERIAL_IN : in std_logic;  START_BIT : out std_logic);
   end component;
   
   signal RBUF_FULL_port, START_BIT, CHK_ERROR, OE, SB_DETECT, STOP_RCVING, 
      RBUF_LOAD, SBC_CLR, SBC_EN, SET_RBUF_FULL, TIMER_TRIG, LOAD_DATA_7_port, 
      LOAD_DATA_6_port, LOAD_DATA_5_port, LOAD_DATA_4_port, LOAD_DATA_3_port, 
      LOAD_DATA_2_port, LOAD_DATA_1_port, LOAD_DATA_0_port, RCV_DATA_7_port, 
      RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, RCV_DATA_3_port, 
      RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, CLR_RBUF, 
      STOP_DATA_1_port, STOP_DATA_0_port, SBE, SHIFT_STROBE, n1, n2 : std_logic
      ;

begin
   RBUF_FULL <= RBUF_FULL_port;
   
   U_0 : uart_edge_detector_0 port map( CLK => CLK, RST => n1, SERIAL_IN => 
                           SERIAL_IN, START_BIT => START_BIT);
   U_1 : uart_error_0 port map( RST => n1, CLK => CLK, RBUF_FULL => 
                           RBUF_FULL_port, CHK_ERROR => CHK_ERROR, OE => OE);
   U_2 : uart_rcu_0 port map( CLK => CLK, RST => n1, START_BIT => START_BIT, 
                           STOP_RCVING => STOP_RCVING, SB_DETECT => SB_DETECT, 
                           RBUF_LOAD => RBUF_LOAD, TIMER_TRIG => TIMER_TRIG, 
                           CHK_ERROR => CHK_ERROR, SET_RBUF_FULL => 
                           SET_RBUF_FULL, SBC_EN => SBC_EN, SBC_CLR => SBC_CLR)
                           ;
   U_3 : uart_rcv_buf_0 port map( CLK => CLK, RST => n1, LOAD_RBUF => RBUF_LOAD
                           , LOAD_DATA(7) => LOAD_DATA_7_port, LOAD_DATA(6) => 
                           LOAD_DATA_6_port, LOAD_DATA(5) => LOAD_DATA_5_port, 
                           LOAD_DATA(4) => LOAD_DATA_4_port, LOAD_DATA(3) => 
                           LOAD_DATA_3_port, LOAD_DATA(2) => LOAD_DATA_2_port, 
                           LOAD_DATA(1) => LOAD_DATA_1_port, LOAD_DATA(0) => 
                           LOAD_DATA_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port);
   U_4 : uart_rcv_buf_full_0 port map( CLK => CLK, RST => n1, CLR_RBUF => 
                           CLR_RBUF, SET_RBUF_FULL => SET_RBUF_FULL, RBUF_FULL 
                           => RBUF_FULL_port);
   U_5 : uart_sb_check_0 port map( RST => n1, CLK => CLK, SBC_CLR => SBC_CLR, 
                           SBC_EN => SBC_EN, STOP_DATA(1) => STOP_DATA_1_port, 
                           STOP_DATA(0) => STOP_DATA_0_port, SB_DETECT => 
                           SB_DETECT, SBE => SBE);
   U_6 : uart_sr_10bit_0 port map( CLK => CLK, RST => n1, SHIFT_STROBE => 
                           SHIFT_STROBE, SERIAL_IN => SERIAL_IN, LOAD_DATA(7) 
                           => LOAD_DATA_7_port, LOAD_DATA(6) => 
                           LOAD_DATA_6_port, LOAD_DATA(5) => LOAD_DATA_5_port, 
                           LOAD_DATA(4) => LOAD_DATA_4_port, LOAD_DATA(3) => 
                           LOAD_DATA_3_port, LOAD_DATA(2) => LOAD_DATA_2_port, 
                           LOAD_DATA(1) => LOAD_DATA_1_port, LOAD_DATA(0) => 
                           LOAD_DATA_0_port, STOP_DATA(1) => STOP_DATA_1_port, 
                           STOP_DATA(0) => STOP_DATA_0_port);
   U_8 : keyreg_0 port map( CLK => CLK, RST => n1, SBE => SBE, OE => OE, 
                           RBUF_FULL => RBUF_FULL_port, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           PLAINKEY(63) => PLAINKEY(63), PLAINKEY(62) => 
                           PLAINKEY(62), PLAINKEY(61) => PLAINKEY(61), 
                           PLAINKEY(60) => PLAINKEY(60), PLAINKEY(59) => 
                           PLAINKEY(59), PLAINKEY(58) => PLAINKEY(58), 
                           PLAINKEY(57) => PLAINKEY(57), PLAINKEY(56) => 
                           PLAINKEY(56), PLAINKEY(55) => PLAINKEY(55), 
                           PLAINKEY(54) => PLAINKEY(54), PLAINKEY(53) => 
                           PLAINKEY(53), PLAINKEY(52) => PLAINKEY(52), 
                           PLAINKEY(51) => PLAINKEY(51), PLAINKEY(50) => 
                           PLAINKEY(50), PLAINKEY(49) => PLAINKEY(49), 
                           PLAINKEY(48) => PLAINKEY(48), PLAINKEY(47) => 
                           PLAINKEY(47), PLAINKEY(46) => PLAINKEY(46), 
                           PLAINKEY(45) => PLAINKEY(45), PLAINKEY(44) => 
                           PLAINKEY(44), PLAINKEY(43) => PLAINKEY(43), 
                           PLAINKEY(42) => PLAINKEY(42), PLAINKEY(41) => 
                           PLAINKEY(41), PLAINKEY(40) => PLAINKEY(40), 
                           PLAINKEY(39) => PLAINKEY(39), PLAINKEY(38) => 
                           PLAINKEY(38), PLAINKEY(37) => PLAINKEY(37), 
                           PLAINKEY(36) => PLAINKEY(36), PLAINKEY(35) => 
                           PLAINKEY(35), PLAINKEY(34) => PLAINKEY(34), 
                           PLAINKEY(33) => PLAINKEY(33), PLAINKEY(32) => 
                           PLAINKEY(32), PLAINKEY(31) => PLAINKEY(31), 
                           PLAINKEY(30) => PLAINKEY(30), PLAINKEY(29) => 
                           PLAINKEY(29), PLAINKEY(28) => PLAINKEY(28), 
                           PLAINKEY(27) => PLAINKEY(27), PLAINKEY(26) => 
                           PLAINKEY(26), PLAINKEY(25) => PLAINKEY(25), 
                           PLAINKEY(24) => PLAINKEY(24), PLAINKEY(23) => 
                           PLAINKEY(23), PLAINKEY(22) => PLAINKEY(22), 
                           PLAINKEY(21) => PLAINKEY(21), PLAINKEY(20) => 
                           PLAINKEY(20), PLAINKEY(19) => PLAINKEY(19), 
                           PLAINKEY(18) => PLAINKEY(18), PLAINKEY(17) => 
                           PLAINKEY(17), PLAINKEY(16) => PLAINKEY(16), 
                           PLAINKEY(15) => PLAINKEY(15), PLAINKEY(14) => 
                           PLAINKEY(14), PLAINKEY(13) => PLAINKEY(13), 
                           PLAINKEY(12) => PLAINKEY(12), PLAINKEY(11) => 
                           PLAINKEY(11), PLAINKEY(10) => PLAINKEY(10), 
                           PLAINKEY(9) => PLAINKEY(9), PLAINKEY(8) => 
                           PLAINKEY(8), PLAINKEY(7) => PLAINKEY(7), PLAINKEY(6)
                           => PLAINKEY(6), PLAINKEY(5) => PLAINKEY(5), 
                           PLAINKEY(4) => PLAINKEY(4), PLAINKEY(3) => 
                           PLAINKEY(3), PLAINKEY(2) => PLAINKEY(2), PLAINKEY(1)
                           => PLAINKEY(1), PLAINKEY(0) => PLAINKEY(0), 
                           KEY_ERROR => KEY_ERROR, PROG_ERROR => PROG_ERROR, 
                           CLR_RBUFF => CLR_RBUF, PARITY_ERROR => PARITY_ERROR)
                           ;
   U_7 : uart_timer_0 port map( CLK => CLK, RST => n1, TIMER_TRIG => TIMER_TRIG
                           , STOP_RCVING => STOP_RCVING, SHIFT_STROBE => 
                           SHIFT_STROBE);
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct1;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_0 is

   port( KEY : in std_logic_vector (63 downto 0);  CLK, RST, KEY_ERROR, 
         BYTE_READY : in std_logic;  BYTE : in std_logic_vector (7 downto 0);  
         OPCODE : in std_logic_vector (1 downto 0);  DATA_IN : in 
         std_logic_vector (7 downto 0);  PROCESSED_DATA : out std_logic_vector 
         (7 downto 0);  PDATA_READY, W_ENABLE, R_ENABLE : out std_logic;  ADDR,
         DATA : out std_logic_vector (7 downto 0));

end KSA_0;

architecture SYN_bksa of KSA_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUFX1
      port( A, EN : in std_logic;  Y : out std_logic);
   end component;
   
   component KSA_0_DW01_add_2
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_0_DW01_add_3
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_0_DW01_inc_2
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_0_DW01_inc_1
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_0_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_0_DW01_add_1
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_0_DW01_add_0
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, PROCESSED_DATA_5_port, 
      PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, PROCESSED_DATA_2_port, 
      PROCESSED_DATA_1_port, PROCESSED_DATA_0_port, W_ENABLE_port, 
      R_ENABLE_port, ADDR_7_port, ADDR_6_port, ADDR_5_port, ADDR_4_port, 
      ADDR_3_port, ADDR_2_port, ADDR_1_port, ADDR_0_port, DATA_7_port, 
      DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, DATA_2_port, 
      DATA_1_port, DATA_0_port, state_4_port, state_3_port, state_2_port, 
      state_1_port, state_0_port, si_7_port, si_6_port, si_5_port, si_4_port, 
      si_3_port, si_2_port, si_1_port, si_0_port, sj_7_port, sj_6_port, 
      sj_5_port, sj_4_port, sj_3_port, sj_2_port, sj_1_port, sj_0_port, 
      currentProcessedData_7_port, currentProcessedData_6_port, 
      currentProcessedData_5_port, currentProcessedData_4_port, 
      currentProcessedData_3_port, currentProcessedData_2_port, 
      currentProcessedData_1_port, currentProcessedData_0_port, 
      nextState_4_port, nextState_3_port, nextState_2_port, nextState_1_port, 
      nextState_0_port, inti_7_port, inti_6_port, inti_5_port, inti_4_port, 
      inti_3_port, inti_2_port, inti_1_port, inti_0_port, intj_7_port, 
      intj_6_port, intj_5_port, intj_4_port, intj_3_port, intj_2_port, 
      intj_1_port, intj_0_port, keyi_2_port, keyi_1_port, keyi_0_port, 
      permuteComplete, temp_7_port, temp_6_port, temp_5_port, temp_4_port, 
      temp_3_port, temp_2_port, temp_1_port, temp_0_port, extratemp_7_port, 
      extratemp_6_port, extratemp_5_port, extratemp_4_port, extratemp_3_port, 
      extratemp_2_port, extratemp_1_port, extratemp_0_port, 
      nextProcessedData_7_port, nextProcessedData_6_port, 
      nextProcessedData_5_port, nextProcessedData_4_port, 
      nextProcessedData_3_port, nextProcessedData_2_port, 
      nextProcessedData_1_port, nextProcessedData_0_port, keyTable_0_7_port, 
      keyTable_0_6_port, keyTable_0_5_port, keyTable_0_4_port, 
      keyTable_0_3_port, keyTable_0_2_port, keyTable_0_1_port, 
      keyTable_0_0_port, keyTable_1_7_port, keyTable_1_6_port, 
      keyTable_1_5_port, keyTable_1_4_port, keyTable_1_3_port, 
      keyTable_1_2_port, keyTable_1_1_port, keyTable_1_0_port, 
      keyTable_2_7_port, keyTable_2_6_port, keyTable_2_5_port, 
      keyTable_2_4_port, keyTable_2_3_port, keyTable_2_2_port, 
      keyTable_2_1_port, keyTable_2_0_port, keyTable_3_7_port, 
      keyTable_3_6_port, keyTable_3_5_port, keyTable_3_4_port, 
      keyTable_3_3_port, keyTable_3_2_port, keyTable_3_1_port, 
      keyTable_3_0_port, keyTable_4_7_port, keyTable_4_6_port, 
      keyTable_4_5_port, keyTable_4_4_port, keyTable_4_3_port, 
      keyTable_4_2_port, keyTable_4_1_port, keyTable_4_0_port, 
      keyTable_5_7_port, keyTable_5_6_port, keyTable_5_5_port, 
      keyTable_5_4_port, keyTable_5_3_port, keyTable_5_2_port, 
      keyTable_5_1_port, keyTable_5_0_port, keyTable_6_7_port, 
      keyTable_6_6_port, keyTable_6_5_port, keyTable_6_4_port, 
      keyTable_6_3_port, keyTable_6_2_port, keyTable_6_1_port, 
      keyTable_6_0_port, keyTable_7_7_port, keyTable_7_6_port, 
      keyTable_7_5_port, keyTable_7_4_port, keyTable_7_3_port, 
      keyTable_7_2_port, keyTable_7_1_port, keyTable_7_0_port, delaydata_7_port
      , delaydata_6_port, delaydata_5_port, delaydata_4_port, delaydata_3_port,
      delaydata_2_port, delaydata_1_port, delaydata_0_port, 
      prefillCounter_7_port, prefillCounter_6_port, prefillCounter_5_port, 
      prefillCounter_4_port, prefillCounter_3_port, prefillCounter_2_port, 
      prefillCounter_1_port, prefillCounter_0_port, faddr_7_port, faddr_6_port,
      faddr_5_port, faddr_4_port, faddr_3_port, faddr_2_port, faddr_1_port, 
      faddr_0_port, nfaddr_7_port, nfaddr_6_port, nfaddr_5_port, nfaddr_4_port,
      nfaddr_3_port, nfaddr_2_port, nfaddr_1_port, nfaddr_0_port, fdata_7_port,
      fdata_6_port, fdata_5_port, fdata_4_port, fdata_3_port, fdata_2_port, 
      fdata_1_port, fdata_0_port, nfdata_7_port, nfdata_6_port, nfdata_5_port, 
      nfdata_4_port, nfdata_3_port, nfdata_2_port, nfdata_1_port, nfdata_0_port
      , fw_enable, fr_enable, N407, N408, N409, N410, N411, N412, N413, N414, 
      N424, N425, N426, N427, N428, N429, N430, N431, N442, N443, N444, N445, 
      N446, N447, N448, N472, N473, N474, N475, N476, N477, N478, N479, N480, 
      N481, N482, N483, N484, N485, N486, N487, N496, N497, N498, N499, N500, 
      N501, N502, N503, N512, N513, N514, N515, N516, N517, N518, N519, N520, 
      N521, N522, N523, N524, N525, N526, N527, N456, N455, N454, N453, N452, 
      N451, N450, N449, n3, n4, n5, n6, n7, n8, n9, n10, n12, n14, n15, n16, 
      n17, n20, n22, n24, n27, n29, n32, n34, n37, n39, n42, n44, n47, n49, n52
      , n54, n62, n64, n117, n121, n122, n129, n131, n135, n136, n141, n151, 
      n160, n161, n172, n175, n177, n180, n185, n187, n188, n196, n203, n206, 
      n208, n210, n212, n214, n216, n218, n220, n230, n235, n237, n238, n239, 
      n240, n241, n244, n246, n247, n249, n250, n252, n253, n255, n256, n258, 
      n259, n261, n262, n264, n265, n267, n268, n270, n271, n275, n277, n280, 
      n282, n285, n287, n290, n292, n295, n297, n300, n302, n305, n307, n311, 
      n317, n318, n326, n327, n329, n331, n333, n335, n337, n339, n341, n343, 
      n345, n347, n349, n351, n353, n355, n357, n359, n361, n363, n365, n367, 
      n369, n371, n373, n375, n377, n379, n381, n383, n385, n387, n389, n391, 
      n393, n395, n397, n399, n401, n403, n405, n407_port, n409_port, n411_port
      , n413_port, n415, n417, n419, n421, n423, n425_port, n427_port, 
      n429_port, n431_port, n433, n435, n437, n439, n441, n443_port, n445_port,
      n447_port, n449_port, n451_port, n453_port, n455_port, n458, n459, n462, 
      n463, n465, n467, n469, n471, n473_port, n475_port, n480_port, n482_port,
      n488, n498_port, n500_port, n501_port, n503_port, n504, n505, n506, n507,
      n509, n512_port, n514_port, n516_port, n518_port, n520_port, n522_port, 
      n524_port, n528, n540, n541, n542, n543, n545, n547, n549, n551, n553, 
      n555, n557, n562, n569, n571, n572, n575, n577, n579, n581, n592, n594, 
      n600, n604, n605, n606, n610, n612, n614, n616, n618, n624, n626, n629, 
      n630, n632, n636, n637, n638, n648, n649, n650, n651, n692, n701, n746, 
      n748, n750, n752, n754, n756, n758, n760, n761, n762, n763, n764, n765, 
      n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, 
      n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, 
      n790, n791, n864, n865, n866, n867, n868, n869, n870, n871, n883, n884, 
      n885, n886, n887, n888, n889, n890, n916, n917, n918, n919, n920, n921, 
      n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, 
      n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, 
      n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, 
      n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
      n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, 
      n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, 
      n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, 
      n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, 
      n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, 
      n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, 
      n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, 
      n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, 
      n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, 
      n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
      n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
      n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
      n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, 
      n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
      n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
      n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
      n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
      n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, 
      n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
      n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
      n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
      n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
      n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, 
      n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, 
      n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, 
      n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
      n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, 
      n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, 
      n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, 
      n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, 
      n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, 
      n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, 
      n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, 
      n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
      n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, 
      n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, 
      n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, 
      n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, 
      n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, 
      n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, 
      n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, 
      n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, 
      n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, 
      n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, 
      n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, 
      n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
      n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, 
      n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, 
      n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
      n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, 
      n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, 
      n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, 
      n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, 
      n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, 
      n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, 
      n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, 
      n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, 
      n_1021, n_1022, n_1023, n_1024 : std_logic;

begin
   PROCESSED_DATA <= ( PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, 
      PROCESSED_DATA_5_port, PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, 
      PROCESSED_DATA_2_port, PROCESSED_DATA_1_port, PROCESSED_DATA_0_port );
   W_ENABLE <= W_ENABLE_port;
   R_ENABLE <= R_ENABLE_port;
   ADDR <= ( ADDR_7_port, ADDR_6_port, ADDR_5_port, ADDR_4_port, ADDR_3_port, 
      ADDR_2_port, ADDR_1_port, ADDR_0_port );
   DATA <= ( DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, 
      DATA_2_port, DATA_1_port, DATA_0_port );
   
   n1604 <= '0';
   n1603 <= '0';
   prefillCounter_reg_0_inst : DFFPOSX1 port map( D => n986, CLK => CLK, Q => 
                           prefillCounter_0_port);
   permuteComplete_reg : DFFPOSX1 port map( D => n1002, CLK => CLK, Q => 
                           permuteComplete);
   extratemp_reg_7_inst : DFFPOSX1 port map( D => n482_port, CLK => CLK, Q => 
                           extratemp_7_port);
   extratemp_reg_6_inst : DFFPOSX1 port map( D => n480_port, CLK => CLK, Q => 
                           extratemp_6_port);
   extratemp_reg_5_inst : DFFPOSX1 port map( D => n475_port, CLK => CLK, Q => 
                           extratemp_5_port);
   extratemp_reg_4_inst : DFFPOSX1 port map( D => n473_port, CLK => CLK, Q => 
                           extratemp_4_port);
   extratemp_reg_3_inst : DFFPOSX1 port map( D => n471, CLK => CLK, Q => 
                           extratemp_3_port);
   extratemp_reg_2_inst : DFFPOSX1 port map( D => n469, CLK => CLK, Q => 
                           extratemp_2_port);
   extratemp_reg_1_inst : DFFPOSX1 port map( D => n467, CLK => CLK, Q => 
                           extratemp_1_port);
   extratemp_reg_0_inst : DFFPOSX1 port map( D => n465, CLK => CLK, Q => 
                           extratemp_0_port);
   keyTable_reg_7_0_inst : DFFPOSX1 port map( D => n1093, CLK => CLK, Q => 
                           keyTable_7_0_port);
   keyTable_reg_7_1_inst : DFFPOSX1 port map( D => n1092, CLK => CLK, Q => 
                           keyTable_7_1_port);
   keyTable_reg_7_2_inst : DFFPOSX1 port map( D => n1091, CLK => CLK, Q => 
                           keyTable_7_2_port);
   keyTable_reg_7_3_inst : DFFPOSX1 port map( D => n1090, CLK => CLK, Q => 
                           keyTable_7_3_port);
   keyTable_reg_7_4_inst : DFFPOSX1 port map( D => n1089, CLK => CLK, Q => 
                           keyTable_7_4_port);
   keyTable_reg_7_5_inst : DFFPOSX1 port map( D => n1088, CLK => CLK, Q => 
                           keyTable_7_5_port);
   keyTable_reg_7_6_inst : DFFPOSX1 port map( D => n1087, CLK => CLK, Q => 
                           keyTable_7_6_port);
   keyTable_reg_7_7_inst : DFFPOSX1 port map( D => n1086, CLK => CLK, Q => 
                           keyTable_7_7_port);
   keyTable_reg_6_0_inst : DFFPOSX1 port map( D => n1085, CLK => CLK, Q => 
                           keyTable_6_0_port);
   keyTable_reg_6_1_inst : DFFPOSX1 port map( D => n1084, CLK => CLK, Q => 
                           keyTable_6_1_port);
   keyTable_reg_6_2_inst : DFFPOSX1 port map( D => n1083, CLK => CLK, Q => 
                           keyTable_6_2_port);
   keyTable_reg_6_3_inst : DFFPOSX1 port map( D => n1082, CLK => CLK, Q => 
                           keyTable_6_3_port);
   keyTable_reg_6_4_inst : DFFPOSX1 port map( D => n1081, CLK => CLK, Q => 
                           keyTable_6_4_port);
   keyTable_reg_6_5_inst : DFFPOSX1 port map( D => n1080, CLK => CLK, Q => 
                           keyTable_6_5_port);
   keyTable_reg_6_6_inst : DFFPOSX1 port map( D => n1079, CLK => CLK, Q => 
                           keyTable_6_6_port);
   keyTable_reg_6_7_inst : DFFPOSX1 port map( D => n1078, CLK => CLK, Q => 
                           keyTable_6_7_port);
   keyTable_reg_5_0_inst : DFFPOSX1 port map( D => n1077, CLK => CLK, Q => 
                           keyTable_5_0_port);
   keyTable_reg_5_1_inst : DFFPOSX1 port map( D => n1076, CLK => CLK, Q => 
                           keyTable_5_1_port);
   keyTable_reg_5_2_inst : DFFPOSX1 port map( D => n1075, CLK => CLK, Q => 
                           keyTable_5_2_port);
   keyTable_reg_5_3_inst : DFFPOSX1 port map( D => n1074, CLK => CLK, Q => 
                           keyTable_5_3_port);
   keyTable_reg_5_4_inst : DFFPOSX1 port map( D => n1073, CLK => CLK, Q => 
                           keyTable_5_4_port);
   keyTable_reg_5_5_inst : DFFPOSX1 port map( D => n1072, CLK => CLK, Q => 
                           keyTable_5_5_port);
   keyTable_reg_5_6_inst : DFFPOSX1 port map( D => n1071, CLK => CLK, Q => 
                           keyTable_5_6_port);
   keyTable_reg_5_7_inst : DFFPOSX1 port map( D => n1070, CLK => CLK, Q => 
                           keyTable_5_7_port);
   keyTable_reg_4_0_inst : DFFPOSX1 port map( D => n1069, CLK => CLK, Q => 
                           keyTable_4_0_port);
   keyTable_reg_4_1_inst : DFFPOSX1 port map( D => n1068, CLK => CLK, Q => 
                           keyTable_4_1_port);
   keyTable_reg_4_2_inst : DFFPOSX1 port map( D => n1067, CLK => CLK, Q => 
                           keyTable_4_2_port);
   keyTable_reg_4_3_inst : DFFPOSX1 port map( D => n1066, CLK => CLK, Q => 
                           keyTable_4_3_port);
   keyTable_reg_4_4_inst : DFFPOSX1 port map( D => n1065, CLK => CLK, Q => 
                           keyTable_4_4_port);
   keyTable_reg_4_5_inst : DFFPOSX1 port map( D => n1064, CLK => CLK, Q => 
                           keyTable_4_5_port);
   keyTable_reg_4_6_inst : DFFPOSX1 port map( D => n1063, CLK => CLK, Q => 
                           keyTable_4_6_port);
   keyTable_reg_4_7_inst : DFFPOSX1 port map( D => n1062, CLK => CLK, Q => 
                           keyTable_4_7_port);
   keyTable_reg_3_0_inst : DFFPOSX1 port map( D => n1061, CLK => CLK, Q => 
                           keyTable_3_0_port);
   keyTable_reg_3_1_inst : DFFPOSX1 port map( D => n1060, CLK => CLK, Q => 
                           keyTable_3_1_port);
   keyTable_reg_3_2_inst : DFFPOSX1 port map( D => n1059, CLK => CLK, Q => 
                           keyTable_3_2_port);
   keyTable_reg_3_3_inst : DFFPOSX1 port map( D => n1058, CLK => CLK, Q => 
                           keyTable_3_3_port);
   keyTable_reg_3_4_inst : DFFPOSX1 port map( D => n1057, CLK => CLK, Q => 
                           keyTable_3_4_port);
   keyTable_reg_3_5_inst : DFFPOSX1 port map( D => n1056, CLK => CLK, Q => 
                           keyTable_3_5_port);
   keyTable_reg_3_6_inst : DFFPOSX1 port map( D => n1055, CLK => CLK, Q => 
                           keyTable_3_6_port);
   keyTable_reg_3_7_inst : DFFPOSX1 port map( D => n1054, CLK => CLK, Q => 
                           keyTable_3_7_port);
   keyTable_reg_2_0_inst : DFFPOSX1 port map( D => n1053, CLK => CLK, Q => 
                           keyTable_2_0_port);
   keyTable_reg_2_1_inst : DFFPOSX1 port map( D => n1052, CLK => CLK, Q => 
                           keyTable_2_1_port);
   keyTable_reg_2_2_inst : DFFPOSX1 port map( D => n1051, CLK => CLK, Q => 
                           keyTable_2_2_port);
   keyTable_reg_2_3_inst : DFFPOSX1 port map( D => n1050, CLK => CLK, Q => 
                           keyTable_2_3_port);
   keyTable_reg_2_4_inst : DFFPOSX1 port map( D => n1049, CLK => CLK, Q => 
                           keyTable_2_4_port);
   keyTable_reg_2_5_inst : DFFPOSX1 port map( D => n1048, CLK => CLK, Q => 
                           keyTable_2_5_port);
   keyTable_reg_2_6_inst : DFFPOSX1 port map( D => n1047, CLK => CLK, Q => 
                           keyTable_2_6_port);
   keyTable_reg_2_7_inst : DFFPOSX1 port map( D => n1046, CLK => CLK, Q => 
                           keyTable_2_7_port);
   keyTable_reg_1_0_inst : DFFPOSX1 port map( D => n1045, CLK => CLK, Q => 
                           keyTable_1_0_port);
   keyTable_reg_1_1_inst : DFFPOSX1 port map( D => n1044, CLK => CLK, Q => 
                           keyTable_1_1_port);
   keyTable_reg_1_2_inst : DFFPOSX1 port map( D => n1043, CLK => CLK, Q => 
                           keyTable_1_2_port);
   keyTable_reg_1_3_inst : DFFPOSX1 port map( D => n1042, CLK => CLK, Q => 
                           keyTable_1_3_port);
   keyTable_reg_1_4_inst : DFFPOSX1 port map( D => n1041, CLK => CLK, Q => 
                           keyTable_1_4_port);
   keyTable_reg_1_5_inst : DFFPOSX1 port map( D => n1040, CLK => CLK, Q => 
                           keyTable_1_5_port);
   keyTable_reg_1_6_inst : DFFPOSX1 port map( D => n1039, CLK => CLK, Q => 
                           keyTable_1_6_port);
   keyTable_reg_0_6_inst : DFFPOSX1 port map( D => n1038, CLK => CLK, Q => 
                           keyTable_0_6_port);
   keyTable_reg_0_5_inst : DFFPOSX1 port map( D => n1037, CLK => CLK, Q => 
                           keyTable_0_5_port);
   keyTable_reg_0_4_inst : DFFPOSX1 port map( D => n1036, CLK => CLK, Q => 
                           keyTable_0_4_port);
   keyTable_reg_0_3_inst : DFFPOSX1 port map( D => n1035, CLK => CLK, Q => 
                           keyTable_0_3_port);
   keyTable_reg_0_2_inst : DFFPOSX1 port map( D => n1034, CLK => CLK, Q => 
                           keyTable_0_2_port);
   keyTable_reg_0_1_inst : DFFPOSX1 port map( D => n1033, CLK => CLK, Q => 
                           keyTable_0_1_port);
   keyTable_reg_0_0_inst : DFFPOSX1 port map( D => n1032, CLK => CLK, Q => 
                           keyTable_0_0_port);
   keyTable_reg_1_7_inst : DFFPOSX1 port map( D => n1031, CLK => CLK, Q => 
                           keyTable_1_7_port);
   keyTable_reg_0_7_inst : DFFPOSX1 port map( D => n1030, CLK => CLK, Q => 
                           keyTable_0_7_port);
   prefillCounter_reg_7_inst : DFFPOSX1 port map( D => n987, CLK => CLK, Q => 
                           prefillCounter_7_port);
   prefillCounter_reg_1_inst : DFFPOSX1 port map( D => n988, CLK => CLK, Q => 
                           prefillCounter_1_port);
   prefillCounter_reg_2_inst : DFFPOSX1 port map( D => n989, CLK => CLK, Q => 
                           prefillCounter_2_port);
   prefillCounter_reg_3_inst : DFFPOSX1 port map( D => n990, CLK => CLK, Q => 
                           prefillCounter_3_port);
   prefillCounter_reg_4_inst : DFFPOSX1 port map( D => n991, CLK => CLK, Q => 
                           prefillCounter_4_port);
   prefillCounter_reg_5_inst : DFFPOSX1 port map( D => n992, CLK => CLK, Q => 
                           prefillCounter_5_port);
   prefillCounter_reg_6_inst : DFFPOSX1 port map( D => n993, CLK => CLK, Q => 
                           prefillCounter_6_port);
   temp_reg_7_inst : DFFPOSX1 port map( D => n1029, CLK => CLK, Q => 
                           temp_7_port);
   temp_reg_0_inst : DFFPOSX1 port map( D => n1022, CLK => CLK, Q => 
                           temp_0_port);
   temp_reg_1_inst : DFFPOSX1 port map( D => n1023, CLK => CLK, Q => 
                           temp_1_port);
   temp_reg_2_inst : DFFPOSX1 port map( D => n1024, CLK => CLK, Q => 
                           temp_2_port);
   temp_reg_3_inst : DFFPOSX1 port map( D => n1025, CLK => CLK, Q => 
                           temp_3_port);
   temp_reg_4_inst : DFFPOSX1 port map( D => n1026, CLK => CLK, Q => 
                           temp_4_port);
   temp_reg_5_inst : DFFPOSX1 port map( D => n1027, CLK => CLK, Q => 
                           temp_5_port);
   temp_reg_6_inst : DFFPOSX1 port map( D => n1028, CLK => CLK, Q => 
                           temp_6_port);
   delaydata_reg_7_inst : DFFPOSX1 port map( D => n383, CLK => CLK, Q => 
                           delaydata_7_port);
   delaydata_reg_0_inst : DFFPOSX1 port map( D => n411_port, CLK => CLK, Q => 
                           delaydata_0_port);
   delaydata_reg_1_inst : DFFPOSX1 port map( D => n407_port, CLK => CLK, Q => 
                           delaydata_1_port);
   delaydata_reg_2_inst : DFFPOSX1 port map( D => n403, CLK => CLK, Q => 
                           delaydata_2_port);
   delaydata_reg_3_inst : DFFPOSX1 port map( D => n399, CLK => CLK, Q => 
                           delaydata_3_port);
   delaydata_reg_4_inst : DFFPOSX1 port map( D => n395, CLK => CLK, Q => 
                           delaydata_4_port);
   delaydata_reg_5_inst : DFFPOSX1 port map( D => n391, CLK => CLK, Q => 
                           delaydata_5_port);
   delaydata_reg_6_inst : DFFPOSX1 port map( D => n387, CLK => CLK, Q => 
                           delaydata_6_port);
   intj_reg_7_inst : DFFPOSX1 port map( D => n1018, CLK => CLK, Q => 
                           intj_7_port);
   intj_reg_0_inst : DFFPOSX1 port map( D => n1011, CLK => CLK, Q => 
                           intj_0_port);
   intj_reg_1_inst : DFFPOSX1 port map( D => n1012, CLK => CLK, Q => 
                           intj_1_port);
   intj_reg_2_inst : DFFPOSX1 port map( D => n1013, CLK => CLK, Q => 
                           intj_2_port);
   intj_reg_3_inst : DFFPOSX1 port map( D => n1014, CLK => CLK, Q => 
                           intj_3_port);
   intj_reg_4_inst : DFFPOSX1 port map( D => n1015, CLK => CLK, Q => 
                           intj_4_port);
   intj_reg_5_inst : DFFPOSX1 port map( D => n1016, CLK => CLK, Q => 
                           intj_5_port);
   intj_reg_6_inst : DFFPOSX1 port map( D => n1017, CLK => CLK, Q => 
                           intj_6_port);
   keyi_reg_2_inst : DFFPOSX1 port map( D => n1019, CLK => CLK, Q => 
                           keyi_2_port);
   keyi_reg_1_inst : DFFPOSX1 port map( D => n1020, CLK => CLK, Q => 
                           keyi_1_port);
   keyi_reg_0_inst : DFFPOSX1 port map( D => n1021, CLK => CLK, Q => 
                           keyi_0_port);
   inti_reg_7_inst : DFFPOSX1 port map( D => n437, CLK => CLK, Q => inti_7_port
                           );
   inti_reg_0_inst : DFFPOSX1 port map( D => n423, CLK => CLK, Q => inti_0_port
                           );
   inti_reg_1_inst : DFFPOSX1 port map( D => n425_port, CLK => CLK, Q => 
                           inti_1_port);
   inti_reg_2_inst : DFFPOSX1 port map( D => n427_port, CLK => CLK, Q => 
                           inti_2_port);
   inti_reg_3_inst : DFFPOSX1 port map( D => n429_port, CLK => CLK, Q => 
                           inti_3_port);
   inti_reg_4_inst : DFFPOSX1 port map( D => n431_port, CLK => CLK, Q => 
                           inti_4_port);
   inti_reg_5_inst : DFFPOSX1 port map( D => n433, CLK => CLK, Q => inti_5_port
                           );
   inti_reg_6_inst : DFFPOSX1 port map( D => n435, CLK => CLK, Q => inti_6_port
                           );
   PROCESSED_DATA_reg_0_inst : DFFPOSX1 port map( D => n1094, CLK => CLK, Q => 
                           PROCESSED_DATA_0_port);
   PROCESSED_DATA_reg_1_inst : DFFPOSX1 port map( D => n1095, CLK => CLK, Q => 
                           PROCESSED_DATA_1_port);
   PROCESSED_DATA_reg_2_inst : DFFPOSX1 port map( D => n1096, CLK => CLK, Q => 
                           PROCESSED_DATA_2_port);
   PROCESSED_DATA_reg_3_inst : DFFPOSX1 port map( D => n1097, CLK => CLK, Q => 
                           PROCESSED_DATA_3_port);
   PROCESSED_DATA_reg_4_inst : DFFPOSX1 port map( D => n1098, CLK => CLK, Q => 
                           PROCESSED_DATA_4_port);
   PROCESSED_DATA_reg_5_inst : DFFPOSX1 port map( D => n1099, CLK => CLK, Q => 
                           PROCESSED_DATA_5_port);
   PROCESSED_DATA_reg_6_inst : DFFPOSX1 port map( D => n1100, CLK => CLK, Q => 
                           PROCESSED_DATA_6_port);
   PROCESSED_DATA_reg_7_inst : DFFPOSX1 port map( D => n1101, CLK => CLK, Q => 
                           PROCESSED_DATA_7_port);
   faddr_reg_7_inst : DFFPOSX1 port map( D => n1102, CLK => CLK, Q => 
                           faddr_7_port);
   ADDR_reg_7_inst : DFFPOSX1 port map( D => n1103, CLK => CLK, Q => 
                           ADDR_7_port);
   faddr_reg_6_inst : DFFPOSX1 port map( D => n1104, CLK => CLK, Q => 
                           faddr_6_port);
   ADDR_reg_6_inst : DFFPOSX1 port map( D => n1105, CLK => CLK, Q => 
                           ADDR_6_port);
   faddr_reg_5_inst : DFFPOSX1 port map( D => n1106, CLK => CLK, Q => 
                           faddr_5_port);
   ADDR_reg_5_inst : DFFPOSX1 port map( D => n1107, CLK => CLK, Q => 
                           ADDR_5_port);
   faddr_reg_4_inst : DFFPOSX1 port map( D => n1108, CLK => CLK, Q => 
                           faddr_4_port);
   ADDR_reg_4_inst : DFFPOSX1 port map( D => n1109, CLK => CLK, Q => 
                           ADDR_4_port);
   faddr_reg_3_inst : DFFPOSX1 port map( D => n1110, CLK => CLK, Q => 
                           faddr_3_port);
   ADDR_reg_3_inst : DFFPOSX1 port map( D => n1111, CLK => CLK, Q => 
                           ADDR_3_port);
   faddr_reg_2_inst : DFFPOSX1 port map( D => n1112, CLK => CLK, Q => 
                           faddr_2_port);
   ADDR_reg_2_inst : DFFPOSX1 port map( D => n1113, CLK => CLK, Q => 
                           ADDR_2_port);
   faddr_reg_1_inst : DFFPOSX1 port map( D => n1114, CLK => CLK, Q => 
                           faddr_1_port);
   ADDR_reg_1_inst : DFFPOSX1 port map( D => n1115, CLK => CLK, Q => 
                           ADDR_1_port);
   faddr_reg_0_inst : DFFPOSX1 port map( D => n1116, CLK => CLK, Q => 
                           faddr_0_port);
   ADDR_reg_0_inst : DFFPOSX1 port map( D => n1117, CLK => CLK, Q => 
                           ADDR_0_port);
   fdata_reg_7_inst : DFFPOSX1 port map( D => n1118, CLK => CLK, Q => 
                           fdata_7_port);
   fdata_reg_6_inst : DFFPOSX1 port map( D => n1119, CLK => CLK, Q => 
                           fdata_6_port);
   fdata_reg_5_inst : DFFPOSX1 port map( D => n1120, CLK => CLK, Q => 
                           fdata_5_port);
   fdata_reg_4_inst : DFFPOSX1 port map( D => n1121, CLK => CLK, Q => 
                           fdata_4_port);
   fdata_reg_3_inst : DFFPOSX1 port map( D => n1122, CLK => CLK, Q => 
                           fdata_3_port);
   fdata_reg_2_inst : DFFPOSX1 port map( D => n1123, CLK => CLK, Q => 
                           fdata_2_port);
   fdata_reg_1_inst : DFFPOSX1 port map( D => n1124, CLK => CLK, Q => 
                           fdata_1_port);
   fdata_reg_0_inst : DFFPOSX1 port map( D => n1125, CLK => CLK, Q => 
                           fdata_0_port);
   fw_enable_reg : DFFPOSX1 port map( D => n1126, CLK => CLK, Q => fw_enable);
   fr_enable_reg : DFFPOSX1 port map( D => n1127, CLK => CLK, Q => fr_enable);
   W_ENABLE_reg : DFFPOSX1 port map( D => n1128, CLK => CLK, Q => W_ENABLE_port
                           );
   R_ENABLE_reg : DFFPOSX1 port map( D => n1129, CLK => CLK, Q => R_ENABLE_port
                           );
   DATA_reg_7_inst : DFFPOSX1 port map( D => n1130, CLK => CLK, Q => 
                           DATA_7_port);
   DATA_reg_6_inst : DFFPOSX1 port map( D => n1131, CLK => CLK, Q => 
                           DATA_6_port);
   DATA_reg_5_inst : DFFPOSX1 port map( D => n1132, CLK => CLK, Q => 
                           DATA_5_port);
   DATA_reg_4_inst : DFFPOSX1 port map( D => n1133, CLK => CLK, Q => 
                           DATA_4_port);
   DATA_reg_3_inst : DFFPOSX1 port map( D => n1134, CLK => CLK, Q => 
                           DATA_3_port);
   DATA_reg_2_inst : DFFPOSX1 port map( D => n1135, CLK => CLK, Q => 
                           DATA_2_port);
   DATA_reg_1_inst : DFFPOSX1 port map( D => n1136, CLK => CLK, Q => 
                           DATA_1_port);
   DATA_reg_0_inst : DFFPOSX1 port map( D => n1137, CLK => CLK, Q => 
                           DATA_0_port);
   U3 : NOR2X1 port map( A => n1602, B => n577, Y => n1153);
   U7 : AOI22X1 port map( A => n271, B => extratemp_7_port, C => n604, D => 
                           temp_7_port, Y => n1601);
   U8 : OAI21X1 port map( A => n463, B => n976, C => n1600, Y => n1602);
   U9 : AOI22X1 port map( A => DATA_IN(7), B => n1599, C => 
                           prefillCounter_7_port, D => n275, Y => n1600);
   U10 : NOR2X1 port map( A => n1598, B => n575, Y => n1152);
   U12 : AOI22X1 port map( A => n271, B => extratemp_6_port, C => n604, D => 
                           temp_6_port, Y => n1597);
   U13 : OAI21X1 port map( A => n463, B => n977, C => n1596, Y => n1598);
   U14 : AOI22X1 port map( A => DATA_IN(6), B => n1599, C => 
                           prefillCounter_6_port, D => n275, Y => n1596);
   U15 : NOR2X1 port map( A => n1595, B => n572, Y => n1151);
   U17 : AOI22X1 port map( A => n271, B => extratemp_5_port, C => n604, D => 
                           temp_5_port, Y => n1594);
   U18 : OAI21X1 port map( A => n463, B => n978, C => n1593, Y => n1595);
   U19 : AOI22X1 port map( A => DATA_IN(5), B => n1599, C => 
                           prefillCounter_5_port, D => n275, Y => n1593);
   U20 : NOR2X1 port map( A => n1592, B => n571, Y => n1150);
   U22 : AOI22X1 port map( A => n271, B => extratemp_4_port, C => n604, D => 
                           temp_4_port, Y => n1591);
   U23 : OAI21X1 port map( A => n463, B => n979, C => n1590, Y => n1592);
   U24 : AOI22X1 port map( A => DATA_IN(4), B => n1599, C => 
                           prefillCounter_4_port, D => n275, Y => n1590);
   U25 : NOR2X1 port map( A => n1589, B => n569, Y => n1149);
   U27 : AOI22X1 port map( A => n271, B => extratemp_3_port, C => n604, D => 
                           temp_3_port, Y => n1588);
   U28 : OAI21X1 port map( A => n463, B => n980, C => n1587, Y => n1589);
   U29 : AOI22X1 port map( A => DATA_IN(3), B => n1599, C => 
                           prefillCounter_3_port, D => n275, Y => n1587);
   U30 : NOR2X1 port map( A => n1586, B => n562, Y => n1148);
   U32 : AOI22X1 port map( A => n271, B => extratemp_2_port, C => n604, D => 
                           temp_2_port, Y => n1585);
   U33 : OAI21X1 port map( A => n463, B => n981, C => n1584, Y => n1586);
   U34 : AOI22X1 port map( A => DATA_IN(2), B => n1599, C => 
                           prefillCounter_2_port, D => n275, Y => n1584);
   U35 : NOR2X1 port map( A => n1583, B => n557, Y => n1147);
   U37 : AOI22X1 port map( A => n271, B => extratemp_1_port, C => n604, D => 
                           temp_1_port, Y => n1582);
   U38 : OAI21X1 port map( A => n463, B => n982, C => n1581, Y => n1583);
   U39 : AOI22X1 port map( A => DATA_IN(1), B => n1599, C => 
                           prefillCounter_1_port, D => n275, Y => n1581);
   U40 : NOR2X1 port map( A => n1580, B => n555, Y => n1146);
   U42 : AOI22X1 port map( A => n271, B => extratemp_0_port, C => n604, D => 
                           temp_0_port, Y => n1579);
   U43 : OAI21X1 port map( A => n463, B => n983, C => n1578, Y => n1580);
   U44 : AOI22X1 port map( A => DATA_IN(0), B => n1599, C => 
                           prefillCounter_0_port, D => n275, Y => n1578);
   U46 : NOR2X1 port map( A => n1576, B => n1575, Y => n1145);
   U47 : NAND2X1 port map( A => n1574, B => n1573, Y => n1575);
   U48 : AOI22X1 port map( A => sj_7_port, B => n1572, C => N448, D => n282, Y 
                           => n1573);
   U49 : AOI22X1 port map( A => intj_7_port, B => n280, C => N503, D => n268, Y
                           => n1574);
   U50 : NAND2X1 port map( A => n1570, B => n1569, Y => n1576);
   U51 : AOI22X1 port map( A => temp_7_port, B => n39, C => inti_7_port, D => 
                           n1567, Y => n1569);
   U52 : AOI22X1 port map( A => prefillCounter_7_port, B => n275, C => 
                           faddr_7_port, D => n300, Y => n1570);
   U53 : NOR2X1 port map( A => n1565, B => n1564, Y => n1144);
   U54 : NAND2X1 port map( A => n1563, B => n1562, Y => n1564);
   U55 : AOI22X1 port map( A => sj_6_port, B => n1572, C => N447, D => n282, Y 
                           => n1562);
   U56 : AOI22X1 port map( A => intj_6_port, B => n280, C => N502, D => n268, Y
                           => n1563);
   U57 : NAND2X1 port map( A => n1561, B => n1560, Y => n1565);
   U58 : AOI22X1 port map( A => temp_6_port, B => n39, C => inti_6_port, D => 
                           n1567, Y => n1560);
   U59 : AOI22X1 port map( A => prefillCounter_6_port, B => n275, C => 
                           faddr_6_port, D => n300, Y => n1561);
   U60 : NOR2X1 port map( A => n1559, B => n1558, Y => n1143);
   U61 : NAND2X1 port map( A => n1557, B => n1556, Y => n1558);
   U62 : AOI22X1 port map( A => sj_5_port, B => n1572, C => N446, D => n282, Y 
                           => n1556);
   U63 : AOI22X1 port map( A => intj_5_port, B => n280, C => N501, D => n268, Y
                           => n1557);
   U64 : NAND2X1 port map( A => n1555, B => n1554, Y => n1559);
   U65 : AOI22X1 port map( A => temp_5_port, B => n39, C => inti_5_port, D => 
                           n1567, Y => n1554);
   U66 : AOI22X1 port map( A => prefillCounter_5_port, B => n275, C => 
                           faddr_5_port, D => n300, Y => n1555);
   U67 : NOR2X1 port map( A => n1553, B => n1552, Y => n1142);
   U68 : NAND2X1 port map( A => n1551, B => n1550, Y => n1552);
   U69 : AOI22X1 port map( A => sj_4_port, B => n1572, C => N445, D => n282, Y 
                           => n1550);
   U70 : AOI22X1 port map( A => intj_4_port, B => n280, C => N500, D => n268, Y
                           => n1551);
   U71 : NAND2X1 port map( A => n1549, B => n1548, Y => n1553);
   U72 : AOI22X1 port map( A => temp_4_port, B => n39, C => inti_4_port, D => 
                           n1567, Y => n1548);
   U73 : AOI22X1 port map( A => prefillCounter_4_port, B => n275, C => 
                           faddr_4_port, D => n300, Y => n1549);
   U74 : NOR2X1 port map( A => n1547, B => n1546, Y => n1141);
   U75 : NAND2X1 port map( A => n1545, B => n1544, Y => n1546);
   U76 : AOI22X1 port map( A => sj_3_port, B => n1572, C => N444, D => n282, Y 
                           => n1544);
   U77 : AOI22X1 port map( A => intj_3_port, B => n280, C => N499, D => n268, Y
                           => n1545);
   U78 : NAND2X1 port map( A => n1543, B => n1542, Y => n1547);
   U79 : AOI22X1 port map( A => temp_3_port, B => n39, C => inti_3_port, D => 
                           n1567, Y => n1542);
   U80 : AOI22X1 port map( A => prefillCounter_3_port, B => n275, C => 
                           faddr_3_port, D => n300, Y => n1543);
   U81 : NOR2X1 port map( A => n1541, B => n1540, Y => n1140);
   U82 : NAND2X1 port map( A => n1539, B => n1538, Y => n1540);
   U83 : AOI22X1 port map( A => sj_2_port, B => n1572, C => N443, D => n282, Y 
                           => n1538);
   U84 : AOI22X1 port map( A => intj_2_port, B => n280, C => N498, D => n268, Y
                           => n1539);
   U85 : NAND2X1 port map( A => n1537, B => n1536, Y => n1541);
   U86 : AOI22X1 port map( A => temp_2_port, B => n39, C => inti_2_port, D => 
                           n1567, Y => n1536);
   U87 : AOI22X1 port map( A => prefillCounter_2_port, B => n275, C => 
                           faddr_2_port, D => n300, Y => n1537);
   U88 : NOR2X1 port map( A => n1535, B => n1534, Y => n1139);
   U89 : NAND2X1 port map( A => n1533, B => n1532, Y => n1534);
   U90 : AOI22X1 port map( A => sj_1_port, B => n1572, C => N442, D => n282, Y 
                           => n1532);
   U91 : AOI22X1 port map( A => intj_1_port, B => n280, C => N497, D => n268, Y
                           => n1533);
   U92 : NAND2X1 port map( A => n1531, B => n1530, Y => n1535);
   U93 : AOI22X1 port map( A => temp_1_port, B => n39, C => inti_1_port, D => 
                           n1567, Y => n1530);
   U94 : AOI22X1 port map( A => prefillCounter_1_port, B => n275, C => 
                           faddr_1_port, D => n300, Y => n1531);
   U95 : NOR2X1 port map( A => n1529, B => n1528, Y => n1138);
   U96 : NAND2X1 port map( A => n1527, B => n1526, Y => n1528);
   U97 : AOI22X1 port map( A => sj_0_port, B => n1572, C => n932, D => n282, Y 
                           => n1526);
   U98 : OAI21X1 port map( A => n1525, B => n1524, C => n1523, Y => n1572);
   U99 : AOI22X1 port map( A => intj_0_port, B => n280, C => N496, D => n268, Y
                           => n1527);
   U100 : NAND2X1 port map( A => n1522, B => n1521, Y => n1529);
   U101 : AOI22X1 port map( A => temp_0_port, B => n39, C => inti_0_port, D => 
                           n1567, Y => n1521);
   U102 : OAI21X1 port map( A => n1520, B => n1519, C => n516_port, Y => n1567)
                           ;
   U104 : AOI22X1 port map( A => prefillCounter_0_port, B => n275, C => 
                           faddr_0_port, D => n300, Y => n1522);
   U106 : OAI21X1 port map( A => n252, B => n630, C => n277, Y => n1516);
   U108 : OAI21X1 port map( A => n1515, B => n1514, C => n1513, Y => n1517);
   U109 : AOI21X1 port map( A => n1512, B => n1511, C => n553, Y => n1513);
   U110 : NOR2X1 port map( A => KEY_ERROR, B => n1510, Y => n1512);
   U111 : OAI21X1 port map( A => n373, B => n1509, C => n371, Y => n1514);
   U112 : NAND3X1 port map( A => n1508, B => n1507, C => n1506, Y => 
                           nextState_3_port);
   U113 : AOI21X1 port map( A => n600, B => n629, C => n1505, Y => n1506);
   U114 : NAND2X1 port map( A => n1504, B => n1503, Y => n1505);
   U115 : AOI22X1 port map( A => n1502, B => n371, C => n547, D => n1501, Y => 
                           n1508);
   U116 : NAND3X1 port map( A => n1500, B => n1499, C => n1498, Y => 
                           nextState_2_port);
   U117 : NOR2X1 port map( A => n1497, B => n1496, Y => n1498);
   U118 : OAI21X1 port map( A => n1495, B => n1525, C => n1507, Y => n1496);
   U119 : AOI21X1 port map( A => n1494, B => permuteComplete, C => n1493, Y => 
                           n1507);
   U120 : NAND2X1 port map( A => n249, B => n1492, Y => n1493);
   U121 : OAI22X1 port map( A => n1519, B => n1491, C => KEY_ERROR, D => n1490,
                           Y => n1497);
   U122 : AOI22X1 port map( A => n1489, B => n1488, C => n1487, D => n1486, Y 
                           => n1490);
   U123 : NOR2X1 port map( A => n1485, B => n373, Y => n1489);
   U124 : NOR2X1 port map( A => n271, B => n618, Y => n1499);
   U125 : NOR2X1 port map( A => n616, B => n1484, Y => n1500);
   U126 : NAND3X1 port map( A => n1483, B => n1482, C => n1481, Y => 
                           nextState_1_port);
   U127 : NOR2X1 port map( A => n1480, B => n1479, Y => n1481);
   U128 : OAI21X1 port map( A => n1478, B => n1477, C => n220, Y => n1479);
   U129 : NAND3X1 port map( A => n1475, B => n413_port, C => n1474, Y => n1477)
                           ;
   U130 : NOR2X1 port map( A => prefillCounter_2_port, B => 
                           prefillCounter_1_port, Y => n1474);
   U131 : NAND3X1 port map( A => n1473, B => n922, C => n1472, Y => n1478);
   U132 : NOR2X1 port map( A => prefillCounter_4_port, B => 
                           prefillCounter_3_port, Y => n1472);
   U133 : NOR2X1 port map( A => prefillCounter_7_port, B => 
                           prefillCounter_6_port, Y => n1473);
   U135 : AOI22X1 port map( A => n1471, B => state_0_port, C => n1470, D => 
                           n371, Y => n1483);
   U137 : OAI21X1 port map( A => n542, B => n1486, C => n1469, Y => n1470);
   U138 : NAND2X1 port map( A => n1501, B => n1468, Y => n1469);
   U139 : OAI21X1 port map( A => n1467, B => n1486, C => n1466, Y => n1468);
   U140 : OAI21X1 port map( A => n1485, B => n373, C => n594, Y => n1466);
   U143 : NAND3X1 port map( A => n379, B => n377, C => BYTE_READY, Y => n1486);
   U145 : NOR2X1 port map( A => state_1_port, B => n1519, Y => n1471);
   U146 : NAND3X1 port map( A => n1464, B => n1463, C => n1462, Y => 
                           nextState_0_port);
   U147 : NOR2X1 port map( A => n282, B => n1461, Y => n1462);
   U148 : OAI21X1 port map( A => KEY_ERROR, B => n1460, C => n1482, Y => n1461)
                           ;
   U149 : NOR2X1 port map( A => n1459, B => n1458, Y => n1482);
   U150 : OAI21X1 port map( A => permuteComplete, B => n592, C => n1457, Y => 
                           n1458);
   U151 : NAND3X1 port map( A => n1492, B => n1456, C => n1455, Y => n1459);
   U152 : AOI21X1 port map( A => n1488, B => n1510, C => n1454, Y => n1460);
   U153 : OAI21X1 port map( A => n252, B => n1453, C => n1452, Y => n1454);
   U154 : NAND3X1 port map( A => BYTE_READY, B => n1487, C => n375, Y => n1452)
                           ;
   U156 : NAND2X1 port map( A => OPCODE(0), B => n377, Y => n1509);
   U158 : NAND2X1 port map( A => BYTE_READY, B => n1451, Y => n1510);
   U159 : OAI21X1 port map( A => OPCODE(0), B => OPCODE(1), C => n1465, Y => 
                           n1451);
   U160 : NAND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n1465);
   U161 : NOR2X1 port map( A => n553, B => n271, Y => n1463);
   U162 : NOR2X1 port map( A => n1475, B => n1450, Y => n1464);
   U163 : OAI21X1 port map( A => n318, B => n415, C => n1449, Y => n1137);
   U164 : NAND2X1 port map( A => DATA_0_port, B => n305, Y => n1449);
   U165 : OAI21X1 port map( A => n326, B => n462, C => n1448, Y => n1136);
   U166 : NAND2X1 port map( A => DATA_1_port, B => n327, Y => n1448);
   U167 : OAI21X1 port map( A => n326, B => n459, C => n1447, Y => n1135);
   U168 : NAND2X1 port map( A => DATA_2_port, B => n327, Y => n1447);
   U169 : OAI21X1 port map( A => n326, B => n458, C => n1446, Y => n1134);
   U170 : NAND2X1 port map( A => DATA_3_port, B => n327, Y => n1446);
   U171 : OAI21X1 port map( A => n326, B => n455_port, C => n1445, Y => n1133);
   U172 : NAND2X1 port map( A => DATA_4_port, B => RST, Y => n1445);
   U173 : OAI21X1 port map( A => n326, B => n453_port, C => n1444, Y => n1132);
   U174 : NAND2X1 port map( A => DATA_5_port, B => n327, Y => n1444);
   U175 : OAI21X1 port map( A => n326, B => n451_port, C => n1443, Y => n1131);
   U176 : NAND2X1 port map( A => DATA_6_port, B => n327, Y => n1443);
   U177 : OAI21X1 port map( A => n326, B => n449_port, C => n1442, Y => n1130);
   U178 : NAND2X1 port map( A => DATA_7_port, B => n327, Y => n1442);
   U179 : OAI21X1 port map( A => n326, B => n1441, C => n1440, Y => n1129);
   U180 : NAND2X1 port map( A => R_ENABLE_port, B => n327, Y => n1440);
   U181 : AOI21X1 port map( A => fr_enable, B => n1439, C => n1438, Y => n1441)
                           ;
   U182 : OAI21X1 port map( A => n318, B => n1437, C => n1436, Y => n1128);
   U183 : NAND2X1 port map( A => W_ENABLE_port, B => n326, Y => n1436);
   U184 : AOI21X1 port map( A => fw_enable, B => n1435, C => n1434, Y => n1437)
                           ;
   U185 : OAI21X1 port map( A => n318, B => n518_port, C => n1433, Y => n1127);
   U186 : OAI21X1 port map( A => n318, B => n1439, C => fr_enable, Y => n1433);
   U187 : NAND3X1 port map( A => n1432, B => n1431, C => n1430, Y => n1439);
   U188 : NOR2X1 port map( A => n606, B => n1429, Y => n1430);
   U189 : NAND2X1 port map( A => n247, B => n44, Y => n1429);
   U191 : NAND2X1 port map( A => n610, B => n624, Y => n1523);
   U192 : OAI21X1 port map( A => n318, B => n528, C => n1428, Y => n1126);
   U193 : OAI21X1 port map( A => n318, B => n1435, C => fw_enable, Y => n1428);
   U195 : NAND3X1 port map( A => n247, B => n44, C => n1427, Y => n1434);
   U196 : NOR2X1 port map( A => n1599, B => n604, Y => n1427);
   U197 : OAI22X1 port map( A => n343, B => n983, C => n317, D => n415, Y => 
                           n1125);
   U200 : OAI22X1 port map( A => n343, B => n982, C => n311, D => n462, Y => 
                           n1124);
   U203 : OAI22X1 port map( A => n343, B => n981, C => n317, D => n459, Y => 
                           n1123);
   U206 : OAI22X1 port map( A => n343, B => n980, C => n311, D => n458, Y => 
                           n1122);
   U209 : OAI22X1 port map( A => n345, B => n979, C => n317, D => n455_port, Y 
                           => n1121);
   U212 : OAI22X1 port map( A => n341, B => n978, C => n311, D => n453_port, Y 
                           => n1120);
   U215 : OAI22X1 port map( A => n341, B => n977, C => n317, D => n451_port, Y 
                           => n1119);
   U218 : OAI22X1 port map( A => n341, B => n976, C => n311, D => n449_port, Y 
                           => n1118);
   U221 : OAI21X1 port map( A => n318, B => n417, C => n1426, Y => n1117);
   U222 : NAND2X1 port map( A => ADDR_0_port, B => n326, Y => n1426);
   U223 : OAI22X1 port map( A => n337, B => n975, C => n311, D => n417, Y => 
                           n1116);
   U226 : OAI21X1 port map( A => n318, B => n501_port, C => n1425, Y => n1115);
   U227 : NAND2X1 port map( A => ADDR_1_port, B => n327, Y => n1425);
   U228 : OAI22X1 port map( A => n347, B => n974, C => n311, D => n501_port, Y 
                           => n1114);
   U231 : OAI21X1 port map( A => n318, B => n503_port, C => n1424, Y => n1113);
   U232 : NAND2X1 port map( A => ADDR_2_port, B => n326, Y => n1424);
   U233 : OAI22X1 port map( A => n349, B => n973, C => n311, D => n503_port, Y 
                           => n1112);
   U236 : OAI21X1 port map( A => n318, B => n504, C => n1423, Y => n1111);
   U237 : NAND2X1 port map( A => ADDR_3_port, B => n327, Y => n1423);
   U238 : OAI22X1 port map( A => n339, B => n972, C => n311, D => n504, Y => 
                           n1110);
   U241 : OAI21X1 port map( A => n318, B => n505, C => n1422, Y => n1109);
   U242 : NAND2X1 port map( A => ADDR_4_port, B => n327, Y => n1422);
   U243 : OAI22X1 port map( A => n329, B => n971, C => n311, D => n505, Y => 
                           n1108);
   U246 : OAI21X1 port map( A => n318, B => n506, C => n1421, Y => n1107);
   U247 : NAND2X1 port map( A => ADDR_5_port, B => n327, Y => n1421);
   U248 : OAI22X1 port map( A => n335, B => n970, C => n311, D => n506, Y => 
                           n1106);
   U251 : OAI21X1 port map( A => n317, B => n507, C => n1420, Y => n1105);
   U252 : NAND2X1 port map( A => ADDR_6_port, B => n327, Y => n1420);
   U253 : OAI22X1 port map( A => n333, B => n969, C => n311, D => n507, Y => 
                           n1104);
   U256 : OAI21X1 port map( A => n317, B => n509, C => n1419, Y => n1103);
   U257 : NAND2X1 port map( A => ADDR_7_port, B => n327, Y => n1419);
   U258 : OAI22X1 port map( A => n331, B => n968, C => n311, D => n509, Y => 
                           n1102);
   U261 : OAI21X1 port map( A => n317, B => n381, C => n1418, Y => n1101);
   U262 : NAND2X1 port map( A => PROCESSED_DATA_7_port, B => n327, Y => n1418);
   U264 : OAI21X1 port map( A => n512_port, B => n967, C => n1417, Y => 
                           nextProcessedData_7_port);
   U265 : AOI22X1 port map( A => n37, B => n1415, C => BYTE(7), D => n605, Y =>
                           n1417);
   U266 : XOR2X1 port map( A => temp_7_port, B => delaydata_7_port, Y => n1415)
                           ;
   U268 : OAI21X1 port map( A => n317, B => n385, C => n1414, Y => n1100);
   U269 : NAND2X1 port map( A => PROCESSED_DATA_6_port, B => n327, Y => n1414);
   U271 : OAI21X1 port map( A => n512_port, B => n966, C => n1413, Y => 
                           nextProcessedData_6_port);
   U272 : AOI22X1 port map( A => n37, B => n1412, C => BYTE(6), D => n605, Y =>
                           n1413);
   U273 : XOR2X1 port map( A => temp_6_port, B => delaydata_6_port, Y => n1412)
                           ;
   U275 : OAI21X1 port map( A => n317, B => n389, C => n1411, Y => n1099);
   U276 : NAND2X1 port map( A => PROCESSED_DATA_5_port, B => n327, Y => n1411);
   U278 : OAI21X1 port map( A => n512_port, B => n965, C => n1410, Y => 
                           nextProcessedData_5_port);
   U279 : AOI22X1 port map( A => n37, B => n1409, C => BYTE(5), D => n605, Y =>
                           n1410);
   U280 : XOR2X1 port map( A => temp_5_port, B => delaydata_5_port, Y => n1409)
                           ;
   U282 : OAI21X1 port map( A => n317, B => n393, C => n1408, Y => n1098);
   U283 : NAND2X1 port map( A => PROCESSED_DATA_4_port, B => n327, Y => n1408);
   U285 : OAI21X1 port map( A => n512_port, B => n964, C => n1407, Y => 
                           nextProcessedData_4_port);
   U286 : AOI22X1 port map( A => n37, B => n1406, C => BYTE(4), D => n605, Y =>
                           n1407);
   U287 : XOR2X1 port map( A => temp_4_port, B => delaydata_4_port, Y => n1406)
                           ;
   U289 : OAI21X1 port map( A => n318, B => n397, C => n1405, Y => n1097);
   U290 : NAND2X1 port map( A => PROCESSED_DATA_3_port, B => n327, Y => n1405);
   U292 : OAI21X1 port map( A => n512_port, B => n963, C => n1404, Y => 
                           nextProcessedData_3_port);
   U293 : AOI22X1 port map( A => n37, B => n1403, C => BYTE(3), D => n605, Y =>
                           n1404);
   U294 : XOR2X1 port map( A => temp_3_port, B => delaydata_3_port, Y => n1403)
                           ;
   U296 : OAI21X1 port map( A => n317, B => n401, C => n1402, Y => n1096);
   U297 : NAND2X1 port map( A => PROCESSED_DATA_2_port, B => n327, Y => n1402);
   U299 : OAI21X1 port map( A => n512_port, B => n962, C => n1401, Y => 
                           nextProcessedData_2_port);
   U300 : AOI22X1 port map( A => n37, B => n1400, C => BYTE(2), D => n605, Y =>
                           n1401);
   U301 : XOR2X1 port map( A => temp_2_port, B => delaydata_2_port, Y => n1400)
                           ;
   U303 : OAI21X1 port map( A => n317, B => n405, C => n1399, Y => n1095);
   U304 : NAND2X1 port map( A => PROCESSED_DATA_1_port, B => RST, Y => n1399);
   U306 : OAI21X1 port map( A => n512_port, B => n961, C => n1398, Y => 
                           nextProcessedData_1_port);
   U307 : AOI22X1 port map( A => n37, B => n1397, C => BYTE(1), D => n605, Y =>
                           n1398);
   U308 : XOR2X1 port map( A => temp_1_port, B => delaydata_1_port, Y => n1397)
                           ;
   U310 : OAI21X1 port map( A => n317, B => n409_port, C => n1396, Y => n1094);
   U311 : NAND2X1 port map( A => PROCESSED_DATA_0_port, B => RST, Y => n1396);
   U313 : OAI21X1 port map( A => n512_port, B => n960, C => n1395, Y => 
                           nextProcessedData_0_port);
   U314 : AOI22X1 port map( A => n37, B => n1394, C => BYTE(0), D => n605, Y =>
                           n1395);
   U315 : XOR2X1 port map( A => temp_0_port, B => delaydata_0_port, Y => n1394)
                           ;
   U318 : NAND3X1 port map( A => n285, B => n520_port, C => n1392, Y => n1393);
   U319 : NOR2X1 port map( A => n1391, B => n1390, Y => n1392);
   U322 : AOI22X1 port map( A => BYTE(7), B => n241, C => n302, D => 
                           delaydata_7_port, Y => n1388);
   U324 : AOI22X1 port map( A => BYTE(0), B => n241, C => n302, D => 
                           delaydata_0_port, Y => n1387);
   U326 : AOI22X1 port map( A => BYTE(1), B => n241, C => n302, D => 
                           delaydata_1_port, Y => n1386);
   U328 : AOI22X1 port map( A => BYTE(2), B => n241, C => n302, D => 
                           delaydata_2_port, Y => n1385);
   U330 : AOI22X1 port map( A => BYTE(3), B => n241, C => n302, D => 
                           delaydata_3_port, Y => n1384);
   U332 : AOI22X1 port map( A => BYTE(4), B => n241, C => n302, D => 
                           delaydata_4_port, Y => n1383);
   U334 : AOI22X1 port map( A => BYTE(5), B => n241, C => n302, D => 
                           delaydata_5_port, Y => n1382);
   U336 : AOI22X1 port map( A => BYTE(6), B => n241, C => n302, D => 
                           delaydata_6_port, Y => n1381);
   U339 : OAI21X1 port map( A => n20, B => n637, C => n1379, Y => n1093);
   U340 : NAND2X1 port map( A => KEY(56), B => n7, Y => n1379);
   U342 : OAI21X1 port map( A => n12, B => n638, C => n1378, Y => n1092);
   U343 : NAND2X1 port map( A => KEY(57), B => n15, Y => n1378);
   U345 : OAI21X1 port map( A => n10, B => n648, C => n1377, Y => n1091);
   U346 : NAND2X1 port map( A => KEY(58), B => n16, Y => n1377);
   U348 : OAI21X1 port map( A => n9, B => n649, C => n1376, Y => n1090);
   U349 : NAND2X1 port map( A => KEY(59), B => n20, Y => n1376);
   U351 : OAI21X1 port map( A => n8, B => n650, C => n1375, Y => n1089);
   U352 : NAND2X1 port map( A => KEY(60), B => n17, Y => n1375);
   U354 : OAI21X1 port map( A => n7, B => n651, C => n1374, Y => n1088);
   U355 : NAND2X1 port map( A => KEY(61), B => n10, Y => n1374);
   U357 : OAI21X1 port map( A => n12, B => n692, C => n1373, Y => n1087);
   U358 : NAND2X1 port map( A => KEY(62), B => n14, Y => n1373);
   U360 : OAI21X1 port map( A => n10, B => n701, C => n1372, Y => n1086);
   U361 : NAND2X1 port map( A => KEY(63), B => n12, Y => n1372);
   U363 : OAI21X1 port map( A => n9, B => n746, C => n1371, Y => n1085);
   U364 : NAND2X1 port map( A => KEY(48), B => n14, Y => n1371);
   U366 : OAI21X1 port map( A => n8, B => n748, C => n1370, Y => n1084);
   U367 : NAND2X1 port map( A => KEY(49), B => n15, Y => n1370);
   U369 : OAI21X1 port map( A => n9, B => n750, C => n1369, Y => n1083);
   U370 : NAND2X1 port map( A => KEY(50), B => n12, Y => n1369);
   U372 : OAI21X1 port map( A => n8, B => n752, C => n1368, Y => n1082);
   U373 : NAND2X1 port map( A => KEY(51), B => n20, Y => n1368);
   U375 : OAI21X1 port map( A => n7, B => n754, C => n1367, Y => n1081);
   U376 : NAND2X1 port map( A => KEY(52), B => n24, Y => n1367);
   U378 : OAI21X1 port map( A => n6, B => n756, C => n1366, Y => n1080);
   U379 : NAND2X1 port map( A => KEY(53), B => n16, Y => n1366);
   U381 : OAI21X1 port map( A => n20, B => n758, C => n1365, Y => n1079);
   U382 : NAND2X1 port map( A => KEY(54), B => n29, Y => n1365);
   U384 : OAI21X1 port map( A => n17, B => n760, C => n1364, Y => n1078);
   U385 : NAND2X1 port map( A => KEY(55), B => n9, Y => n1364);
   U387 : OAI21X1 port map( A => n16, B => n761, C => n1363, Y => n1077);
   U388 : NAND2X1 port map( A => KEY(40), B => n22, Y => n1363);
   U390 : OAI21X1 port map( A => n17, B => n762, C => n1362, Y => n1076);
   U391 : NAND2X1 port map( A => KEY(41), B => n27, Y => n1362);
   U393 : OAI21X1 port map( A => n16, B => n763, C => n1361, Y => n1075);
   U394 : NAND2X1 port map( A => KEY(42), B => n12, Y => n1361);
   U396 : OAI21X1 port map( A => n15, B => n764, C => n1360, Y => n1074);
   U397 : NAND2X1 port map( A => KEY(43), B => n6, Y => n1360);
   U399 : OAI21X1 port map( A => n14, B => n765, C => n1359, Y => n1073);
   U400 : NAND2X1 port map( A => KEY(44), B => n14, Y => n1359);
   U402 : OAI21X1 port map( A => n15, B => n766, C => n1358, Y => n1072);
   U403 : NAND2X1 port map( A => KEY(45), B => n15, Y => n1358);
   U405 : OAI21X1 port map( A => n14, B => n767, C => n1357, Y => n1071);
   U406 : NAND2X1 port map( A => KEY(46), B => n10, Y => n1357);
   U408 : OAI21X1 port map( A => n12, B => n768, C => n1356, Y => n1070);
   U409 : NAND2X1 port map( A => KEY(47), B => n17, Y => n1356);
   U411 : OAI21X1 port map( A => n10, B => n769, C => n1355, Y => n1069);
   U412 : NAND2X1 port map( A => KEY(32), B => n9, Y => n1355);
   U414 : OAI21X1 port map( A => n15, B => n770, C => n1354, Y => n1068);
   U415 : NAND2X1 port map( A => KEY(33), B => n10, Y => n1354);
   U417 : OAI21X1 port map( A => n14, B => n771, C => n1353, Y => n1067);
   U418 : NAND2X1 port map( A => KEY(34), B => n27, Y => n1353);
   U420 : OAI21X1 port map( A => n6, B => n772, C => n1352, Y => n1066);
   U421 : NAND2X1 port map( A => KEY(35), B => n6, Y => n1352);
   U423 : OAI21X1 port map( A => n29, B => n773, C => n1351, Y => n1065);
   U424 : NAND2X1 port map( A => KEY(36), B => n16, Y => n1351);
   U426 : OAI21X1 port map( A => n27, B => n774, C => n1350, Y => n1064);
   U427 : NAND2X1 port map( A => KEY(37), B => n8, Y => n1350);
   U429 : OAI21X1 port map( A => n24, B => n775, C => n1349, Y => n1063);
   U430 : NAND2X1 port map( A => KEY(38), B => n6, Y => n1349);
   U432 : OAI21X1 port map( A => n22, B => n776, C => n1348, Y => n1062);
   U433 : NAND2X1 port map( A => KEY(39), B => n9, Y => n1348);
   U435 : OAI21X1 port map( A => n15, B => n777, C => n1347, Y => n1061);
   U436 : NAND2X1 port map( A => KEY(24), B => n6, Y => n1347);
   U437 : OAI21X1 port map( A => n17, B => n778, C => n1346, Y => n1060);
   U438 : NAND2X1 port map( A => KEY(25), B => n7, Y => n1346);
   U439 : OAI21X1 port map( A => n7, B => n779, C => n1345, Y => n1059);
   U440 : NAND2X1 port map( A => KEY(26), B => n29, Y => n1345);
   U441 : OAI21X1 port map( A => n6, B => n780, C => n1344, Y => n1058);
   U442 : NAND2X1 port map( A => KEY(27), B => n8, Y => n1344);
   U443 : OAI21X1 port map( A => n29, B => n781, C => n1343, Y => n1057);
   U444 : NAND2X1 port map( A => KEY(28), B => n7, Y => n1343);
   U445 : OAI21X1 port map( A => n27, B => n782, C => n1342, Y => n1056);
   U446 : NAND2X1 port map( A => KEY(29), B => n29, Y => n1342);
   U447 : OAI21X1 port map( A => n29, B => n783, C => n1341, Y => n1055);
   U448 : NAND2X1 port map( A => KEY(30), B => n7, Y => n1341);
   U449 : OAI21X1 port map( A => n27, B => n784, C => n1340, Y => n1054);
   U450 : NAND2X1 port map( A => KEY(31), B => n8, Y => n1340);
   U451 : OAI21X1 port map( A => n24, B => n785, C => n1339, Y => n1053);
   U452 : NAND2X1 port map( A => KEY(16), B => n24, Y => n1339);
   U453 : OAI21X1 port map( A => n22, B => n786, C => n1338, Y => n1052);
   U454 : NAND2X1 port map( A => KEY(17), B => n16, Y => n1338);
   U455 : OAI21X1 port map( A => n16, B => n787, C => n1337, Y => n1051);
   U456 : NAND2X1 port map( A => KEY(18), B => n22, Y => n1337);
   U457 : OAI21X1 port map( A => n12, B => n788, C => n1336, Y => n1050);
   U458 : NAND2X1 port map( A => KEY(19), B => n27, Y => n1336);
   U459 : OAI21X1 port map( A => n10, B => n789, C => n1335, Y => n1049);
   U460 : NAND2X1 port map( A => KEY(20), B => n24, Y => n1335);
   U461 : OAI21X1 port map( A => n20, B => n790, C => n1334, Y => n1048);
   U462 : NAND2X1 port map( A => KEY(21), B => n20, Y => n1334);
   U463 : OAI21X1 port map( A => n14, B => n791, C => n1333, Y => n1047);
   U464 : NAND2X1 port map( A => KEY(22), B => n29, Y => n1333);
   U465 : OAI21X1 port map( A => n9, B => n864, C => n1332, Y => n1046);
   U466 : NAND2X1 port map( A => KEY(23), B => n27, Y => n1332);
   U467 : OAI21X1 port map( A => n9, B => n865, C => n1331, Y => n1045);
   U468 : NAND2X1 port map( A => KEY(8), B => n6, Y => n1331);
   U469 : OAI21X1 port map( A => n8, B => n866, C => n1330, Y => n1044);
   U470 : NAND2X1 port map( A => KEY(9), B => n12, Y => n1330);
   U471 : OAI21X1 port map( A => n22, B => n867, C => n1329, Y => n1043);
   U472 : NAND2X1 port map( A => KEY(10), B => n20, Y => n1329);
   U473 : OAI21X1 port map( A => n7, B => n868, C => n1328, Y => n1042);
   U474 : NAND2X1 port map( A => KEY(11), B => n14, Y => n1328);
   U475 : OAI21X1 port map( A => n6, B => n869, C => n1327, Y => n1041);
   U476 : NAND2X1 port map( A => KEY(12), B => n15, Y => n1327);
   U477 : OAI21X1 port map( A => n8, B => n870, C => n1326, Y => n1040);
   U478 : NAND2X1 port map( A => KEY(13), B => n24, Y => n1326);
   U479 : OAI21X1 port map( A => n24, B => n871, C => n1325, Y => n1039);
   U480 : NAND2X1 port map( A => KEY(14), B => n22, Y => n1325);
   U481 : OAI21X1 port map( A => n24, B => n883, C => n1324, Y => n1038);
   U482 : NAND2X1 port map( A => KEY(6), B => n10, Y => n1324);
   U483 : OAI21X1 port map( A => n17, B => n884, C => n1323, Y => n1037);
   U484 : NAND2X1 port map( A => KEY(5), B => n17, Y => n1323);
   U485 : OAI21X1 port map( A => n15, B => n885, C => n1322, Y => n1036);
   U486 : NAND2X1 port map( A => KEY(4), B => n8, Y => n1322);
   U487 : OAI21X1 port map( A => n14, B => n886, C => n1321, Y => n1035);
   U488 : NAND2X1 port map( A => KEY(3), B => n9, Y => n1321);
   U489 : OAI21X1 port map( A => n27, B => n887, C => n1320, Y => n1034);
   U490 : NAND2X1 port map( A => KEY(2), B => n7, Y => n1320);
   U491 : OAI21X1 port map( A => n29, B => n888, C => n1319, Y => n1033);
   U492 : NAND2X1 port map( A => KEY(1), B => n22, Y => n1319);
   U493 : OAI21X1 port map( A => n12, B => n889, C => n1318, Y => n1032);
   U494 : NAND2X1 port map( A => KEY(0), B => n20, Y => n1318);
   U495 : OAI21X1 port map( A => n22, B => n890, C => n1317, Y => n1031);
   U496 : NAND2X1 port map( A => KEY(15), B => n17, Y => n1317);
   U497 : OAI21X1 port map( A => n10, B => n916, C => n1316, Y => n1030);
   U498 : NAND2X1 port map( A => KEY(7), B => n16, Y => n1316);
   U499 : NOR2X1 port map( A => n1315, B => n1391, Y => n1380);
   U500 : OAI21X1 port map( A => n500_port, B => n924, C => n1314, Y => n1029);
   U501 : AOI22X1 port map( A => N527, B => n1313, C => n237, D => DATA_IN(7), 
                           Y => n1314);
   U503 : OAI21X1 port map( A => n500_port, B => n931, C => n1312, Y => n1028);
   U504 : AOI22X1 port map( A => N526, B => n1313, C => n237, D => DATA_IN(6), 
                           Y => n1312);
   U506 : OAI21X1 port map( A => n500_port, B => n930, C => n1311, Y => n1027);
   U507 : AOI22X1 port map( A => N525, B => n1313, C => n237, D => DATA_IN(5), 
                           Y => n1311);
   U509 : OAI21X1 port map( A => n500_port, B => n929, C => n1310, Y => n1026);
   U510 : AOI22X1 port map( A => N524, B => n1313, C => n237, D => DATA_IN(4), 
                           Y => n1310);
   U512 : OAI21X1 port map( A => n500_port, B => n928, C => n1309, Y => n1025);
   U513 : AOI22X1 port map( A => N523, B => n1313, C => n237, D => DATA_IN(3), 
                           Y => n1309);
   U515 : OAI21X1 port map( A => n500_port, B => n927, C => n1308, Y => n1024);
   U516 : AOI22X1 port map( A => N522, B => n1313, C => n237, D => DATA_IN(2), 
                           Y => n1308);
   U518 : OAI21X1 port map( A => n500_port, B => n926, C => n1307, Y => n1023);
   U519 : AOI22X1 port map( A => N521, B => n1313, C => n237, D => DATA_IN(1), 
                           Y => n1307);
   U521 : OAI21X1 port map( A => n500_port, B => n925, C => n1306, Y => n1022);
   U522 : AOI22X1 port map( A => N520, B => n1313, C => n237, D => DATA_IN(0), 
                           Y => n1306);
   U527 : NAND3X1 port map( A => n1303, B => n522_port, C => n1302, Y => n1305)
                           ;
   U528 : NOR2X1 port map( A => n1389, B => n300, Y => n1302);
   U529 : NAND2X1 port map( A => n1431, B => n545, Y => n1566);
   U530 : NAND3X1 port map( A => n1301, B => n247, C => n1300, Y => n1389);
   U532 : NOR2X1 port map( A => n326, B => n1475, Y => n1303);
   U534 : AOI22X1 port map( A => n295, B => extratemp_0_port, C => DATA_IN(0), 
                           D => n292, Y => n1298);
   U536 : AOI22X1 port map( A => n295, B => extratemp_1_port, C => DATA_IN(1), 
                           D => n292, Y => n1296);
   U538 : AOI22X1 port map( A => n295, B => extratemp_2_port, C => DATA_IN(2), 
                           D => n292, Y => n1295);
   U540 : AOI22X1 port map( A => n295, B => extratemp_3_port, C => DATA_IN(3), 
                           D => n292, Y => n1294);
   U542 : AOI22X1 port map( A => n295, B => extratemp_4_port, C => DATA_IN(4), 
                           D => n292, Y => n1293);
   U544 : AOI22X1 port map( A => n295, B => extratemp_5_port, C => DATA_IN(5), 
                           D => n292, Y => n1292);
   U546 : AOI22X1 port map( A => n295, B => extratemp_6_port, C => DATA_IN(6), 
                           D => n292, Y => n1291);
   U548 : AOI22X1 port map( A => n295, B => extratemp_7_port, C => DATA_IN(7), 
                           D => n292, Y => n1290);
   U550 : NAND3X1 port map( A => n1504, B => n247, C => n1289, Y => n1297);
   U551 : NOR2X1 port map( A => n1288, B => n1577, Y => n1289);
   U552 : NAND3X1 port map( A => n498_port, B => n545, C => n1432, Y => n1577);
   U553 : NAND2X1 port map( A => n610, B => n1501, Y => n1504);
   U555 : OAI22X1 port map( A => n441, B => n932, C => n1286, D => n959, Y => 
                           n1021);
   U556 : OAI22X1 port map( A => n441, B => n369, C => n1286, D => n259, Y => 
                           n1020);
   U557 : OAI22X1 port map( A => n441, B => n933, C => n1286, D => n953, Y => 
                           n1019);
   U559 : NOR2X1 port map( A => n1285, B => n1391, Y => n1286);
   U560 : OAI21X1 port map( A => n240, B => n938, C => n1284, Y => n1018);
   U561 : NAND2X1 port map( A => N519, B => n1283, Y => n1284);
   U563 : OAI21X1 port map( A => n240, B => n945, C => n1282, Y => n1017);
   U564 : NAND2X1 port map( A => N518, B => n1283, Y => n1282);
   U566 : OAI21X1 port map( A => n240, B => n944, C => n1281, Y => n1016);
   U567 : NAND2X1 port map( A => N517, B => n1283, Y => n1281);
   U569 : OAI21X1 port map( A => n240, B => n943, C => n1280, Y => n1015);
   U570 : NAND2X1 port map( A => N516, B => n1283, Y => n1280);
   U572 : OAI21X1 port map( A => n240, B => n942, C => n1279, Y => n1014);
   U573 : NAND2X1 port map( A => N515, B => n1283, Y => n1279);
   U575 : OAI21X1 port map( A => n240, B => n941, C => n1278, Y => n1013);
   U576 : NAND2X1 port map( A => N514, B => n1283, Y => n1278);
   U578 : OAI21X1 port map( A => n240, B => n940, C => n1277, Y => n1012);
   U579 : NAND2X1 port map( A => N513, B => n1283, Y => n1277);
   U581 : OAI21X1 port map( A => n240, B => n939, C => n1276, Y => n1011);
   U582 : NAND2X1 port map( A => N512, B => n1283, Y => n1276);
   U583 : NOR2X1 port map( A => n1492, B => n1275, Y => n1283);
   U586 : NAND3X1 port map( A => n1274, B => n551, C => n1273, Y => n1275);
   U587 : NOR2X1 port map( A => n326, B => n616, Y => n1273);
   U589 : AOI22X1 port map( A => n290, B => inti_7_port, C => N503, D => n255, 
                           Y => n1272);
   U591 : AOI22X1 port map( A => n290, B => inti_6_port, C => N502, D => n255, 
                           Y => n1269);
   U593 : AOI22X1 port map( A => n290, B => inti_5_port, C => N501, D => n255, 
                           Y => n1268);
   U595 : AOI22X1 port map( A => n290, B => inti_4_port, C => N500, D => n255, 
                           Y => n1267);
   U597 : AOI22X1 port map( A => n290, B => inti_3_port, C => N499, D => n253, 
                           Y => n1266);
   U599 : AOI22X1 port map( A => n290, B => inti_2_port, C => N498, D => n253, 
                           Y => n1265);
   U601 : AOI22X1 port map( A => n290, B => inti_1_port, C => N497, D => n253, 
                           Y => n1264);
   U603 : AOI22X1 port map( A => n290, B => inti_0_port, C => N496, D => n253, 
                           Y => n1263);
   U604 : NOR2X1 port map( A => n290, B => n249, Y => n1270);
   U605 : NAND3X1 port map( A => n581, B => n545, C => n443_port, Y => n1271);
   U606 : OAI21X1 port map( A => n419, B => n256, C => n1262, Y => n1010);
   U607 : NAND2X1 port map( A => N480, B => n616, Y => n1262);
   U609 : OAI21X1 port map( A => n419, B => n952, C => n1261, Y => n1009);
   U610 : NAND2X1 port map( A => N481, B => n616, Y => n1261);
   U612 : OAI21X1 port map( A => n419, B => n951, C => n1260, Y => n1008);
   U613 : NAND2X1 port map( A => N482, B => n616, Y => n1260);
   U615 : OAI21X1 port map( A => n419, B => n950, C => n1259, Y => n1007);
   U616 : NAND2X1 port map( A => N483, B => n616, Y => n1259);
   U618 : OAI21X1 port map( A => n419, B => n949, C => n1258, Y => n1006);
   U619 : NAND2X1 port map( A => N484, B => n616, Y => n1258);
   U621 : OAI21X1 port map( A => n419, B => n948, C => n1257, Y => n1005);
   U622 : NAND2X1 port map( A => N485, B => n616, Y => n1257);
   U624 : OAI21X1 port map( A => n419, B => n947, C => n1256, Y => n1004);
   U625 : NAND2X1 port map( A => N486, B => n616, Y => n1256);
   U628 : NAND2X1 port map( A => N487, B => n616, Y => n1255);
   U631 : NAND3X1 port map( A => n551, B => n1492, C => n1274, Y => n1254);
   U632 : NOR2X1 port map( A => n1253, B => n1252, Y => n1274);
   U633 : NAND3X1 port map( A => n1432, B => n581, C => n447_port, Y => n1252);
   U634 : NAND3X1 port map( A => n612, B => n545, C => n1251, Y => n1253);
   U637 : OAI21X1 port map( A => n581, B => n1249, C => n1248, Y => n1002);
   U638 : OAI21X1 port map( A => n1247, B => n1285, C => permuteComplete, Y => 
                           n1248);
   U639 : NAND2X1 port map( A => n1246, B => n439, Y => n1249);
   U641 : NAND3X1 port map( A => n543, B => n249, C => n443_port, Y => n1285);
   U643 : NAND3X1 port map( A => n285, B => n341, C => n447_port, Y => n1245);
   U646 : OAI21X1 port map( A => n445_port, B => n937, C => n1244, Y => n1001);
   U647 : NAND2X1 port map( A => N431, B => n1243, Y => n1244);
   U649 : OAI21X1 port map( A => n445_port, B => n936, C => n1242, Y => n1000);
   U650 : NAND2X1 port map( A => N430, B => n1243, Y => n1242);
   U652 : OAI21X1 port map( A => n445_port, B => n935, C => n1241, Y => n999);
   U653 : NAND2X1 port map( A => N429, B => n1243, Y => n1241);
   U654 : OAI21X1 port map( A => n445_port, B => n934, C => n1240, Y => n998);
   U655 : NAND2X1 port map( A => N428, B => n1243, Y => n1240);
   U656 : OAI21X1 port map( A => n445_port, B => n367, C => n1239, Y => n997);
   U657 : NAND2X1 port map( A => N427, B => n1243, Y => n1239);
   U659 : OAI21X1 port map( A => n445_port, B => n933, C => n1238, Y => n996);
   U660 : NAND2X1 port map( A => N426, B => n1243, Y => n1238);
   U662 : OAI21X1 port map( A => n445_port, B => n369, C => n1237, Y => n995);
   U663 : NAND2X1 port map( A => N425, B => n1243, Y => n1237);
   U664 : OAI21X1 port map( A => n445_port, B => n932, C => n1236, Y => n994);
   U665 : NAND2X1 port map( A => N424, B => n1243, Y => n1236);
   U666 : NOR2X1 port map( A => n581, B => n1246, Y => n1243);
   U667 : NOR2X1 port map( A => n1235, B => n1234, Y => n1246);
   U668 : NAND3X1 port map( A => si_7_port, B => si_6_port, C => n1233, Y => 
                           n1234);
   U669 : NOR2X1 port map( A => n934, B => n935, Y => n1233);
   U672 : NAND3X1 port map( A => si_3_port, B => si_2_port, C => n1232, Y => 
                           n1235);
   U673 : NOR2X1 port map( A => n932, B => n369, Y => n1232);
   U677 : NAND3X1 port map( A => n447_port, B => n285, C => n1230, Y => n1231);
   U678 : NOR2X1 port map( A => n268, B => n1391, Y => n1230);
   U679 : NOR2X1 port map( A => n1453, B => n1519, Y => n1391);
   U681 : OAI21X1 port map( A => n252, B => n1287, C => n549, Y => n1229);
   U684 : NAND3X1 port map( A => n1515, B => n1300, C => n1226, Y => n1227);
   U685 : NOR2X1 port map( A => n1225, B => n1224, Y => n1226);
   U686 : OAI21X1 port map( A => n252, B => n220, C => n1503, Y => n1224);
   U690 : OAI21X1 port map( A => n1524, B => n34, C => n44, Y => n1571);
   U693 : OAI21X1 port map( A => n488, B => n923, C => n1220, Y => n993);
   U694 : NAND2X1 port map( A => N413, B => n1219, Y => n1220);
   U696 : OAI21X1 port map( A => n488, B => n922, C => n1218, Y => n992);
   U697 : NAND2X1 port map( A => N412, B => n1219, Y => n1218);
   U699 : OAI21X1 port map( A => n488, B => n921, C => n1217, Y => n991);
   U700 : NAND2X1 port map( A => N411, B => n1219, Y => n1217);
   U702 : OAI21X1 port map( A => n488, B => n920, C => n1216, Y => n990);
   U703 : NAND2X1 port map( A => N410, B => n1219, Y => n1216);
   U705 : OAI21X1 port map( A => n488, B => n919, C => n1215, Y => n989);
   U706 : NAND2X1 port map( A => N409, B => n1219, Y => n1215);
   U708 : OAI21X1 port map( A => n488, B => n918, C => n1214, Y => n988);
   U709 : NAND2X1 port map( A => N408, B => n1219, Y => n1214);
   U711 : OAI21X1 port map( A => n488, B => n917, C => n1213, Y => n987);
   U712 : NAND2X1 port map( A => N414, B => n1219, Y => n1213);
   U714 : OAI21X1 port map( A => n488, B => n413_port, C => n1212, Y => n986);
   U715 : NAND2X1 port map( A => N407, B => n1219, Y => n1212);
   U716 : NOR2X1 port map( A => n1315, B => n247, Y => n1219);
   U721 : NAND3X1 port map( A => n498_port, B => n1457, C => n1211, Y => n1315)
                           ;
   U722 : NOR2X1 port map( A => n216, B => n1288, Y => n1211);
   U723 : NAND3X1 port map( A => n270, B => n612, C => n1210, Y => n1288);
   U724 : NOR2X1 port map( A => n326, B => n271, Y => n1210);
   U727 : NOR2X1 port map( A => n1519, B => n1287, Y => n1475);
   U732 : NOR2X1 port map( A => n1467, B => n1525, Y => n1484);
   U733 : OAI21X1 port map( A => n1519, B => n1208, C => n524_port, Y => n1299)
                           ;
   U735 : OAI21X1 port map( A => n1476, B => n626, C => n592, Y => n1207);
   U737 : NOR2X1 port map( A => n1524, B => n626, Y => n1494);
   U738 : NAND3X1 port map( A => n1206, B => n624, C => n614, Y => n1457);
   U739 : XOR2X1 port map( A => n42, B => n252, Y => n1206);
   U741 : NAND3X1 port map( A => n1304, B => n1431, C => n518_port, Y => n1435)
                           ;
   U743 : NAND2X1 port map( A => n1301, B => n540, Y => n1438);
   U745 : OAI21X1 port map( A => n1524, B => n34, C => n1223, Y => n1205);
   U746 : NAND2X1 port map( A => n629, B => n541, Y => n1223);
   U748 : NOR2X1 port map( A => n1225, B => n268, Y => n1301);
   U750 : OAI21X1 port map( A => n1525, B => n1524, C => n1204, Y => n1225);
   U751 : NOR2X1 port map( A => n618, B => n1518, Y => n1204);
   U752 : NOR2X1 port map( A => n1467, B => n1519, Y => n1518);
   U754 : NAND2X1 port map( A => n39, B => n42, Y => n1456);
   U755 : NOR2X1 port map( A => n1390, B => n553, Y => n1431);
   U757 : NOR2X1 port map( A => n37, B => n605, Y => n1503);
   U759 : NAND3X1 port map( A => n1501, B => n614, C => n42, Y => n1203);
   U760 : NOR2X1 port map( A => n1209, B => n626, Y => n1416);
   U762 : OAI21X1 port map( A => n220, B => n1525, C => n581, Y => n1202);
   U764 : NOR2X1 port map( A => n1524, B => n1519, Y => n1247);
   U765 : NAND2X1 port map( A => n600, B => n630, Y => n1524);
   U766 : NAND2X1 port map( A => state_0_port, B => n547, Y => n1476);
   U767 : NAND2X1 port map( A => n542, B => n514_port, Y => n1502);
   U769 : AOI21X1 port map( A => n1467, B => n1208, C => n626, Y => n1488);
   U771 : NOR2X1 port map( A => n636, B => state_2_port, Y => n1501);
   U772 : NAND3X1 port map( A => n42, B => n579, C => state_0_port, Y => n1467)
                           ;
   U774 : NAND2X1 port map( A => n543, B => n1221, Y => n1487);
   U778 : NAND2X1 port map( A => n547, B => n632, Y => n1453);
   U780 : NAND2X1 port map( A => n579, B => n630, Y => n1495);
   U781 : NOR2X1 port map( A => n1228, B => n616, Y => n1304);
   U783 : NAND2X1 port map( A => n39, B => n630, Y => n1455);
   U784 : NOR2X1 port map( A => n1525, B => n1520, Y => n1568);
   U785 : NAND3X1 port map( A => n1492, B => n1250, C => n551, Y => n1228);
   U787 : NOR2X1 port map( A => n1519, B => n1209, Y => n1450);
   U788 : NAND3X1 port map( A => n632, B => n579, C => n42, Y => n1209);
   U790 : NAND2X1 port map( A => n624, B => n636, Y => n1519);
   U792 : NAND2X1 port map( A => n594, B => n629, Y => n1250);
   U794 : NAND2X1 port map( A => state_2_port, B => n636, Y => n1525);
   U797 : NAND2X1 port map( A => n600, B => n42, Y => n1208);
   U799 : NAND2X1 port map( A => state_0_port, B => state_1_port, Y => n1491);
   U801 : NAND2X1 port map( A => n614, B => n630, Y => n1287);
   U804 : NAND2X1 port map( A => state_1_port, B => n632, Y => n1520);
   U806 : NAND2X1 port map( A => state_2_port, B => n252, Y => n1222);
   U807 : NAND3X1 port map( A => n1199, B => n1201, C => n1200, Y => N479);
   U808 : NOR2X1 port map( A => n1198, B => n1197, Y => n1199);
   U809 : OAI22X1 port map( A => n865, B => n1196, C => n889, D => n250, Y => 
                           n1197);
   U812 : OAI22X1 port map( A => n777, B => n1194, C => n785, D => n1193, Y => 
                           n1198);
   U815 : AOI22X1 port map( A => n955, B => keyTable_5_0_port, C => n954, D => 
                           keyTable_4_0_port, Y => n1200);
   U816 : AOI22X1 port map( A => n957, B => keyTable_7_0_port, C => 
                           keyTable_6_0_port, D => n956, Y => n1201);
   U817 : NAND3X1 port map( A => n1192, B => n1191, C => n1190, Y => N478);
   U818 : NOR2X1 port map( A => n1189, B => n1188, Y => n1190);
   U819 : OAI22X1 port map( A => n866, B => n1196, C => n888, D => n250, Y => 
                           n1188);
   U822 : OAI22X1 port map( A => n778, B => n1194, C => n786, D => n1193, Y => 
                           n1189);
   U825 : AOI22X1 port map( A => n955, B => keyTable_5_1_port, C => n954, D => 
                           keyTable_4_1_port, Y => n1191);
   U826 : AOI22X1 port map( A => n957, B => keyTable_7_1_port, C => n956, D => 
                           keyTable_6_1_port, Y => n1192);
   U827 : NAND3X1 port map( A => n1187, B => n1186, C => n1185, Y => N477);
   U828 : NOR2X1 port map( A => n1184, B => n1183, Y => n1185);
   U829 : OAI22X1 port map( A => n867, B => n1196, C => n887, D => n250, Y => 
                           n1183);
   U832 : OAI22X1 port map( A => n779, B => n1194, C => n787, D => n264, Y => 
                           n1184);
   U835 : AOI22X1 port map( A => n955, B => keyTable_5_2_port, C => n954, D => 
                           keyTable_4_2_port, Y => n1186);
   U836 : AOI22X1 port map( A => n957, B => keyTable_7_2_port, C => n956, D => 
                           keyTable_6_2_port, Y => n1187);
   U837 : NAND3X1 port map( A => n1182, B => n1181, C => n1180, Y => N476);
   U838 : NOR2X1 port map( A => n1179, B => n1178, Y => n1180);
   U839 : OAI22X1 port map( A => n868, B => n1196, C => n886, D => n250, Y => 
                           n1178);
   U842 : OAI22X1 port map( A => n780, B => n1194, C => n788, D => n264, Y => 
                           n1179);
   U845 : AOI22X1 port map( A => n955, B => keyTable_5_3_port, C => n954, D => 
                           keyTable_4_3_port, Y => n1181);
   U846 : AOI22X1 port map( A => n957, B => keyTable_7_3_port, C => n956, D => 
                           keyTable_6_3_port, Y => n1182);
   U847 : NAND3X1 port map( A => n1177, B => n1176, C => n1175, Y => N475);
   U848 : NOR2X1 port map( A => n1174, B => n1173, Y => n1175);
   U849 : OAI22X1 port map( A => n869, B => n1196, C => n885, D => n250, Y => 
                           n1173);
   U852 : OAI22X1 port map( A => n781, B => n1194, C => n789, D => n264, Y => 
                           n1174);
   U855 : AOI22X1 port map( A => n955, B => keyTable_5_4_port, C => n954, D => 
                           keyTable_4_4_port, Y => n1176);
   U856 : AOI22X1 port map( A => n957, B => keyTable_7_4_port, C => n956, D => 
                           keyTable_6_4_port, Y => n1177);
   U857 : NAND3X1 port map( A => n1172, B => n1171, C => n1170, Y => N474);
   U858 : NOR2X1 port map( A => n1169, B => n1168, Y => n1170);
   U859 : OAI22X1 port map( A => n870, B => n1196, C => n884, D => n250, Y => 
                           n1168);
   U862 : OAI22X1 port map( A => n782, B => n1194, C => n790, D => n264, Y => 
                           n1169);
   U865 : AOI22X1 port map( A => n955, B => keyTable_5_5_port, C => n954, D => 
                           keyTable_4_5_port, Y => n1171);
   U866 : AOI22X1 port map( A => n957, B => keyTable_7_5_port, C => n956, D => 
                           keyTable_6_5_port, Y => n1172);
   U867 : NAND3X1 port map( A => n1167, B => n1166, C => n1165, Y => N473);
   U868 : NOR2X1 port map( A => n1164, B => n1163, Y => n1165);
   U869 : OAI22X1 port map( A => n871, B => n1196, C => n883, D => n250, Y => 
                           n1163);
   U872 : OAI22X1 port map( A => n783, B => n1194, C => n791, D => n264, Y => 
                           n1164);
   U875 : AOI22X1 port map( A => n955, B => keyTable_5_6_port, C => n954, D => 
                           keyTable_4_6_port, Y => n1166);
   U876 : AOI22X1 port map( A => n957, B => keyTable_7_6_port, C => n956, D => 
                           keyTable_6_6_port, Y => n1167);
   U877 : NAND3X1 port map( A => n1162, B => n1161, C => n1160, Y => N472);
   U878 : NOR2X1 port map( A => n1159, B => n1158, Y => n1160);
   U879 : OAI22X1 port map( A => n890, B => n1196, C => n916, D => n250, Y => 
                           n1158);
   U880 : NAND3X1 port map( A => n953, B => n958, C => n959, Y => n1195);
   U882 : NAND3X1 port map( A => n958, B => keyi_0_port, C => n953, Y => n1196)
                           ;
   U884 : OAI22X1 port map( A => n784, B => n1194, C => n864, D => n264, Y => 
                           n1159);
   U885 : NAND3X1 port map( A => n959, B => n953, C => n265, Y => n1193);
   U887 : NAND3X1 port map( A => keyi_1_port, B => keyi_0_port, C => n953, Y =>
                           n1194);
   U890 : AOI22X1 port map( A => n955, B => keyTable_5_7_port, C => n954, D => 
                           keyTable_4_7_port, Y => n1161);
   U892 : NAND3X1 port map( A => n959, B => n259, C => n261, Y => n1157);
   U894 : NAND3X1 port map( A => n259, B => n258, C => n261, Y => n1156);
   U896 : AOI22X1 port map( A => n957, B => keyTable_7_7_port, C => n956, D => 
                           keyTable_6_7_port, Y => n1162);
   U898 : NAND3X1 port map( A => keyi_1_port, B => n959, C => n261, Y => n1155)
                           ;
   U901 : NAND3X1 port map( A => n265, B => n258, C => n261, Y => n1154);
   U105 : OR2X2 port map( A => n1517, B => n1516, Y => nextState_4_port);
   U134 : OR2X2 port map( A => n1484, B => n605, Y => n1480);
   U142 : AND2X2 port map( A => n1509, B => n1465, Y => n1485);
   U524 : AND2X2 port map( A => n1484, B => n500_port, Y => n1313);
   U635 : AND2X2 port map( A => n249, B => n1250, Y => n1251);
   U692 : AND2X2 port map( A => n1221, B => n514_port, Y => n1515);
   U761 : OR2X2 port map( A => n1502, B => n1202, Y => n1390);
   U775 : OR2X2 port map( A => n34, B => n1209, Y => n1221);
   U800 : OR2X2 port map( A => n34, B => n1287, Y => n1492);
   add_377 : KSA_0_DW01_add_0 port map( A(7) => temp_7_port, A(6) => 
                           temp_6_port, A(5) => temp_5_port, A(4) => 
                           temp_4_port, A(3) => temp_3_port, A(2) => 
                           temp_2_port, A(1) => temp_1_port, A(0) => 
                           temp_0_port, B(7) => extratemp_7_port, B(6) => 
                           extratemp_6_port, B(5) => extratemp_5_port, B(4) => 
                           extratemp_4_port, B(3) => extratemp_3_port, B(2) => 
                           extratemp_2_port, B(1) => extratemp_1_port, B(0) => 
                           extratemp_0_port, CI => n1604, SUM(7) => N527, 
                           SUM(6) => N526, SUM(5) => N525, SUM(4) => N524, 
                           SUM(3) => N523, SUM(2) => N522, SUM(1) => N521, 
                           SUM(0) => N520, CO => n_1021);
   add_337 : KSA_0_DW01_add_1 port map( A(7) => intj_7_port, A(6) => 
                           intj_6_port, A(5) => intj_5_port, A(4) => 
                           intj_4_port, A(3) => intj_3_port, A(2) => 
                           intj_2_port, A(1) => intj_1_port, A(0) => 
                           intj_0_port, B(7) => DATA_IN(7), B(6) => DATA_IN(6),
                           B(5) => DATA_IN(5), B(4) => DATA_IN(4), B(3) => 
                           DATA_IN(3), B(2) => DATA_IN(2), B(1) => DATA_IN(1), 
                           B(0) => DATA_IN(0), CI => n1603, SUM(7) => N519, 
                           SUM(6) => N518, SUM(5) => N517, SUM(4) => N516, 
                           SUM(3) => N515, SUM(2) => N514, SUM(1) => N513, 
                           SUM(0) => N512, CO => n_1022);
   add_289 : KSA_0_DW01_inc_0 port map( A(7) => si_7_port, A(6) => si_6_port, 
                           A(5) => si_5_port, A(4) => si_4_port, A(3) => 
                           si_3_port, A(2) => si_2_port, A(1) => si_1_port, 
                           A(0) => si_0_port, SUM(7) => N431, SUM(6) => N430, 
                           SUM(5) => N429, SUM(4) => N428, SUM(3) => N427, 
                           SUM(2) => N426, SUM(1) => N425, SUM(0) => N424);
   add_263 : KSA_0_DW01_inc_1 port map( A(7) => prefillCounter_7_port, A(6) => 
                           prefillCounter_6_port, A(5) => prefillCounter_5_port
                           , A(4) => prefillCounter_4_port, A(3) => 
                           prefillCounter_3_port, A(2) => prefillCounter_2_port
                           , A(1) => prefillCounter_1_port, A(0) => 
                           prefillCounter_0_port, SUM(7) => N414, SUM(6) => 
                           N413, SUM(5) => N412, SUM(4) => N411, SUM(3) => N410
                           , SUM(2) => N409, SUM(1) => N408, SUM(0) => N407);
   r126 : KSA_0_DW01_inc_2 port map( A(7) => inti_7_port, A(6) => inti_6_port, 
                           A(5) => inti_5_port, A(4) => inti_4_port, A(3) => 
                           inti_3_port, A(2) => inti_2_port, A(1) => 
                           inti_1_port, A(0) => inti_0_port, SUM(7) => N503, 
                           SUM(6) => N502, SUM(5) => N501, SUM(4) => N500, 
                           SUM(3) => N499, SUM(2) => N498, SUM(1) => N497, 
                           SUM(0) => N496);
   add_1_root_add_0_root_add_302_2 : KSA_0_DW01_add_3 port map( A(7) => 
                           DATA_IN(7), A(6) => DATA_IN(6), A(5) => DATA_IN(5), 
                           A(4) => DATA_IN(4), A(3) => DATA_IN(3), A(2) => 
                           DATA_IN(2), A(1) => DATA_IN(1), A(0) => DATA_IN(0), 
                           B(7) => sj_7_port, B(6) => sj_6_port, B(5) => 
                           sj_5_port, B(4) => sj_4_port, B(3) => sj_3_port, 
                           B(2) => sj_2_port, B(1) => sj_1_port, B(0) => 
                           sj_0_port, CI => n984, SUM(7) => N456, SUM(6) => 
                           N455, SUM(5) => N454, SUM(4) => N453, SUM(3) => N452
                           , SUM(2) => N451, SUM(1) => N450, SUM(0) => N449, CO
                           => n_1023);
   add_0_root_add_0_root_add_302_2 : KSA_0_DW01_add_2 port map( A(7) => N472, 
                           A(6) => N473, A(5) => N474, A(4) => N475, A(3) => 
                           N476, A(2) => N477, A(1) => N478, A(0) => N479, B(7)
                           => N456, B(6) => N455, B(5) => N454, B(4) => N453, 
                           B(3) => N452, B(2) => N451, B(1) => N450, B(0) => 
                           N449, CI => n985, SUM(7) => N487, SUM(6) => N486, 
                           SUM(5) => N485, SUM(4) => N484, SUM(3) => N483, 
                           SUM(2) => N482, SUM(1) => N481, SUM(0) => N480, CO 
                           => n_1024);
   nfaddr_tri_5_inst : TBUFX1 port map( A => n1143, EN => n285, Y => 
                           nfaddr_5_port);
   nfaddr_tri_0_inst : TBUFX1 port map( A => n1138, EN => n285, Y => 
                           nfaddr_0_port);
   nfaddr_tri_1_inst : TBUFX1 port map( A => n1139, EN => n285, Y => 
                           nfaddr_1_port);
   nfaddr_tri_2_inst : TBUFX1 port map( A => n1140, EN => n285, Y => 
                           nfaddr_2_port);
   nfaddr_tri_3_inst : TBUFX1 port map( A => n1141, EN => n285, Y => 
                           nfaddr_3_port);
   nfaddr_tri_4_inst : TBUFX1 port map( A => n1142, EN => n285, Y => 
                           nfaddr_4_port);
   nfaddr_tri_6_inst : TBUFX1 port map( A => n1144, EN => n285, Y => 
                           nfaddr_6_port);
   nfaddr_tri_7_inst : TBUFX1 port map( A => n1145, EN => n285, Y => 
                           nfaddr_7_port);
   nfdata_tri_0_inst : TBUFX1 port map( A => n1146, EN => n612, Y => 
                           nfdata_0_port);
   nfdata_tri_1_inst : TBUFX1 port map( A => n1147, EN => n612, Y => 
                           nfdata_1_port);
   nfdata_tri_2_inst : TBUFX1 port map( A => n1148, EN => n612, Y => 
                           nfdata_2_port);
   nfdata_tri_3_inst : TBUFX1 port map( A => n1149, EN => n612, Y => 
                           nfdata_3_port);
   nfdata_tri_4_inst : TBUFX1 port map( A => n1150, EN => n612, Y => 
                           nfdata_4_port);
   nfdata_tri_5_inst : TBUFX1 port map( A => n1151, EN => n612, Y => 
                           nfdata_5_port);
   nfdata_tri_6_inst : TBUFX1 port map( A => n1152, EN => n612, Y => 
                           nfdata_6_port);
   nfdata_tri_7_inst : TBUFX1 port map( A => n1153, EN => n612, Y => 
                           nfdata_7_port);
   PDATA_READY_reg : DFFSR port map( D => n553, CLK => CLK, R => n307, S => 
                           n214, Q => PDATA_READY);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n307, S => n212, Q => state_1_port);
   state_reg_3_inst : DFFSR port map( D => nextState_3_port, CLK => CLK, R => 
                           n307, S => n210, Q => state_3_port);
   state_reg_4_inst : DFFSR port map( D => nextState_4_port, CLK => CLK, R => 
                           n307, S => n208, Q => state_4_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n307, S => n206, Q => state_2_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n307, S => n203, Q => state_0_port);
   si_reg_7_inst : DFFSR port map( D => n1001, CLK => CLK, R => n307, S => n196
                           , Q => si_7_port);
   si_reg_6_inst : DFFSR port map( D => n1000, CLK => CLK, R => n307, S => n188
                           , Q => si_6_port);
   si_reg_5_inst : DFFSR port map( D => n999, CLK => CLK, R => n307, S => n187,
                           Q => si_5_port);
   si_reg_4_inst : DFFSR port map( D => n998, CLK => CLK, R => n307, S => n185,
                           Q => si_4_port);
   si_reg_3_inst : DFFSR port map( D => n997, CLK => CLK, R => n307, S => n180,
                           Q => si_3_port);
   si_reg_2_inst : DFFSR port map( D => n996, CLK => CLK, R => n307, S => n177,
                           Q => si_2_port);
   si_reg_1_inst : DFFSR port map( D => n995, CLK => CLK, R => n307, S => n175,
                           Q => si_1_port);
   si_reg_0_inst : DFFSR port map( D => n994, CLK => CLK, R => n307, S => n172,
                           Q => si_0_port);
   currentProcessedData_reg_7_inst : DFFSR port map( D => 
                           nextProcessedData_7_port, CLK => CLK, R => n307, S 
                           => n161, Q => currentProcessedData_7_port);
   currentProcessedData_reg_6_inst : DFFSR port map( D => 
                           nextProcessedData_6_port, CLK => CLK, R => n307, S 
                           => n160, Q => currentProcessedData_6_port);
   currentProcessedData_reg_5_inst : DFFSR port map( D => 
                           nextProcessedData_5_port, CLK => CLK, R => n307, S 
                           => n151, Q => currentProcessedData_5_port);
   currentProcessedData_reg_4_inst : DFFSR port map( D => 
                           nextProcessedData_4_port, CLK => CLK, R => n307, S 
                           => n141, Q => currentProcessedData_4_port);
   currentProcessedData_reg_3_inst : DFFSR port map( D => 
                           nextProcessedData_3_port, CLK => CLK, R => n307, S 
                           => n136, Q => currentProcessedData_3_port);
   currentProcessedData_reg_2_inst : DFFSR port map( D => 
                           nextProcessedData_2_port, CLK => CLK, R => n307, S 
                           => n135, Q => currentProcessedData_2_port);
   currentProcessedData_reg_1_inst : DFFSR port map( D => 
                           nextProcessedData_1_port, CLK => CLK, R => n307, S 
                           => n131, Q => currentProcessedData_1_port);
   currentProcessedData_reg_0_inst : DFFSR port map( D => 
                           nextProcessedData_0_port, CLK => CLK, R => n307, S 
                           => n129, Q => currentProcessedData_0_port);
   sj_reg_5_inst : DFFSR port map( D => n1005, CLK => CLK, R => n307, S => n122
                           , Q => sj_5_port);
   sj_reg_4_inst : DFFSR port map( D => n1006, CLK => CLK, R => n307, S => n121
                           , Q => sj_4_port);
   sj_reg_3_inst : DFFSR port map( D => n1007, CLK => CLK, R => n307, S => n117
                           , Q => sj_3_port);
   sj_reg_2_inst : DFFSR port map( D => n1008, CLK => CLK, R => n307, S => n64,
                           Q => sj_2_port);
   sj_reg_1_inst : DFFSR port map( D => n1009, CLK => CLK, R => n307, S => n62,
                           Q => sj_1_port);
   sj_reg_0_inst : DFFSR port map( D => n1010, CLK => CLK, R => n307, S => n54,
                           Q => sj_0_port);
   sj_reg_6_inst : DFFSR port map( D => n1004, CLK => CLK, R => n307, S => n52,
                           Q => sj_6_port);
   sj_reg_7_inst : DFFSR port map( D => n1003, CLK => CLK, R => n307, S => n49,
                           Q => sj_7_port);
   U4 : BUFX4 port map( A => n1195, Y => n250);
   U11 : INVX4 port map( A => n1157, Y => n954);
   U16 : BUFX2 port map( A => n1380, Y => n3);
   U21 : BUFX2 port map( A => n1380, Y => n4);
   U26 : BUFX2 port map( A => n1380, Y => n5);
   U31 : BUFX2 port map( A => n3, Y => n6);
   U36 : BUFX2 port map( A => n3, Y => n7);
   U41 : BUFX2 port map( A => n3, Y => n8);
   U45 : BUFX2 port map( A => n3, Y => n9);
   U103 : BUFX2 port map( A => n3, Y => n10);
   U107 : BUFX2 port map( A => n4, Y => n12);
   U136 : BUFX2 port map( A => n4, Y => n14);
   U141 : BUFX2 port map( A => n4, Y => n15);
   U144 : BUFX2 port map( A => n4, Y => n16);
   U155 : BUFX2 port map( A => n4, Y => n17);
   U157 : BUFX2 port map( A => n5, Y => n20);
   U190 : BUFX2 port map( A => n5, Y => n22);
   U194 : BUFX2 port map( A => n5, Y => n24);
   U198 : BUFX2 port map( A => n5, Y => n27);
   U199 : BUFX2 port map( A => n5, Y => n29);
   U201 : INVX4 port map( A => n297, Y => n300);
   U202 : INVX2 port map( A => n1222, Y => n32);
   U204 : INVX4 port map( A => n32, Y => n34);
   U205 : BUFX2 port map( A => n1416, Y => n37);
   U207 : BUFX4 port map( A => state_3_port, Y => n252);
   U208 : INVX2 port map( A => n1155, Y => n956);
   U210 : BUFX2 port map( A => state_4_port, Y => n42);
   U211 : INVX2 port map( A => n287, Y => n290);
   U213 : INVX2 port map( A => n241, Y => n302);
   U214 : INVX2 port map( A => n1305, Y => n500_port);
   U216 : INVX4 port map( A => n1156, Y => n955);
   U217 : BUFX4 port map( A => n1568, Y => n39);
   U219 : INVX2 port map( A => n44, Y => n271);
   U220 : INVX1 port map( A => sj_0_port, Y => n256);
   U224 : INVX2 port map( A => keyi_0_port, Y => n959);
   U225 : INVX1 port map( A => keyi_1_port, Y => n259);
   U229 : OR2X2 port map( A => n1525, B => n1209, Y => n44);
   U230 : INVX2 port map( A => n292, Y => n295);
   U234 : INVX2 port map( A => n249, Y => n268);
   U235 : OR2X2 port map( A => n34, B => n1476, Y => n249);
   U239 : BUFX2 port map( A => keyi_0_port, Y => n258);
   U240 : AND2X2 port map( A => n270, B => n1223, Y => n47);
   U244 : INVX4 port map( A => RST, Y => n307);
   n49 <= '1';
   n52 <= '1';
   n54 <= '1';
   n62 <= '1';
   n64 <= '1';
   n117 <= '1';
   n121 <= '1';
   n122 <= '1';
   n129 <= '1';
   n131 <= '1';
   n135 <= '1';
   n136 <= '1';
   n141 <= '1';
   n151 <= '1';
   n160 <= '1';
   n161 <= '1';
   n172 <= '1';
   n175 <= '1';
   n177 <= '1';
   n180 <= '1';
   n185 <= '1';
   n187 <= '1';
   n188 <= '1';
   n196 <= '1';
   n203 <= '1';
   n206 <= '1';
   n208 <= '1';
   n210 <= '1';
   n212 <= '1';
   n214 <= '1';
   U331 : OR2X2 port map( A => n1299, B => n1484, Y => n216);
   U333 : INVX2 port map( A => n216, Y => n1432);
   U335 : INVX2 port map( A => n42, Y => n630);
   U337 : INVX1 port map( A => n1476, Y => n218);
   U338 : INVX2 port map( A => n218, Y => n220);
   U341 : BUFX2 port map( A => n244, Y => n237);
   U344 : INVX2 port map( A => n1501, Y => n626);
   U347 : INVX2 port map( A => n34, Y => n230);
   U350 : NOR2X1 port map( A => n1495, B => n235, Y => n1511);
   U353 : NAND2X1 port map( A => n632, B => n230, Y => n235);
   U356 : INVX1 port map( A => n1503, Y => n553);
   U359 : INVX2 port map( A => n238, Y => n1300);
   U362 : INVX2 port map( A => n277, Y => n280);
   U365 : INVX1 port map( A => state_2_port, Y => n624);
   U368 : NAND3X1 port map( A => n277, B => n1457, C => n47, Y => n238);
   U371 : INVX1 port map( A => n47, Y => n282);
   U374 : NOR2X1 port map( A => n1495, B => n239, Y => n1599);
   U377 : NAND2X1 port map( A => n632, B => n1501, Y => n239);
   U380 : INVX2 port map( A => n1275, Y => n240);
   U383 : INVX2 port map( A => n1275, Y => n421);
   U386 : INVX2 port map( A => n337, Y => n317);
   U389 : INVX2 port map( A => n335, Y => n318);
   U392 : INVX2 port map( A => n331, Y => n327);
   U395 : INVX2 port map( A => n333, Y => n326);
   U398 : INVX2 port map( A => n339, Y => n311);
   U401 : BUFX2 port map( A => n345, Y => n341);
   U404 : BUFX2 port map( A => n347, Y => n339);
   U407 : BUFX2 port map( A => n329, Y => n337);
   U410 : BUFX2 port map( A => n347, Y => n335);
   U413 : BUFX2 port map( A => n329, Y => n333);
   U416 : BUFX2 port map( A => n349, Y => n331);
   U419 : BUFX2 port map( A => n349, Y => n329);
   U422 : BUFX2 port map( A => n345, Y => n343);
   U425 : INVX2 port map( A => n1475, Y => n612);
   U428 : AND2X2 port map( A => n421, B => n543, Y => n241);
   U431 : INVX2 port map( A => n1271, Y => n287);
   U434 : NOR2X1 port map( A => n1305, B => n1304, Y => n244);
   U502 : INVX2 port map( A => n1566, Y => n297);
   U505 : INVX2 port map( A => n305, Y => n347);
   U508 : INVX2 port map( A => n305, Y => n345);
   U511 : INVX2 port map( A => n305, Y => n349);
   U514 : INVX1 port map( A => n1193, Y => n262);
   U517 : INVX2 port map( A => n1455, Y => n616);
   U520 : INVX2 port map( A => n1254, Y => n419);
   U523 : INVX2 port map( A => n1599, Y => n270);
   U525 : INVX2 port map( A => n1297, Y => n292);
   U526 : INVX2 port map( A => n247, Y => n275);
   U531 : INVX2 port map( A => n246, Y => n285);
   U533 : INVX2 port map( A => n307, Y => n305);
   U535 : INVX2 port map( A => n1457, Y => n604);
   U537 : OR2X2 port map( A => n216, B => n1229, Y => n246);
   U539 : OR2X2 port map( A => n220, B => n1519, Y => n247);
   U541 : INVX2 port map( A => n1571, Y => n277);
   U543 : INVX2 port map( A => n1203, Y => n605);
   U545 : INVX2 port map( A => keyi_1_port, Y => n958);
   U547 : BUFX2 port map( A => n1270, Y => n253);
   U549 : BUFX2 port map( A => n1270, Y => n255);
   U554 : INVX2 port map( A => keyi_2_port, Y => n953);
   U558 : BUFX2 port map( A => keyi_2_port, Y => n261);
   U562 : INVX2 port map( A => n262, Y => n264);
   U565 : INVX4 port map( A => n1154, Y => n957);
   U568 : BUFX2 port map( A => keyi_1_port, Y => n265);
   U571 : INVX1 port map( A => n1315, Y => n488);
   U574 : INVX1 port map( A => n1453, Y => n541);
   U577 : OR2X2 port map( A => n419, B => n946, Y => n267);
   U580 : NAND2X1 port map( A => n267, B => n1255, Y => n1003);
   U584 : NAND2X1 port map( A => n369, B => n932, Y => n351);
   U585 : OAI21X1 port map( A => n932, B => n369, C => n351, Y => N442);
   U588 : NOR2X1 port map( A => n351, B => si_2_port, Y => n355);
   U590 : AOI21X1 port map( A => n351, B => si_2_port, C => n355, Y => n353);
   U592 : NAND2X1 port map( A => n355, B => n367, Y => n357);
   U594 : OAI21X1 port map( A => n355, B => n367, C => n357, Y => N444);
   U596 : NOR2X1 port map( A => n357, B => si_4_port, Y => n361);
   U598 : AOI21X1 port map( A => n357, B => si_4_port, C => n361, Y => n359);
   U600 : NAND2X1 port map( A => n361, B => n935, Y => n363);
   U602 : OAI21X1 port map( A => n361, B => n935, C => n363, Y => N446);
   U608 : XNOR2X1 port map( A => si_6_port, B => n363, Y => N447);
   U611 : NOR2X1 port map( A => si_6_port, B => n363, Y => n365);
   U614 : XOR2X1 port map( A => si_7_port, B => n365, Y => N448);
   U617 : INVX2 port map( A => si_3_port, Y => n367);
   U620 : INVX2 port map( A => si_1_port, Y => n369);
   U623 : INVX2 port map( A => n359, Y => N445);
   U626 : INVX2 port map( A => n353, Y => N443);
   U627 : INVX2 port map( A => KEY_ERROR, Y => n371);
   U629 : INVX2 port map( A => BYTE_READY, Y => n373);
   U630 : INVX2 port map( A => n1509, Y => n375);
   U636 : INVX2 port map( A => OPCODE(1), Y => n377);
   U640 : INVX2 port map( A => OPCODE(0), Y => n379);
   U642 : INVX2 port map( A => nextProcessedData_7_port, Y => n381);
   U644 : INVX2 port map( A => n1388, Y => n383);
   U645 : INVX2 port map( A => nextProcessedData_6_port, Y => n385);
   U648 : INVX2 port map( A => n1381, Y => n387);
   U651 : INVX2 port map( A => nextProcessedData_5_port, Y => n389);
   U658 : INVX2 port map( A => n1382, Y => n391);
   U661 : INVX2 port map( A => nextProcessedData_4_port, Y => n393);
   U670 : INVX2 port map( A => n1383, Y => n395);
   U671 : INVX2 port map( A => nextProcessedData_3_port, Y => n397);
   U674 : INVX2 port map( A => n1384, Y => n399);
   U675 : INVX2 port map( A => nextProcessedData_2_port, Y => n401);
   U676 : INVX2 port map( A => n1385, Y => n403);
   U680 : INVX2 port map( A => nextProcessedData_1_port, Y => n405);
   U682 : INVX2 port map( A => n1386, Y => n407_port);
   U683 : INVX2 port map( A => nextProcessedData_0_port, Y => n409_port);
   U687 : INVX2 port map( A => n1387, Y => n411_port);
   U688 : INVX2 port map( A => prefillCounter_0_port, Y => n413_port);
   U689 : INVX2 port map( A => nfdata_0_port, Y => n415);
   U691 : INVX2 port map( A => nfaddr_0_port, Y => n417);
   U695 : INVX2 port map( A => n1263, Y => n423);
   U698 : INVX2 port map( A => n1264, Y => n425_port);
   U701 : INVX2 port map( A => n1265, Y => n427_port);
   U704 : INVX2 port map( A => n1266, Y => n429_port);
   U707 : INVX2 port map( A => n1267, Y => n431_port);
   U710 : INVX2 port map( A => n1268, Y => n433);
   U713 : INVX2 port map( A => n1269, Y => n435);
   U717 : INVX2 port map( A => n1272, Y => n437);
   U718 : INVX2 port map( A => n1285, Y => n439);
   U719 : INVX2 port map( A => n1286, Y => n441);
   U720 : INVX2 port map( A => n1245, Y => n443_port);
   U725 : INVX2 port map( A => n1231, Y => n445_port);
   U726 : INVX2 port map( A => n1227, Y => n447_port);
   U728 : INVX2 port map( A => nfdata_7_port, Y => n449_port);
   U729 : INVX2 port map( A => nfdata_6_port, Y => n451_port);
   U730 : INVX2 port map( A => nfdata_5_port, Y => n453_port);
   U731 : INVX2 port map( A => nfdata_4_port, Y => n455_port);
   U734 : INVX2 port map( A => nfdata_3_port, Y => n458);
   U736 : INVX2 port map( A => nfdata_2_port, Y => n459);
   U740 : INVX2 port map( A => nfdata_1_port, Y => n462);
   U742 : INVX2 port map( A => n1577, Y => n463);
   U744 : INVX2 port map( A => n1298, Y => n465);
   U747 : INVX2 port map( A => n1296, Y => n467);
   U749 : INVX2 port map( A => n1295, Y => n469);
   U753 : INVX2 port map( A => n1294, Y => n471);
   U756 : INVX2 port map( A => n1293, Y => n473_port);
   U758 : INVX2 port map( A => n1292, Y => n475_port);
   U763 : INVX2 port map( A => n1291, Y => n480_port);
   U768 : INVX2 port map( A => n1290, Y => n482_port);
   U770 : INVX2 port map( A => n1435, Y => n498_port);
   U773 : INVX2 port map( A => nfaddr_1_port, Y => n501_port);
   U776 : INVX2 port map( A => nfaddr_2_port, Y => n503_port);
   U777 : INVX2 port map( A => nfaddr_3_port, Y => n504);
   U779 : INVX2 port map( A => nfaddr_4_port, Y => n505);
   U782 : INVX2 port map( A => nfaddr_5_port, Y => n506);
   U786 : INVX2 port map( A => nfaddr_6_port, Y => n507);
   U789 : INVX2 port map( A => nfaddr_7_port, Y => n509);
   U791 : INVX2 port map( A => n1393, Y => n512_port);
   U793 : INVX2 port map( A => n1488, Y => n514_port);
   U795 : INVX2 port map( A => n1518, Y => n516_port);
   U796 : INVX2 port map( A => n1438, Y => n518_port);
   U798 : INVX2 port map( A => n1389, Y => n520_port);
   U802 : INVX2 port map( A => n1299, Y => n522_port);
   U803 : INVX2 port map( A => n1207, Y => n524_port);
   U805 : INVX2 port map( A => n1434, Y => n528);
   U810 : INVX2 port map( A => n1205, Y => n540);
   U811 : INVX2 port map( A => n1487, Y => n542);
   U813 : INVX2 port map( A => n1511, Y => n543);
   U814 : INVX2 port map( A => n1391, Y => n545);
   U820 : INVX2 port map( A => n1495, Y => n547);
   U821 : INVX2 port map( A => n1228, Y => n549);
   U823 : INVX2 port map( A => n1450, Y => n551);
   U824 : INVX2 port map( A => n1579, Y => n555);
   U830 : INVX2 port map( A => n1582, Y => n557);
   U831 : INVX2 port map( A => n1585, Y => n562);
   U833 : INVX2 port map( A => n1588, Y => n569);
   U834 : INVX2 port map( A => n1591, Y => n571);
   U840 : INVX2 port map( A => n1594, Y => n572);
   U841 : INVX2 port map( A => n1597, Y => n575);
   U843 : INVX2 port map( A => n1601, Y => n577);
   U844 : INVX2 port map( A => state_1_port, Y => n579);
   U850 : INVX2 port map( A => n1247, Y => n581);
   U851 : INVX2 port map( A => n1494, Y => n592);
   U853 : INVX2 port map( A => n1208, Y => n594);
   U854 : INVX2 port map( A => n1491, Y => n600);
   U860 : INVX2 port map( A => n1523, Y => n606);
   U861 : INVX2 port map( A => n1287, Y => n610);
   U863 : INVX2 port map( A => n1520, Y => n614);
   U864 : INVX2 port map( A => n1456, Y => n618);
   U870 : INVX2 port map( A => n1525, Y => n629);
   U871 : INVX2 port map( A => state_0_port, Y => n632);
   U873 : INVX2 port map( A => state_3_port, Y => n636);
   U874 : INVX2 port map( A => keyTable_7_0_port, Y => n637);
   U881 : INVX2 port map( A => keyTable_7_1_port, Y => n638);
   U883 : INVX2 port map( A => keyTable_7_2_port, Y => n648);
   U886 : INVX2 port map( A => keyTable_7_3_port, Y => n649);
   U888 : INVX2 port map( A => keyTable_7_4_port, Y => n650);
   U889 : INVX2 port map( A => keyTable_7_5_port, Y => n651);
   U891 : INVX2 port map( A => keyTable_7_6_port, Y => n692);
   U893 : INVX2 port map( A => keyTable_7_7_port, Y => n701);
   U895 : INVX2 port map( A => keyTable_6_0_port, Y => n746);
   U897 : INVX2 port map( A => keyTable_6_1_port, Y => n748);
   U899 : INVX2 port map( A => keyTable_6_2_port, Y => n750);
   U900 : INVX2 port map( A => keyTable_6_3_port, Y => n752);
   U902 : INVX2 port map( A => keyTable_6_4_port, Y => n754);
   U903 : INVX2 port map( A => keyTable_6_5_port, Y => n756);
   U904 : INVX2 port map( A => keyTable_6_6_port, Y => n758);
   U905 : INVX2 port map( A => keyTable_6_7_port, Y => n760);
   U906 : INVX2 port map( A => keyTable_5_0_port, Y => n761);
   U907 : INVX2 port map( A => keyTable_5_1_port, Y => n762);
   U908 : INVX2 port map( A => keyTable_5_2_port, Y => n763);
   U909 : INVX2 port map( A => keyTable_5_3_port, Y => n764);
   U910 : INVX2 port map( A => keyTable_5_4_port, Y => n765);
   U911 : INVX2 port map( A => keyTable_5_5_port, Y => n766);
   U912 : INVX2 port map( A => keyTable_5_6_port, Y => n767);
   U913 : INVX2 port map( A => keyTable_5_7_port, Y => n768);
   U914 : INVX2 port map( A => keyTable_4_0_port, Y => n769);
   U915 : INVX2 port map( A => keyTable_4_1_port, Y => n770);
   U916 : INVX2 port map( A => keyTable_4_2_port, Y => n771);
   U917 : INVX2 port map( A => keyTable_4_3_port, Y => n772);
   U918 : INVX2 port map( A => keyTable_4_4_port, Y => n773);
   U919 : INVX2 port map( A => keyTable_4_5_port, Y => n774);
   U920 : INVX2 port map( A => keyTable_4_6_port, Y => n775);
   U921 : INVX2 port map( A => keyTable_4_7_port, Y => n776);
   U922 : INVX2 port map( A => keyTable_3_0_port, Y => n777);
   U923 : INVX2 port map( A => keyTable_3_1_port, Y => n778);
   U924 : INVX2 port map( A => keyTable_3_2_port, Y => n779);
   U925 : INVX2 port map( A => keyTable_3_3_port, Y => n780);
   U926 : INVX2 port map( A => keyTable_3_4_port, Y => n781);
   U927 : INVX2 port map( A => keyTable_3_5_port, Y => n782);
   U928 : INVX2 port map( A => keyTable_3_6_port, Y => n783);
   U929 : INVX2 port map( A => keyTable_3_7_port, Y => n784);
   U930 : INVX2 port map( A => keyTable_2_0_port, Y => n785);
   U931 : INVX2 port map( A => keyTable_2_1_port, Y => n786);
   U932 : INVX2 port map( A => keyTable_2_2_port, Y => n787);
   U933 : INVX2 port map( A => keyTable_2_3_port, Y => n788);
   U934 : INVX2 port map( A => keyTable_2_4_port, Y => n789);
   U935 : INVX2 port map( A => keyTable_2_5_port, Y => n790);
   U936 : INVX2 port map( A => keyTable_2_6_port, Y => n791);
   U937 : INVX2 port map( A => keyTable_2_7_port, Y => n864);
   U938 : INVX2 port map( A => keyTable_1_0_port, Y => n865);
   U939 : INVX2 port map( A => keyTable_1_1_port, Y => n866);
   U940 : INVX2 port map( A => keyTable_1_2_port, Y => n867);
   U941 : INVX2 port map( A => keyTable_1_3_port, Y => n868);
   U942 : INVX2 port map( A => keyTable_1_4_port, Y => n869);
   U943 : INVX2 port map( A => keyTable_1_5_port, Y => n870);
   U944 : INVX2 port map( A => keyTable_1_6_port, Y => n871);
   U945 : INVX2 port map( A => keyTable_0_6_port, Y => n883);
   U946 : INVX2 port map( A => keyTable_0_5_port, Y => n884);
   U947 : INVX2 port map( A => keyTable_0_4_port, Y => n885);
   U948 : INVX2 port map( A => keyTable_0_3_port, Y => n886);
   U949 : INVX2 port map( A => keyTable_0_2_port, Y => n887);
   U950 : INVX2 port map( A => keyTable_0_1_port, Y => n888);
   U951 : INVX2 port map( A => keyTable_0_0_port, Y => n889);
   U952 : INVX2 port map( A => keyTable_1_7_port, Y => n890);
   U953 : INVX2 port map( A => keyTable_0_7_port, Y => n916);
   U954 : INVX2 port map( A => prefillCounter_7_port, Y => n917);
   U955 : INVX2 port map( A => prefillCounter_1_port, Y => n918);
   U956 : INVX2 port map( A => prefillCounter_2_port, Y => n919);
   U957 : INVX2 port map( A => prefillCounter_3_port, Y => n920);
   U958 : INVX2 port map( A => prefillCounter_4_port, Y => n921);
   U959 : INVX2 port map( A => prefillCounter_5_port, Y => n922);
   U960 : INVX2 port map( A => prefillCounter_6_port, Y => n923);
   U961 : INVX2 port map( A => temp_7_port, Y => n924);
   U962 : INVX2 port map( A => temp_0_port, Y => n925);
   U963 : INVX2 port map( A => temp_1_port, Y => n926);
   U964 : INVX2 port map( A => temp_2_port, Y => n927);
   U965 : INVX2 port map( A => temp_3_port, Y => n928);
   U966 : INVX2 port map( A => temp_4_port, Y => n929);
   U967 : INVX2 port map( A => temp_5_port, Y => n930);
   U968 : INVX2 port map( A => temp_6_port, Y => n931);
   U969 : INVX2 port map( A => si_0_port, Y => n932);
   U970 : INVX2 port map( A => si_2_port, Y => n933);
   U971 : INVX2 port map( A => si_4_port, Y => n934);
   U972 : INVX2 port map( A => si_5_port, Y => n935);
   U973 : INVX2 port map( A => si_6_port, Y => n936);
   U974 : INVX2 port map( A => si_7_port, Y => n937);
   U975 : INVX2 port map( A => intj_7_port, Y => n938);
   U976 : INVX2 port map( A => intj_0_port, Y => n939);
   U977 : INVX2 port map( A => intj_1_port, Y => n940);
   U978 : INVX2 port map( A => intj_2_port, Y => n941);
   U979 : INVX2 port map( A => intj_3_port, Y => n942);
   U980 : INVX2 port map( A => intj_4_port, Y => n943);
   U981 : INVX2 port map( A => intj_5_port, Y => n944);
   U982 : INVX2 port map( A => intj_6_port, Y => n945);
   U983 : INVX2 port map( A => sj_7_port, Y => n946);
   U984 : INVX2 port map( A => sj_6_port, Y => n947);
   U985 : INVX2 port map( A => sj_5_port, Y => n948);
   U986 : INVX2 port map( A => sj_4_port, Y => n949);
   U987 : INVX2 port map( A => sj_3_port, Y => n950);
   U988 : INVX2 port map( A => sj_2_port, Y => n951);
   U989 : INVX2 port map( A => sj_1_port, Y => n952);
   U990 : INVX2 port map( A => currentProcessedData_0_port, Y => n960);
   U991 : INVX2 port map( A => currentProcessedData_1_port, Y => n961);
   U992 : INVX2 port map( A => currentProcessedData_2_port, Y => n962);
   U993 : INVX2 port map( A => currentProcessedData_3_port, Y => n963);
   U994 : INVX2 port map( A => currentProcessedData_4_port, Y => n964);
   U995 : INVX2 port map( A => currentProcessedData_5_port, Y => n965);
   U996 : INVX2 port map( A => currentProcessedData_6_port, Y => n966);
   U997 : INVX2 port map( A => currentProcessedData_7_port, Y => n967);
   U998 : INVX2 port map( A => faddr_7_port, Y => n968);
   U999 : INVX2 port map( A => faddr_6_port, Y => n969);
   U1000 : INVX2 port map( A => faddr_5_port, Y => n970);
   U1001 : INVX2 port map( A => faddr_4_port, Y => n971);
   U1002 : INVX2 port map( A => faddr_3_port, Y => n972);
   U1003 : INVX2 port map( A => faddr_2_port, Y => n973);
   U1004 : INVX2 port map( A => faddr_1_port, Y => n974);
   U1005 : INVX2 port map( A => faddr_0_port, Y => n975);
   U1006 : INVX2 port map( A => fdata_7_port, Y => n976);
   U1007 : INVX2 port map( A => fdata_6_port, Y => n977);
   U1008 : INVX2 port map( A => fdata_5_port, Y => n978);
   U1009 : INVX2 port map( A => fdata_4_port, Y => n979);
   U1010 : INVX2 port map( A => fdata_3_port, Y => n980);
   U1011 : INVX2 port map( A => fdata_2_port, Y => n981);
   U1012 : INVX2 port map( A => fdata_1_port, Y => n982);
   U1013 : INVX2 port map( A => fdata_0_port, Y => n983);
   n984 <= '0';
   n985 <= '0';

end SYN_bksa;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity transmitter_block_0 is

   port( PRGA_OUT : in std_logic_vector (7 downto 0);  clk, p_ready : in 
         std_logic;  prga_opcode : in std_logic_vector (1 downto 0);  rst : in 
         std_logic;  SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE : out std_logic);

end transmitter_block_0;

architecture SYN_struct of transmitter_block_0 is

   component tx_timer_0
      port( CLK, RST, SENDING : in std_logic;  SHIFT_ENABLE_R, SHIFT_ENABLE_E :
            out std_logic);
   end component;
   
   component tx_tcu_0
      port( clk, rst, p_ready, t_bitstuff : in std_logic;  PRGA_OUT : in 
            std_logic_vector (7 downto 0);  prga_opcode : in std_logic_vector 
            (1 downto 0);  t_crc : in std_logic_vector (15 downto 0);  sending,
            EOP, next_byte : out std_logic;  send_data : out std_logic_vector 
            (7 downto 0);  t_strobe : out std_logic);
   end component;
   
   component tx_shiftreg_0
      port( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe : in std_logic;  
            send_data : in std_logic_vector (7 downto 0);  d_encode : out 
            std_logic);
   end component;
   
   component tx_encode_0
      port( clk, rst, SHIFT_ENABLE_E, d_encode, EOP : in std_logic;  t_bitstuff
            , dp_tx_out, dm_tx_out : out std_logic);
   end component;
   
   component tx_CRC_CALC_0
      port( CLK, RST, EOP, T_STROBE : in std_logic;  PRGA_OPCODE : in 
            std_logic_vector (1 downto 0);  PRGA_OUT : in std_logic_vector (7 
            downto 0);  TX_CRC : out std_logic_vector (15 downto 0));
   end component;
   
   signal SENDING_port, t_strobe, EOP, TX_CRC_15_port, TX_CRC_14_port, 
      TX_CRC_13_port, TX_CRC_12_port, TX_CRC_11_port, TX_CRC_10_port, 
      TX_CRC_9_port, TX_CRC_8_port, TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port
      , TX_CRC_4_port, TX_CRC_3_port, TX_CRC_2_port, TX_CRC_1_port, 
      TX_CRC_0_port, SHIFT_ENABLE_E, d_encode, t_bitstuff, SHIFT_ENABLE_R, 
      send_data_7_port, send_data_6_port, send_data_5_port, send_data_4_port, 
      send_data_3_port, send_data_2_port, send_data_1_port, send_data_0_port : 
      std_logic;

begin
   SENDING <= SENDING_port;
   
   U_1 : tx_CRC_CALC_0 port map( CLK => clk, RST => rst, EOP => EOP, T_STROBE 
                           => t_strobe, PRGA_OPCODE(1) => prga_opcode(1), 
                           PRGA_OPCODE(0) => prga_opcode(0), PRGA_OUT(7) => 
                           PRGA_OUT(7), PRGA_OUT(6) => PRGA_OUT(6), PRGA_OUT(5)
                           => PRGA_OUT(5), PRGA_OUT(4) => PRGA_OUT(4), 
                           PRGA_OUT(3) => PRGA_OUT(3), PRGA_OUT(2) => 
                           PRGA_OUT(2), PRGA_OUT(1) => PRGA_OUT(1), PRGA_OUT(0)
                           => PRGA_OUT(0), TX_CRC(15) => TX_CRC_15_port, 
                           TX_CRC(14) => TX_CRC_14_port, TX_CRC(13) => 
                           TX_CRC_13_port, TX_CRC(12) => TX_CRC_12_port, 
                           TX_CRC(11) => TX_CRC_11_port, TX_CRC(10) => 
                           TX_CRC_10_port, TX_CRC(9) => TX_CRC_9_port, 
                           TX_CRC(8) => TX_CRC_8_port, TX_CRC(7) => 
                           TX_CRC_7_port, TX_CRC(6) => TX_CRC_6_port, TX_CRC(5)
                           => TX_CRC_5_port, TX_CRC(4) => TX_CRC_4_port, 
                           TX_CRC(3) => TX_CRC_3_port, TX_CRC(2) => 
                           TX_CRC_2_port, TX_CRC(1) => TX_CRC_1_port, TX_CRC(0)
                           => TX_CRC_0_port);
   U_0 : tx_encode_0 port map( clk => clk, rst => rst, SHIFT_ENABLE_E => 
                           SHIFT_ENABLE_E, d_encode => d_encode, EOP => EOP, 
                           t_bitstuff => t_bitstuff, dp_tx_out => dp_tx_out, 
                           dm_tx_out => dm_tx_out);
   U_2 : tx_shiftreg_0 port map( clk => clk, rst => rst, SHIFT_ENABLE_R => 
                           SHIFT_ENABLE_R, t_bitstuff => t_bitstuff, t_strobe 
                           => t_strobe, send_data(7) => send_data_7_port, 
                           send_data(6) => send_data_6_port, send_data(5) => 
                           send_data_5_port, send_data(4) => send_data_4_port, 
                           send_data(3) => send_data_3_port, send_data(2) => 
                           send_data_2_port, send_data(1) => send_data_1_port, 
                           send_data(0) => send_data_0_port, d_encode => 
                           d_encode);
   U_3 : tx_tcu_0 port map( clk => clk, rst => rst, p_ready => p_ready, 
                           t_bitstuff => t_bitstuff, PRGA_OUT(7) => PRGA_OUT(7)
                           , PRGA_OUT(6) => PRGA_OUT(6), PRGA_OUT(5) => 
                           PRGA_OUT(5), PRGA_OUT(4) => PRGA_OUT(4), PRGA_OUT(3)
                           => PRGA_OUT(3), PRGA_OUT(2) => PRGA_OUT(2), 
                           PRGA_OUT(1) => PRGA_OUT(1), PRGA_OUT(0) => 
                           PRGA_OUT(0), prga_opcode(1) => prga_opcode(1), 
                           prga_opcode(0) => prga_opcode(0), t_crc(15) => 
                           TX_CRC_15_port, t_crc(14) => TX_CRC_14_port, 
                           t_crc(13) => TX_CRC_13_port, t_crc(12) => 
                           TX_CRC_12_port, t_crc(11) => TX_CRC_11_port, 
                           t_crc(10) => TX_CRC_10_port, t_crc(9) => 
                           TX_CRC_9_port, t_crc(8) => TX_CRC_8_port, t_crc(7) 
                           => TX_CRC_7_port, t_crc(6) => TX_CRC_6_port, 
                           t_crc(5) => TX_CRC_5_port, t_crc(4) => TX_CRC_4_port
                           , t_crc(3) => TX_CRC_3_port, t_crc(2) => 
                           TX_CRC_2_port, t_crc(1) => TX_CRC_1_port, t_crc(0) 
                           => TX_CRC_0_port, sending => SENDING_port, EOP => 
                           EOP, next_byte => NEXT_BYTE, send_data(7) => 
                           send_data_7_port, send_data(6) => send_data_6_port, 
                           send_data(5) => send_data_5_port, send_data(4) => 
                           send_data_4_port, send_data(3) => send_data_3_port, 
                           send_data(2) => send_data_2_port, send_data(1) => 
                           send_data_1_port, send_data(0) => send_data_0_port, 
                           t_strobe => t_strobe);
   U_4 : tx_timer_0 port map( CLK => clk, RST => rst, SENDING => SENDING_port, 
                           SHIFT_ENABLE_R => SHIFT_ENABLE_R, SHIFT_ENABLE_E => 
                           SHIFT_ENABLE_E);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity receiver_block_rewire_0 is

   port( CLK, DM1_RX, DP1_RX, RST : in std_logic;  BS_ERROR, CRC_ERROR, 
         EOP_external : out std_logic;  OPCODE : out std_logic_vector (1 downto
         0);  RCV_DATA : out std_logic_vector (7 downto 0);  R_ERROR, W_ENABLE 
         : out std_logic);

end receiver_block_rewire_0;

architecture SYN_struct of receiver_block_rewire_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component rx_timer_0
      port( CLK, RST, D_EDGE, RCVING : in std_logic;  SHIFT_ENABLE : out 
            std_logic);
   end component;
   
   component rx_shift_reg_0
      port( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF : in std_logic;  RCV_DATA 
            : out std_logic_vector (7 downto 0));
   end component;
   
   component rx_rcu_0
      port( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR : in 
            std_logic;  RX_CRC, RX_CHECK_CRC : in std_logic_vector (15 downto 
            0);  RCV_DATA : in std_logic_vector (7 downto 0);  RCVING, W_ENABLE
            , R_ERROR, CRC_ERROR : out std_logic;  OPCODE : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component rx_eopdetect_0
      port( DP1_RX, DM1_RX : in std_logic;  EOP : out std_logic);
   end component;
   
   component rx_edgedetect_0
      port( CLK, RST, DP1_RX : in std_logic;  D_EDGE : out std_logic);
   end component;
   
   component rx_decode_0
      port( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP : in std_logic;  D_ORIG, 
            BITSTUFF, BS_ERROR : out std_logic);
   end component;
   
   component rx_accumulator_0
      port( CLK, RST : in std_logic;  RCV_DATA : in std_logic_vector (7 downto 
            0);  W_ENABLE : in std_logic;  rx_CHECK_CRC : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component rx_CRC_CALC_0
      port( CLK, RST, W_ENABLE : in std_logic;  OPCODE : in std_logic_vector (1
            downto 0);  RCV_DATA : in std_logic_vector (7 downto 0);  RX_CRC : 
            out std_logic_vector (15 downto 0));
   end component;
   
   signal BS_ERROR_port, EOP_external_port, OPCODE_1_port, OPCODE_0_port, 
      RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      W_ENABLE_port, RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, 
      RX_CRC_12_port, RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, 
      RX_CRC_8_port, RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port
      , RX_CRC_3_port, RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port, 
      rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, rx_CHECK_CRC_13_port, 
      rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, rx_CHECK_CRC_10_port, 
      rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, rx_CHECK_CRC_7_port, 
      rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, rx_CHECK_CRC_4_port, 
      rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, rx_CHECK_CRC_1_port, 
      rx_CHECK_CRC_0_port, SHIFT_ENABLE, BITSTUFF, D_ORIG, D_EDGE, RCVING, n1, 
      n2 : std_logic;

begin
   BS_ERROR <= BS_ERROR_port;
   EOP_external <= EOP_external_port;
   OPCODE <= ( OPCODE_1_port, OPCODE_0_port );
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   W_ENABLE <= W_ENABLE_port;
   
   U_2 : rx_CRC_CALC_0 port map( CLK => CLK, RST => n1, W_ENABLE => 
                           W_ENABLE_port, OPCODE(1) => OPCODE_1_port, OPCODE(0)
                           => OPCODE_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, RX_CRC(15) => 
                           RX_CRC_15_port, RX_CRC(14) => RX_CRC_14_port, 
                           RX_CRC(13) => RX_CRC_13_port, RX_CRC(12) => 
                           RX_CRC_12_port, RX_CRC(11) => RX_CRC_11_port, 
                           RX_CRC(10) => RX_CRC_10_port, RX_CRC(9) => 
                           RX_CRC_9_port, RX_CRC(8) => RX_CRC_8_port, RX_CRC(7)
                           => RX_CRC_7_port, RX_CRC(6) => RX_CRC_6_port, 
                           RX_CRC(5) => RX_CRC_5_port, RX_CRC(4) => 
                           RX_CRC_4_port, RX_CRC(3) => RX_CRC_3_port, RX_CRC(2)
                           => RX_CRC_2_port, RX_CRC(1) => RX_CRC_1_port, 
                           RX_CRC(0) => RX_CRC_0_port);
   U_3 : rx_accumulator_0 port map( CLK => CLK, RST => n1, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           W_ENABLE => W_ENABLE_port, rx_CHECK_CRC(15) => 
                           rx_CHECK_CRC_15_port, rx_CHECK_CRC(14) => 
                           rx_CHECK_CRC_14_port, rx_CHECK_CRC(13) => 
                           rx_CHECK_CRC_13_port, rx_CHECK_CRC(12) => 
                           rx_CHECK_CRC_12_port, rx_CHECK_CRC(11) => 
                           rx_CHECK_CRC_11_port, rx_CHECK_CRC(10) => 
                           rx_CHECK_CRC_10_port, rx_CHECK_CRC(9) => 
                           rx_CHECK_CRC_9_port, rx_CHECK_CRC(8) => 
                           rx_CHECK_CRC_8_port, rx_CHECK_CRC(7) => 
                           rx_CHECK_CRC_7_port, rx_CHECK_CRC(6) => 
                           rx_CHECK_CRC_6_port, rx_CHECK_CRC(5) => 
                           rx_CHECK_CRC_5_port, rx_CHECK_CRC(4) => 
                           rx_CHECK_CRC_4_port, rx_CHECK_CRC(3) => 
                           rx_CHECK_CRC_3_port, rx_CHECK_CRC(2) => 
                           rx_CHECK_CRC_2_port, rx_CHECK_CRC(1) => 
                           rx_CHECK_CRC_1_port, rx_CHECK_CRC(0) => 
                           rx_CHECK_CRC_0_port);
   U_1 : rx_decode_0 port map( CLK => CLK, RST => n1, DP1_RX => DP1_RX, 
                           SHIFT_ENABLE => SHIFT_ENABLE, EOP => 
                           EOP_external_port, D_ORIG => D_ORIG, BITSTUFF => 
                           BITSTUFF, BS_ERROR => BS_ERROR_port);
   U_0 : rx_edgedetect_0 port map( CLK => CLK, RST => n1, DP1_RX => DP1_RX, 
                           D_EDGE => D_EDGE);
   U_4 : rx_eopdetect_0 port map( DP1_RX => DP1_RX, DM1_RX => DM1_RX, EOP => 
                           EOP_external_port);
   U_5 : rx_rcu_0 port map( CLK => CLK, RST => n1, D_EDGE => D_EDGE, EOP => 
                           EOP_external_port, SHIFT_ENABLE => SHIFT_ENABLE, 
                           BITSTUFF => BITSTUFF, BS_ERROR => BS_ERROR_port, 
                           RX_CRC(15) => RX_CRC_15_port, RX_CRC(14) => 
                           RX_CRC_14_port, RX_CRC(13) => RX_CRC_13_port, 
                           RX_CRC(12) => RX_CRC_12_port, RX_CRC(11) => 
                           RX_CRC_11_port, RX_CRC(10) => RX_CRC_10_port, 
                           RX_CRC(9) => RX_CRC_9_port, RX_CRC(8) => 
                           RX_CRC_8_port, RX_CRC(7) => RX_CRC_7_port, RX_CRC(6)
                           => RX_CRC_6_port, RX_CRC(5) => RX_CRC_5_port, 
                           RX_CRC(4) => RX_CRC_4_port, RX_CRC(3) => 
                           RX_CRC_3_port, RX_CRC(2) => RX_CRC_2_port, RX_CRC(1)
                           => RX_CRC_1_port, RX_CRC(0) => RX_CRC_0_port, 
                           RX_CHECK_CRC(15) => rx_CHECK_CRC_15_port, 
                           RX_CHECK_CRC(14) => rx_CHECK_CRC_14_port, 
                           RX_CHECK_CRC(13) => rx_CHECK_CRC_13_port, 
                           RX_CHECK_CRC(12) => rx_CHECK_CRC_12_port, 
                           RX_CHECK_CRC(11) => rx_CHECK_CRC_11_port, 
                           RX_CHECK_CRC(10) => rx_CHECK_CRC_10_port, 
                           RX_CHECK_CRC(9) => rx_CHECK_CRC_9_port, 
                           RX_CHECK_CRC(8) => rx_CHECK_CRC_8_port, 
                           RX_CHECK_CRC(7) => rx_CHECK_CRC_7_port, 
                           RX_CHECK_CRC(6) => rx_CHECK_CRC_6_port, 
                           RX_CHECK_CRC(5) => rx_CHECK_CRC_5_port, 
                           RX_CHECK_CRC(4) => rx_CHECK_CRC_4_port, 
                           RX_CHECK_CRC(3) => rx_CHECK_CRC_3_port, 
                           RX_CHECK_CRC(2) => rx_CHECK_CRC_2_port, 
                           RX_CHECK_CRC(1) => rx_CHECK_CRC_1_port, 
                           RX_CHECK_CRC(0) => rx_CHECK_CRC_0_port, RCV_DATA(7) 
                           => RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           RCVING => RCVING, W_ENABLE => W_ENABLE_port, R_ERROR
                           => R_ERROR, CRC_ERROR => CRC_ERROR, OPCODE(1) => 
                           OPCODE_1_port, OPCODE(0) => OPCODE_0_port);
   U_6 : rx_shift_reg_0 port map( CLK => CLK, RST => n1, SHIFT_ENABLE => 
                           SHIFT_ENABLE, D_ORIG => D_ORIG, BITSTUFF => BITSTUFF
                           , RCV_DATA(7) => RCV_DATA_7_port, RCV_DATA(6) => 
                           RCV_DATA_6_port, RCV_DATA(5) => RCV_DATA_5_port, 
                           RCV_DATA(4) => RCV_DATA_4_port, RCV_DATA(3) => 
                           RCV_DATA_3_port, RCV_DATA(2) => RCV_DATA_2_port, 
                           RCV_DATA(1) => RCV_DATA_1_port, RCV_DATA(0) => 
                           RCV_DATA_0_port);
   U_7 : rx_timer_0 port map( CLK => CLK, RST => n1, D_EDGE => D_EDGE, RCVING 
                           => RCVING, SHIFT_ENABLE => SHIFT_ENABLE);
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity memoryblock_0 is

   port( CLK, NEXT_BYTE : in std_logic;  RCV_DATA : in std_logic_vector (7 
         downto 0);  RCV_OPCODE : in std_logic_vector (1 downto 0);  RST, 
         W_ENABLE, EOP : in std_logic;  EMPTY, FULL, B_READY : out std_logic;  
         PRGA_IN : out std_logic_vector (7 downto 0);  PRGA_OPCODE : out 
         std_logic_vector (1 downto 0));

end memoryblock_0;

architecture SYN_struct of memoryblock_0 is

   component RFIFO_0
      port( CLK, RST, W_ENABLE, R_ENABLE : in std_logic;  RCV_DATA : in 
            std_logic_vector (7 downto 0);  RCV_OPCODE : in std_logic_vector (1
            downto 0);  DATA : out std_logic_vector (7 downto 0);  OUT_OPCODE :
            out std_logic_vector (1 downto 0);  BYTE_COUNT : out 
            std_logic_vector (4 downto 0);  EMPTY, FULL : out std_logic);
   end component;
   
   component RBUFFER_0
      port( CLK, RST, NEXT_BYTE : in std_logic;  DATA : in std_logic_vector (7 
            downto 0);  OPCODE : in std_logic_vector (1 downto 0);  BYTE_COUNT 
            : in std_logic_vector (4 downto 0);  EOP : in std_logic;  B_READY, 
            R_ENABLE : out std_logic;  PRGA_IN : out std_logic_vector (7 downto
            0);  PRGA_OPCODE : out std_logic_vector (1 downto 0));
   end component;
   
   signal BYTE_COUNT_4_port, BYTE_COUNT_3_port, BYTE_COUNT_2_port, 
      BYTE_COUNT_1_port, BYTE_COUNT_0_port, DATA_7_port, DATA_6_port, 
      DATA_5_port, DATA_4_port, DATA_3_port, DATA_2_port, DATA_1_port, 
      DATA_0_port, OUT_OPCODE_1_port, OUT_OPCODE_0_port, R_ENABLE : std_logic;

begin
   
   U_0 : RBUFFER_0 port map( CLK => CLK, RST => RST, NEXT_BYTE => NEXT_BYTE, 
                           DATA(7) => DATA_7_port, DATA(6) => DATA_6_port, 
                           DATA(5) => DATA_5_port, DATA(4) => DATA_4_port, 
                           DATA(3) => DATA_3_port, DATA(2) => DATA_2_port, 
                           DATA(1) => DATA_1_port, DATA(0) => DATA_0_port, 
                           OPCODE(1) => OUT_OPCODE_1_port, OPCODE(0) => 
                           OUT_OPCODE_0_port, BYTE_COUNT(4) => 
                           BYTE_COUNT_4_port, BYTE_COUNT(3) => 
                           BYTE_COUNT_3_port, BYTE_COUNT(2) => 
                           BYTE_COUNT_2_port, BYTE_COUNT(1) => 
                           BYTE_COUNT_1_port, BYTE_COUNT(0) => 
                           BYTE_COUNT_0_port, EOP => EOP, B_READY => B_READY, 
                           R_ENABLE => R_ENABLE, PRGA_IN(7) => PRGA_IN(7), 
                           PRGA_IN(6) => PRGA_IN(6), PRGA_IN(5) => PRGA_IN(5), 
                           PRGA_IN(4) => PRGA_IN(4), PRGA_IN(3) => PRGA_IN(3), 
                           PRGA_IN(2) => PRGA_IN(2), PRGA_IN(1) => PRGA_IN(1), 
                           PRGA_IN(0) => PRGA_IN(0), PRGA_OPCODE(1) => 
                           PRGA_OPCODE(1), PRGA_OPCODE(0) => PRGA_OPCODE(0));
   U_1 : RFIFO_0 port map( CLK => CLK, RST => RST, W_ENABLE => W_ENABLE, 
                           R_ENABLE => R_ENABLE, RCV_DATA(7) => RCV_DATA(7), 
                           RCV_DATA(6) => RCV_DATA(6), RCV_DATA(5) => 
                           RCV_DATA(5), RCV_DATA(4) => RCV_DATA(4), RCV_DATA(3)
                           => RCV_DATA(3), RCV_DATA(2) => RCV_DATA(2), 
                           RCV_DATA(1) => RCV_DATA(1), RCV_DATA(0) => 
                           RCV_DATA(0), RCV_OPCODE(1) => RCV_OPCODE(1), 
                           RCV_OPCODE(0) => RCV_OPCODE(0), DATA(7) => 
                           DATA_7_port, DATA(6) => DATA_6_port, DATA(5) => 
                           DATA_5_port, DATA(4) => DATA_4_port, DATA(3) => 
                           DATA_3_port, DATA(2) => DATA_2_port, DATA(1) => 
                           DATA_1_port, DATA(0) => DATA_0_port, OUT_OPCODE(1) 
                           => OUT_OPCODE_1_port, OUT_OPCODE(0) => 
                           OUT_OPCODE_0_port, BYTE_COUNT(4) => 
                           BYTE_COUNT_4_port, BYTE_COUNT(3) => 
                           BYTE_COUNT_3_port, BYTE_COUNT(2) => 
                           BYTE_COUNT_2_port, BYTE_COUNT(1) => 
                           BYTE_COUNT_1_port, BYTE_COUNT(0) => 
                           BYTE_COUNT_0_port, EMPTY => EMPTY, FULL => FULL);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity EDBlock_0 is

   port( BYTE : in std_logic_vector (7 downto 0);  BYTE_READY, CLK : in 
         std_logic;  OPCODE : in std_logic_vector (1 downto 0);  RST, SERIAL_IN
         : in std_logic;  DATA_IN : in std_logic_vector (7 downto 0);  
         KEY_ERROR, PARITY_ERROR, PDATA_READY : out std_logic;  PROCESSED_DATA 
         : out std_logic_vector (7 downto 0);  PROG_ERROR, RBUF_FULL, W_ENABLE,
         R_ENABLE : out std_logic;  DATA, ADDR : out std_logic_vector (7 downto
         0));

end EDBlock_0;

architecture SYN_struct of EDBlock_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component uart_rcv_block_0
      port( CLK, RST, SERIAL_IN : in std_logic;  KEY_ERROR, PROG_ERROR : out 
            std_logic;  PLAINKEY : out std_logic_vector (63 downto 0);  
            RBUF_FULL, PARITY_ERROR : out std_logic);
   end component;
   
   component KSA_0
      port( KEY : in std_logic_vector (63 downto 0);  CLK, RST, KEY_ERROR, 
            BYTE_READY : in std_logic;  BYTE : in std_logic_vector (7 downto 0)
            ;  OPCODE : in std_logic_vector (1 downto 0);  DATA_IN : in 
            std_logic_vector (7 downto 0);  PROCESSED_DATA : out 
            std_logic_vector (7 downto 0);  PDATA_READY, W_ENABLE, R_ENABLE : 
            out std_logic;  ADDR, DATA : out std_logic_vector (7 downto 0));
   end component;
   
   signal KEY_ERROR_port, PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port,
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port, n1, n2 : std_logic;

begin
   KEY_ERROR <= KEY_ERROR_port;
   
   U_0 : KSA_0 port map( KEY(63) => PLAINKEY_63_port, KEY(62) => 
                           PLAINKEY_62_port, KEY(61) => PLAINKEY_61_port, 
                           KEY(60) => PLAINKEY_60_port, KEY(59) => 
                           PLAINKEY_59_port, KEY(58) => PLAINKEY_58_port, 
                           KEY(57) => PLAINKEY_57_port, KEY(56) => 
                           PLAINKEY_56_port, KEY(55) => PLAINKEY_55_port, 
                           KEY(54) => PLAINKEY_54_port, KEY(53) => 
                           PLAINKEY_53_port, KEY(52) => PLAINKEY_52_port, 
                           KEY(51) => PLAINKEY_51_port, KEY(50) => 
                           PLAINKEY_50_port, KEY(49) => PLAINKEY_49_port, 
                           KEY(48) => PLAINKEY_48_port, KEY(47) => 
                           PLAINKEY_47_port, KEY(46) => PLAINKEY_46_port, 
                           KEY(45) => PLAINKEY_45_port, KEY(44) => 
                           PLAINKEY_44_port, KEY(43) => PLAINKEY_43_port, 
                           KEY(42) => PLAINKEY_42_port, KEY(41) => 
                           PLAINKEY_41_port, KEY(40) => PLAINKEY_40_port, 
                           KEY(39) => PLAINKEY_39_port, KEY(38) => 
                           PLAINKEY_38_port, KEY(37) => PLAINKEY_37_port, 
                           KEY(36) => PLAINKEY_36_port, KEY(35) => 
                           PLAINKEY_35_port, KEY(34) => PLAINKEY_34_port, 
                           KEY(33) => PLAINKEY_33_port, KEY(32) => 
                           PLAINKEY_32_port, KEY(31) => PLAINKEY_31_port, 
                           KEY(30) => PLAINKEY_30_port, KEY(29) => 
                           PLAINKEY_29_port, KEY(28) => PLAINKEY_28_port, 
                           KEY(27) => PLAINKEY_27_port, KEY(26) => 
                           PLAINKEY_26_port, KEY(25) => PLAINKEY_25_port, 
                           KEY(24) => PLAINKEY_24_port, KEY(23) => 
                           PLAINKEY_23_port, KEY(22) => PLAINKEY_22_port, 
                           KEY(21) => PLAINKEY_21_port, KEY(20) => 
                           PLAINKEY_20_port, KEY(19) => PLAINKEY_19_port, 
                           KEY(18) => PLAINKEY_18_port, KEY(17) => 
                           PLAINKEY_17_port, KEY(16) => PLAINKEY_16_port, 
                           KEY(15) => PLAINKEY_15_port, KEY(14) => 
                           PLAINKEY_14_port, KEY(13) => PLAINKEY_13_port, 
                           KEY(12) => PLAINKEY_12_port, KEY(11) => 
                           PLAINKEY_11_port, KEY(10) => PLAINKEY_10_port, 
                           KEY(9) => PLAINKEY_9_port, KEY(8) => PLAINKEY_8_port
                           , KEY(7) => PLAINKEY_7_port, KEY(6) => 
                           PLAINKEY_6_port, KEY(5) => PLAINKEY_5_port, KEY(4) 
                           => PLAINKEY_4_port, KEY(3) => PLAINKEY_3_port, 
                           KEY(2) => PLAINKEY_2_port, KEY(1) => PLAINKEY_1_port
                           , KEY(0) => PLAINKEY_0_port, CLK => CLK, RST => n1, 
                           KEY_ERROR => KEY_ERROR_port, BYTE_READY => 
                           BYTE_READY, BYTE(7) => BYTE(7), BYTE(6) => BYTE(6), 
                           BYTE(5) => BYTE(5), BYTE(4) => BYTE(4), BYTE(3) => 
                           BYTE(3), BYTE(2) => BYTE(2), BYTE(1) => BYTE(1), 
                           BYTE(0) => BYTE(0), OPCODE(1) => OPCODE(1), 
                           OPCODE(0) => OPCODE(0), DATA_IN(7) => DATA_IN(7), 
                           DATA_IN(6) => DATA_IN(6), DATA_IN(5) => DATA_IN(5), 
                           DATA_IN(4) => DATA_IN(4), DATA_IN(3) => DATA_IN(3), 
                           DATA_IN(2) => DATA_IN(2), DATA_IN(1) => DATA_IN(1), 
                           DATA_IN(0) => DATA_IN(0), PROCESSED_DATA(7) => 
                           PROCESSED_DATA(7), PROCESSED_DATA(6) => 
                           PROCESSED_DATA(6), PROCESSED_DATA(5) => 
                           PROCESSED_DATA(5), PROCESSED_DATA(4) => 
                           PROCESSED_DATA(4), PROCESSED_DATA(3) => 
                           PROCESSED_DATA(3), PROCESSED_DATA(2) => 
                           PROCESSED_DATA(2), PROCESSED_DATA(1) => 
                           PROCESSED_DATA(1), PROCESSED_DATA(0) => 
                           PROCESSED_DATA(0), PDATA_READY => PDATA_READY, 
                           W_ENABLE => W_ENABLE, R_ENABLE => R_ENABLE, ADDR(7) 
                           => ADDR(7), ADDR(6) => ADDR(6), ADDR(5) => ADDR(5), 
                           ADDR(4) => ADDR(4), ADDR(3) => ADDR(3), ADDR(2) => 
                           ADDR(2), ADDR(1) => ADDR(1), ADDR(0) => ADDR(0), 
                           DATA(7) => DATA(7), DATA(6) => DATA(6), DATA(5) => 
                           DATA(5), DATA(4) => DATA(4), DATA(3) => DATA(3), 
                           DATA(2) => DATA(2), DATA(1) => DATA(1), DATA(0) => 
                           DATA(0));
   U_1 : uart_rcv_block_0 port map( CLK => CLK, RST => n1, SERIAL_IN => 
                           SERIAL_IN, KEY_ERROR => KEY_ERROR_port, PROG_ERROR 
                           => PROG_ERROR, PLAINKEY(63) => PLAINKEY_63_port, 
                           PLAINKEY(62) => PLAINKEY_62_port, PLAINKEY(61) => 
                           PLAINKEY_61_port, PLAINKEY(60) => PLAINKEY_60_port, 
                           PLAINKEY(59) => PLAINKEY_59_port, PLAINKEY(58) => 
                           PLAINKEY_58_port, PLAINKEY(57) => PLAINKEY_57_port, 
                           PLAINKEY(56) => PLAINKEY_56_port, PLAINKEY(55) => 
                           PLAINKEY_55_port, PLAINKEY(54) => PLAINKEY_54_port, 
                           PLAINKEY(53) => PLAINKEY_53_port, PLAINKEY(52) => 
                           PLAINKEY_52_port, PLAINKEY(51) => PLAINKEY_51_port, 
                           PLAINKEY(50) => PLAINKEY_50_port, PLAINKEY(49) => 
                           PLAINKEY_49_port, PLAINKEY(48) => PLAINKEY_48_port, 
                           PLAINKEY(47) => PLAINKEY_47_port, PLAINKEY(46) => 
                           PLAINKEY_46_port, PLAINKEY(45) => PLAINKEY_45_port, 
                           PLAINKEY(44) => PLAINKEY_44_port, PLAINKEY(43) => 
                           PLAINKEY_43_port, PLAINKEY(42) => PLAINKEY_42_port, 
                           PLAINKEY(41) => PLAINKEY_41_port, PLAINKEY(40) => 
                           PLAINKEY_40_port, PLAINKEY(39) => PLAINKEY_39_port, 
                           PLAINKEY(38) => PLAINKEY_38_port, PLAINKEY(37) => 
                           PLAINKEY_37_port, PLAINKEY(36) => PLAINKEY_36_port, 
                           PLAINKEY(35) => PLAINKEY_35_port, PLAINKEY(34) => 
                           PLAINKEY_34_port, PLAINKEY(33) => PLAINKEY_33_port, 
                           PLAINKEY(32) => PLAINKEY_32_port, PLAINKEY(31) => 
                           PLAINKEY_31_port, PLAINKEY(30) => PLAINKEY_30_port, 
                           PLAINKEY(29) => PLAINKEY_29_port, PLAINKEY(28) => 
                           PLAINKEY_28_port, PLAINKEY(27) => PLAINKEY_27_port, 
                           PLAINKEY(26) => PLAINKEY_26_port, PLAINKEY(25) => 
                           PLAINKEY_25_port, PLAINKEY(24) => PLAINKEY_24_port, 
                           PLAINKEY(23) => PLAINKEY_23_port, PLAINKEY(22) => 
                           PLAINKEY_22_port, PLAINKEY(21) => PLAINKEY_21_port, 
                           PLAINKEY(20) => PLAINKEY_20_port, PLAINKEY(19) => 
                           PLAINKEY_19_port, PLAINKEY(18) => PLAINKEY_18_port, 
                           PLAINKEY(17) => PLAINKEY_17_port, PLAINKEY(16) => 
                           PLAINKEY_16_port, PLAINKEY(15) => PLAINKEY_15_port, 
                           PLAINKEY(14) => PLAINKEY_14_port, PLAINKEY(13) => 
                           PLAINKEY_13_port, PLAINKEY(12) => PLAINKEY_12_port, 
                           PLAINKEY(11) => PLAINKEY_11_port, PLAINKEY(10) => 
                           PLAINKEY_10_port, PLAINKEY(9) => PLAINKEY_9_port, 
                           PLAINKEY(8) => PLAINKEY_8_port, PLAINKEY(7) => 
                           PLAINKEY_7_port, PLAINKEY(6) => PLAINKEY_6_port, 
                           PLAINKEY(5) => PLAINKEY_5_port, PLAINKEY(4) => 
                           PLAINKEY_4_port, PLAINKEY(3) => PLAINKEY_3_port, 
                           PLAINKEY(2) => PLAINKEY_2_port, PLAINKEY(1) => 
                           PLAINKEY_1_port, PLAINKEY(0) => PLAINKEY_0_port, 
                           RBUF_FULL => RBUF_FULL, PARITY_ERROR => PARITY_ERROR
                           );
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RMEDT_REWIRE_0 is

   port( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN : in std_logic;  DATA_IN : in 
         std_logic_vector (7 downto 0);  BS_ERROR, CRC_ERROR, EMPTY, FULL, 
         KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, R_ERROR, SENDING, 
         dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE : out std_logic;  DATA, 
         ADDR : out std_logic_vector (7 downto 0));

end RMEDT_REWIRE_0;

architecture SYN_struct of RMEDT_REWIRE_0 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component transmitter_block_0
      port( PRGA_OUT : in std_logic_vector (7 downto 0);  clk, p_ready : in 
            std_logic;  prga_opcode : in std_logic_vector (1 downto 0);  rst : 
            in std_logic;  SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE : out 
            std_logic);
   end component;
   
   component receiver_block_rewire_0
      port( CLK, DM1_RX, DP1_RX, RST : in std_logic;  BS_ERROR, CRC_ERROR, 
            EOP_external : out std_logic;  OPCODE : out std_logic_vector (1 
            downto 0);  RCV_DATA : out std_logic_vector (7 downto 0);  R_ERROR,
            W_ENABLE : out std_logic);
   end component;
   
   component memoryblock_0
      port( CLK, NEXT_BYTE : in std_logic;  RCV_DATA : in std_logic_vector (7 
            downto 0);  RCV_OPCODE : in std_logic_vector (1 downto 0);  RST, 
            W_ENABLE, EOP : in std_logic;  EMPTY, FULL, B_READY : out std_logic
            ;  PRGA_IN : out std_logic_vector (7 downto 0);  PRGA_OPCODE : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component EDBlock_0
      port( BYTE : in std_logic_vector (7 downto 0);  BYTE_READY, CLK : in 
            std_logic;  OPCODE : in std_logic_vector (1 downto 0);  RST, 
            SERIAL_IN : in std_logic;  DATA_IN : in std_logic_vector (7 downto 
            0);  KEY_ERROR, PARITY_ERROR, PDATA_READY : out std_logic;  
            PROCESSED_DATA : out std_logic_vector (7 downto 0);  PROG_ERROR, 
            RBUF_FULL, W_ENABLE, R_ENABLE : out std_logic;  DATA, ADDR : out 
            std_logic_vector (7 downto 0));
   end component;
   
   signal PRGA_IN_7_port, PRGA_IN_6_port, PRGA_IN_5_port, PRGA_IN_4_port, 
      PRGA_IN_3_port, PRGA_IN_2_port, PRGA_IN_1_port, PRGA_IN_0_port, B_READY, 
      PRGA_OPCODE_1_port, PRGA_OPCODE_0_port, PDATA_READY, 
      PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, PROCESSED_DATA_5_port, 
      PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, PROCESSED_DATA_2_port, 
      PROCESSED_DATA_1_port, PROCESSED_DATA_0_port, EOP_external, NEXT_BYTE, 
      RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      OPCODE_1_port, OPCODE_0_port, W_ENABLE, n1, n2 : std_logic;

begin
   
   U_0 : EDBlock_0 port map( BYTE(7) => PRGA_IN_7_port, BYTE(6) => 
                           PRGA_IN_6_port, BYTE(5) => PRGA_IN_5_port, BYTE(4) 
                           => PRGA_IN_4_port, BYTE(3) => PRGA_IN_3_port, 
                           BYTE(2) => PRGA_IN_2_port, BYTE(1) => PRGA_IN_1_port
                           , BYTE(0) => PRGA_IN_0_port, BYTE_READY => B_READY, 
                           CLK => CLK, OPCODE(1) => PRGA_OPCODE_1_port, 
                           OPCODE(0) => PRGA_OPCODE_0_port, RST => n1, 
                           SERIAL_IN => SERIAL_IN, DATA_IN(7) => DATA_IN(7), 
                           DATA_IN(6) => DATA_IN(6), DATA_IN(5) => DATA_IN(5), 
                           DATA_IN(4) => DATA_IN(4), DATA_IN(3) => DATA_IN(3), 
                           DATA_IN(2) => DATA_IN(2), DATA_IN(1) => DATA_IN(1), 
                           DATA_IN(0) => DATA_IN(0), KEY_ERROR => KEY_ERROR, 
                           PARITY_ERROR => PARITY_ERROR, PDATA_READY => 
                           PDATA_READY, PROCESSED_DATA(7) => 
                           PROCESSED_DATA_7_port, PROCESSED_DATA(6) => 
                           PROCESSED_DATA_6_port, PROCESSED_DATA(5) => 
                           PROCESSED_DATA_5_port, PROCESSED_DATA(4) => 
                           PROCESSED_DATA_4_port, PROCESSED_DATA(3) => 
                           PROCESSED_DATA_3_port, PROCESSED_DATA(2) => 
                           PROCESSED_DATA_2_port, PROCESSED_DATA(1) => 
                           PROCESSED_DATA_1_port, PROCESSED_DATA(0) => 
                           PROCESSED_DATA_0_port, PROG_ERROR => PROG_ERROR, 
                           RBUF_FULL => RBUF_FULL, W_ENABLE => W_ENABLE_R, 
                           R_ENABLE => R_ENABLE, DATA(7) => DATA(7), DATA(6) =>
                           DATA(6), DATA(5) => DATA(5), DATA(4) => DATA(4), 
                           DATA(3) => DATA(3), DATA(2) => DATA(2), DATA(1) => 
                           DATA(1), DATA(0) => DATA(0), ADDR(7) => ADDR(7), 
                           ADDR(6) => ADDR(6), ADDR(5) => ADDR(5), ADDR(4) => 
                           ADDR(4), ADDR(3) => ADDR(3), ADDR(2) => ADDR(2), 
                           ADDR(1) => ADDR(1), ADDR(0) => ADDR(0));
   U_1 : memoryblock_0 port map( CLK => CLK, NEXT_BYTE => NEXT_BYTE, 
                           RCV_DATA(7) => RCV_DATA_7_port, RCV_DATA(6) => 
                           RCV_DATA_6_port, RCV_DATA(5) => RCV_DATA_5_port, 
                           RCV_DATA(4) => RCV_DATA_4_port, RCV_DATA(3) => 
                           RCV_DATA_3_port, RCV_DATA(2) => RCV_DATA_2_port, 
                           RCV_DATA(1) => RCV_DATA_1_port, RCV_DATA(0) => 
                           RCV_DATA_0_port, RCV_OPCODE(1) => OPCODE_1_port, 
                           RCV_OPCODE(0) => OPCODE_0_port, RST => n1, W_ENABLE 
                           => W_ENABLE, EOP => EOP_external, EMPTY => EMPTY, 
                           FULL => FULL, B_READY => B_READY, PRGA_IN(7) => 
                           PRGA_IN_7_port, PRGA_IN(6) => PRGA_IN_6_port, 
                           PRGA_IN(5) => PRGA_IN_5_port, PRGA_IN(4) => 
                           PRGA_IN_4_port, PRGA_IN(3) => PRGA_IN_3_port, 
                           PRGA_IN(2) => PRGA_IN_2_port, PRGA_IN(1) => 
                           PRGA_IN_1_port, PRGA_IN(0) => PRGA_IN_0_port, 
                           PRGA_OPCODE(1) => PRGA_OPCODE_1_port, PRGA_OPCODE(0)
                           => PRGA_OPCODE_0_port);
   U_2 : receiver_block_rewire_0 port map( CLK => CLK, DM1_RX => DM1_RX, DP1_RX
                           => DP1_RX, RST => n1, BS_ERROR => BS_ERROR, 
                           CRC_ERROR => CRC_ERROR, EOP_external => EOP_external
                           , OPCODE(1) => OPCODE_1_port, OPCODE(0) => 
                           OPCODE_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, R_ERROR => R_ERROR, 
                           W_ENABLE => W_ENABLE);
   U_3 : transmitter_block_0 port map( PRGA_OUT(7) => PROCESSED_DATA_7_port, 
                           PRGA_OUT(6) => PROCESSED_DATA_6_port, PRGA_OUT(5) =>
                           PROCESSED_DATA_5_port, PRGA_OUT(4) => 
                           PROCESSED_DATA_4_port, PRGA_OUT(3) => 
                           PROCESSED_DATA_3_port, PRGA_OUT(2) => 
                           PROCESSED_DATA_2_port, PRGA_OUT(1) => 
                           PROCESSED_DATA_1_port, PRGA_OUT(0) => 
                           PROCESSED_DATA_0_port, clk => CLK, p_ready => 
                           PDATA_READY, prga_opcode(1) => PRGA_OPCODE_1_port, 
                           prga_opcode(0) => PRGA_OPCODE_0_port, rst => n1, 
                           SENDING => SENDING, dm_tx_out => dm_tx_out, 
                           dp_tx_out => dp_tx_out, NEXT_BYTE => NEXT_BYTE);
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_timer_1 is

   port( CLK, RST, TIMER_TRIG : in std_logic;  STOP_RCVING, SHIFT_STROBE : out 
         std_logic);

end uart_timer_1;

architecture SYN_timerB of uart_timer_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component uart_timer_1_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal state_7_port, state_6_port, state_5_port, state_4_port, state_3_port,
      state_2_port, state_1_port, state_0_port, nextState_7_port, 
      nextState_6_port, nextState_5_port, nextState_4_port, nextState_3_port, 
      nextState_2_port, nextState_1_port, nextState_0_port, N26, N27, N28, N29,
      N30, N31, N32, N33, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n1, n2, 
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26_port, n27_port, n28_port, n29_port
      , n30_port, n31_port, n32_port, n33_port, n34 : std_logic;

begin
   
   U21 : OR2X2 port map( A => state_7_port, B => n50, Y => n49);
   U38 : OAI21X1 port map( A => n20, B => n27_port, C => n35, Y => n64);
   U39 : NAND2X1 port map( A => N33, B => n36, Y => n35);
   U40 : OAI21X1 port map( A => n26_port, B => n20, C => n37, Y => n65);
   U41 : NAND2X1 port map( A => N32, B => n36, Y => n37);
   U42 : OAI21X1 port map( A => n25, B => n20, C => n38, Y => n66);
   U43 : NAND2X1 port map( A => N31, B => n36, Y => n38);
   U44 : OAI21X1 port map( A => n20, B => n24, C => n39, Y => n67);
   U45 : NAND2X1 port map( A => N30, B => n36, Y => n39);
   U46 : OAI21X1 port map( A => n23, B => n20, C => n40, Y => n68);
   U47 : NAND2X1 port map( A => N29, B => n36, Y => n40);
   U48 : OAI21X1 port map( A => n22, B => n20, C => n41, Y => n69);
   U49 : NAND2X1 port map( A => N28, B => n36, Y => n41);
   U50 : OAI21X1 port map( A => n20, B => n21, C => n42, Y => n70);
   U51 : NAND2X1 port map( A => N27, B => n36, Y => n42);
   U52 : OAI21X1 port map( A => n19, B => n20, C => n43, Y => n71);
   U53 : NAND2X1 port map( A => N26, B => n36, Y => n43);
   U54 : NOR2X1 port map( A => n44, B => n72, Y => n36);
   U55 : NOR2X1 port map( A => n72, B => TIMER_TRIG, Y => n44);
   U56 : NOR2X1 port map( A => n45, B => n46, Y => n72);
   U57 : NAND3X1 port map( A => nextState_6_port, B => nextState_5_port, C => 
                           n47, Y => n46);
   U58 : NOR2X1 port map( A => n22, B => n23, Y => n47);
   U59 : NAND3X1 port map( A => nextState_0_port, B => n21, C => n48, Y => n45)
                           ;
   U60 : NOR2X1 port map( A => nextState_7_port, B => nextState_4_port, Y => 
                           n48);
   U61 : NOR2X1 port map( A => state_0_port, B => n49, Y => SHIFT_STROBE);
   U62 : AOI21X1 port map( A => n51, B => n32_port, C => n52, Y => n50);
   U63 : OAI21X1 port map( A => n33_port, B => n53, C => n54, Y => n52);
   U64 : NAND3X1 port map( A => state_6_port, B => state_1_port, C => n55, Y =>
                           n54);
   U65 : AOI21X1 port map( A => n56, B => n57, C => state_3_port, Y => n55);
   U66 : NAND3X1 port map( A => n33_port, B => n31_port, C => state_4_port, Y 
                           => n57);
   U67 : NAND3X1 port map( A => state_2_port, B => n32_port, C => state_5_port,
                           Y => n56);
   U68 : NAND2X1 port map( A => state_4_port, B => n58, Y => n53);
   U69 : OAI21X1 port map( A => state_2_port, B => n28_port, C => n59, Y => n51
                           );
   U70 : NAND3X1 port map( A => state_2_port, B => n29_port, C => n30_port, Y 
                           => n59);
   U71 : OAI22X1 port map( A => state_6_port, B => n61, C => n29_port, D => n60
                           , Y => n58);
   U72 : NAND3X1 port map( A => n34, B => n31_port, C => state_3_port, Y => n60
                           );
   U73 : AOI22X1 port map( A => n62, B => state_1_port, C => n63, D => 
                           state_5_port, Y => n61);
   U74 : XOR2X1 port map( A => n34, B => state_3_port, Y => n63);
   U75 : NOR2X1 port map( A => state_5_port, B => state_3_port, Y => n62);
   add_39 : uart_timer_1_DW01_inc_0 port map( A(7) => nextState_7_port, A(6) =>
                           nextState_6_port, A(5) => nextState_5_port, A(4) => 
                           nextState_4_port, A(3) => nextState_3_port, A(2) => 
                           nextState_2_port, A(1) => nextState_1_port, A(0) => 
                           nextState_0_port, SUM(7) => N33, SUM(6) => N32, 
                           SUM(5) => N31, SUM(4) => N30, SUM(3) => N29, SUM(2) 
                           => N28, SUM(1) => N27, SUM(0) => N26);
   state_reg_3_inst : DFFSR port map( D => nextState_3_port, CLK => CLK, R => 
                           n18, S => n17, Q => state_3_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n18, S => n16, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n18, S => n15, Q => state_1_port);
   state_reg_5_inst : DFFSR port map( D => nextState_5_port, CLK => CLK, R => 
                           n18, S => n14, Q => state_5_port);
   state_reg_6_inst : DFFSR port map( D => nextState_6_port, CLK => CLK, R => 
                           n18, S => n13, Q => state_6_port);
   state_reg_4_inst : DFFSR port map( D => nextState_4_port, CLK => CLK, R => 
                           n18, S => n12, Q => state_4_port);
   state_reg_7_inst : DFFSR port map( D => nextState_7_port, CLK => CLK, R => 
                           n18, S => n11, Q => state_7_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n18, S => n10, Q => state_0_port);
   STOP_RCVING_reg : DFFSR port map( D => n72, CLK => CLK, R => n18, S => n9, Q
                           => STOP_RCVING);
   nextState_reg_3_inst : DFFSR port map( D => n68, CLK => CLK, R => n18, S => 
                           n8, Q => nextState_3_port);
   nextState_reg_2_inst : DFFSR port map( D => n69, CLK => CLK, R => n18, S => 
                           n7, Q => nextState_2_port);
   nextState_reg_0_inst : DFFSR port map( D => n71, CLK => CLK, R => n18, S => 
                           n6, Q => nextState_0_port);
   nextState_reg_4_inst : DFFSR port map( D => n67, CLK => CLK, R => n18, S => 
                           n5, Q => nextState_4_port);
   nextState_reg_1_inst : DFFSR port map( D => n70, CLK => CLK, R => n18, S => 
                           n4, Q => nextState_1_port);
   nextState_reg_5_inst : DFFSR port map( D => n66, CLK => CLK, R => n18, S => 
                           n3, Q => nextState_5_port);
   nextState_reg_6_inst : DFFSR port map( D => n65, CLK => CLK, R => n18, S => 
                           n2, Q => nextState_6_port);
   nextState_reg_7_inst : DFFSR port map( D => n64, CLK => CLK, R => n18, S => 
                           n1, Q => nextState_7_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   U20 : INVX2 port map( A => RST, Y => n18);
   U22 : INVX2 port map( A => nextState_0_port, Y => n19);
   U23 : INVX2 port map( A => n44, Y => n20);
   U24 : INVX2 port map( A => nextState_1_port, Y => n21);
   U25 : INVX2 port map( A => nextState_2_port, Y => n22);
   U26 : INVX2 port map( A => nextState_3_port, Y => n23);
   U27 : INVX2 port map( A => nextState_4_port, Y => n24);
   U28 : INVX2 port map( A => nextState_5_port, Y => n25);
   U29 : INVX2 port map( A => nextState_6_port, Y => n26_port);
   U30 : INVX2 port map( A => nextState_7_port, Y => n27_port);
   U31 : INVX2 port map( A => n58, Y => n28_port);
   U32 : INVX2 port map( A => state_6_port, Y => n29_port);
   U33 : INVX2 port map( A => n60, Y => n30_port);
   U34 : INVX2 port map( A => state_5_port, Y => n31_port);
   U35 : INVX2 port map( A => state_4_port, Y => n32_port);
   U36 : INVX2 port map( A => state_2_port, Y => n33_port);
   U37 : INVX2 port map( A => state_1_port, Y => n34);

end SYN_timerB;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity keyreg_1 is

   port( CLK, RST, SBE, OE, RBUF_FULL : in std_logic;  RCV_DATA : in 
         std_logic_vector (7 downto 0);  PLAINKEY : out std_logic_vector (63 
         downto 0);  KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR : out 
         std_logic);

end keyreg_1;

architecture SYN_keyb of keyreg_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component keyreg_1_DW01_add_0
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port, 
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port, CLR_RBUFF_port, state_3_port, state_2_port, state_1_port
      , state_0_port, parityError, keyCount_3_port, keyCount_2_port, 
      keyCount_1_port, keyCount_0_port, address_7_port, address_6_port, 
      address_5_port, address_4_port, address_3_port, address_2_port, 
      address_1_port, address_0_port, currentPlainKey_63_port, 
      currentPlainKey_62_port, currentPlainKey_61_port, currentPlainKey_60_port
      , currentPlainKey_59_port, currentPlainKey_58_port, 
      currentPlainKey_57_port, currentPlainKey_56_port, currentPlainKey_55_port
      , currentPlainKey_54_port, currentPlainKey_53_port, 
      currentPlainKey_52_port, currentPlainKey_51_port, currentPlainKey_50_port
      , currentPlainKey_49_port, currentPlainKey_48_port, 
      currentPlainKey_47_port, currentPlainKey_46_port, currentPlainKey_45_port
      , currentPlainKey_44_port, currentPlainKey_43_port, 
      currentPlainKey_42_port, currentPlainKey_41_port, currentPlainKey_40_port
      , currentPlainKey_39_port, currentPlainKey_38_port, 
      currentPlainKey_37_port, currentPlainKey_36_port, currentPlainKey_35_port
      , currentPlainKey_34_port, currentPlainKey_33_port, 
      currentPlainKey_32_port, currentPlainKey_31_port, currentPlainKey_30_port
      , currentPlainKey_29_port, currentPlainKey_28_port, 
      currentPlainKey_27_port, currentPlainKey_26_port, currentPlainKey_25_port
      , currentPlainKey_24_port, currentPlainKey_23_port, 
      currentPlainKey_22_port, currentPlainKey_21_port, currentPlainKey_20_port
      , currentPlainKey_19_port, currentPlainKey_18_port, 
      currentPlainKey_17_port, currentPlainKey_16_port, currentPlainKey_15_port
      , currentPlainKey_14_port, currentPlainKey_13_port, 
      currentPlainKey_12_port, currentPlainKey_11_port, currentPlainKey_10_port
      , currentPlainKey_9_port, currentPlainKey_8_port, currentPlainKey_7_port,
      currentPlainKey_6_port, currentPlainKey_5_port, currentPlainKey_4_port, 
      currentPlainKey_3_port, currentPlainKey_2_port, currentPlainKey_1_port, 
      currentPlainKey_0_port, parityAccumulator_7_port, 
      parityAccumulator_6_port, parityAccumulator_5_port, 
      parityAccumulator_4_port, parityAccumulator_3_port, 
      parityAccumulator_2_port, parityAccumulator_1_port, 
      parityAccumulator_0_port, nextParityError, N694, N1792, N1793, N1794, 
      N1795, N1796, N1797, N1798, N1799, n3, n12, n13, n15, n18, n22, n24, n26,
      n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56
      , n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, n80, n82, n84, 
      n86, n88, n90, n92, n94, n96, n98, n100, n102, n104, n106, n108, n110, 
      n112, n114, n116, n118, n120, n122, n124, n126, n128, n130, n132, n134, 
      n136, n138, n140, n142, n144, n146, n148, n152, n155, n157, n159, n162, 
      n163, n164, n167, n169, n170, n171, n174, n176, n179, n182, n190, n191, 
      n194, n196, n198, n199, n200, n201, n202, n204, n211, n212, n213, n214, 
      n215, n216, n218, n220, n235, n236, n237, n238, n239, n246, n251, n252, 
      n253, n254, n256, n272, n273, n274, n276, n283, n288, n290, n292, n293, 
      n294, n306, n307, n308, n309, n310, n318, n323, n325, n328, n329, n341, 
      n342, n349, n354, n356, n358, n359, n371, n372, n379, n384, n386, n388, 
      n389, n401, n402, n403, n410, n415, n417, n420, n421, n433, n434, n442, 
      n447, n449, n451, n463, n464, n470, n475, n477, n478, n490, n491, n497, 
      n502, n504, n505, n517, n518, n524, n529, n531, n532, n544, n545, n546, 
      n553, n558, n560, n562, n574, n575, n581, n586, n588, n589, n601, n602, 
      n608, n613, n615, n616, n628, n629, n635, n640, n642, n643, n655, n656, 
      n664, n669, n671, n673, n685, n686, n692, n697, n699, n700, n712, n713, 
      n719, n724, n726, n727, n739, n740, n746, n751, n753, n754, n766, n767, 
      n768, n775, n780, n782, n784, n796, n797, n803, n808, n810, n811, n823, 
      n824, n830, n835, n837, n838, n850, n851, n857, n862, n864, n865, n877, 
      n878, n886, n891, n893, n895, n907, n908, n914, n919, n921, n922, n934, 
      n935, n941, n946, n948, n949, n961, n962, n968, n973, n975, n976, n988, 
      n989, n990, n1002, n1004, n1006, n1011, n1018, n1019, n1031, n1033, n1034
      , n1038, n1046, n1047, n1062, n1063, n1077, n1078, n1089, n1090, n1101, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1143, n1144, n1160, n1178, 
      n1186, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, 
      n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
      n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, 
      n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
      n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1269, n1270, n1271, n1272, n1273, 
      n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
      n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, 
      n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, 
      n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, 
      n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, 
      n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, 
      n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, 
      n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, 
      n1354, n1355, n1356, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n14, n16, 
      n17, n19, n20, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, n41, n43
      , n45, n47, n49, n51, n53, n55, n57, n59, n61, n63, n65, n67, n69, n71, 
      n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95, n97, n99, 
      n101, n103, n105, n107, n109, n111, n113, n115, n117, n119, n121, n123, 
      n125, n127, n129, n131, n133, n135, n137, n139, n141, n143, n145, n147, 
      n149, n150, n151, n153, n154, n156, n158, n160, n161, n165, n166, n168, 
      n172, n173, n175, n177, n178, n180, n181, n183, n184, n185, n186, n187, 
      n188, n189, n192, n193, n195, n197, n203, n205, n206, n207, n208, n209, 
      n210, n217, n219, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n240, n241, n242, n243, n244, n245, n247, 
      n248, n249, n250, n255, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n275, n277, n278, n279, n280, 
      n281, n282, n284, n285, n286, n287, n289, n291, n295, n296, n297, n298, 
      n299, n300, n301, n302, n303, n304, n305, n311, n312, n313, n314, n315, 
      n316, n317, n319, n320, n321, n322, n324, n326, n327, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n343, n344, n345, n346, 
      n347, n348, n350, n351, n352, n353, n355, n357, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n373, n374, n375, n376, n377, 
      n378, n380, n381, n382, n383, n385, n387, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n404, n405, n406, n407, n408, n409, 
      n411, n412, n413, n414, n416, n418, n419, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n435, n436, n437, n438, n439, n440, 
      n441, n443, n444, n445, n446, n448, n450, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n465, n466, n467, n468, n469, n471, 
      n472, n473, n474, n476, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n492, n493, n494, n495, n496, n498, n499, n500, n501, 
      n503, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n519, n520, n521, n522, n523, n525, n526, n527, n528, n530, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n547, n548, n549, 
      n550, n551, n552, n554, n555, n556, n557, n559, n561, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n576, n577, n578, n579, 
      n580, n582, n583, n584, n585, n587, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n603, n604, n605, n606, n607, n609, n610, 
      n611, n612, n614, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n630, n631, n632, n633, n634, n636, n637, n638, n639, n641, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n657, 
      n658, n659, n660, n661, n662, n663, n665, n666, n667, n668, n670, n672, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n687, 
      n688, n689, n690, n691, n693, n694_port, n695, n696, n698, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n714, n715, n716, 
      n717, n718, n720, n721, n722, n723, n725, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n741, n742, n743, n744, n745, n747, 
      n748, n749, n750, n752, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n769, n770, n771, n772, n773, n774, n776, n777, n778, 
      n779, n781, n783, n785, n786, n787, n788, n789, n790, n791, n792, n793, 
      n794, n795, n798, n799, n800, n801, n802, n804, n805, n806, n807, n809, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n825, 
      n826, n827, n828, n829, n831, n832, n833, n834, n836, n839, n840, n841, 
      n842, n843, n844, n845, n846, n847, n848, n849, n852, n853, n854, n855, 
      n856, n858, n859, n860, n861, n863, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n879, n880, n881, n882, n883, n884, n885, 
      n887, n888, n889, n890, n892, n894, n896, n897, n898, n899, n900, n901, 
      n902, n903, n904, n905, n906, n909, n910, n911, n912, n913, n915, n916, 
      n917, n918, n920, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n936, n937, n938, n939, n940, n942, n943, n944, n945, n947, 
      n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n963, 
      n964, n965, n966, n967, n969, n970, n971, n972, n974, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n991, n992, n993, n994, 
      n995, n996, n997, n998, n999, n1000, n1001, n1003, n1005, n1007, n1008, 
      n1009, n1010, n1012, n1013, n1014, n1015, n1016, n1017, n1020, n1021, 
      n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1032, 
      n1035, n1036, n1037, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1079, n1080, n1081, 
      n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1102, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1179, n1180, n1181, n1182, n1183, n1184, 
      n1185, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, 
      n1196, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1357, 
      n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
      n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, 
      n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, PROG_ERROR_port, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n_1025 : std_logic;

begin
   PLAINKEY <= ( PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port, 
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port );
   PROG_ERROR <= PROG_ERROR_port;
   CLR_RBUFF <= CLR_RBUFF_port;
   
   n3 <= '0';
   keyCount_reg_0_inst : DFFPOSX1 port map( D => n1356, CLK => CLK, Q => 
                           keyCount_0_port);
   keyCount_reg_2_inst : DFFPOSX1 port map( D => n1349, CLK => CLK, Q => 
                           keyCount_2_port);
   keyCount_reg_3_inst : DFFPOSX1 port map( D => n1355, CLK => CLK, Q => 
                           keyCount_3_port);
   parityAccumulator_reg_0_inst : DFFPOSX1 port map( D => n1348, CLK => CLK, Q 
                           => parityAccumulator_0_port);
   parityAccumulator_reg_1_inst : DFFPOSX1 port map( D => n1347, CLK => CLK, Q 
                           => parityAccumulator_1_port);
   parityAccumulator_reg_2_inst : DFFPOSX1 port map( D => n1346, CLK => CLK, Q 
                           => parityAccumulator_2_port);
   parityAccumulator_reg_3_inst : DFFPOSX1 port map( D => n1345, CLK => CLK, Q 
                           => parityAccumulator_3_port);
   parityAccumulator_reg_4_inst : DFFPOSX1 port map( D => n1344, CLK => CLK, Q 
                           => parityAccumulator_4_port);
   parityAccumulator_reg_5_inst : DFFPOSX1 port map( D => n1343, CLK => CLK, Q 
                           => parityAccumulator_5_port);
   parityAccumulator_reg_6_inst : DFFPOSX1 port map( D => n1342, CLK => CLK, Q 
                           => parityAccumulator_6_port);
   parityAccumulator_reg_7_inst : DFFPOSX1 port map( D => n1341, CLK => CLK, Q 
                           => parityAccumulator_7_port);
   keyCount_reg_1_inst : DFFPOSX1 port map( D => n1350, CLK => CLK, Q => 
                           keyCount_1_port);
   address_reg_7_inst : DFFPOSX1 port map( D => n1340, CLK => CLK, Q => 
                           address_7_port);
   address_reg_6_inst : DFFPOSX1 port map( D => n1339, CLK => CLK, Q => 
                           address_6_port);
   address_reg_5_inst : DFFPOSX1 port map( D => n1338, CLK => CLK, Q => 
                           address_5_port);
   address_reg_4_inst : DFFPOSX1 port map( D => n1337, CLK => CLK, Q => 
                           address_4_port);
   address_reg_3_inst : DFFPOSX1 port map( D => n1336, CLK => CLK, Q => 
                           address_3_port);
   address_reg_2_inst : DFFPOSX1 port map( D => n1335, CLK => CLK, Q => 
                           address_2_port);
   address_reg_1_inst : DFFPOSX1 port map( D => n1334, CLK => CLK, Q => 
                           address_1_port);
   address_reg_0_inst : DFFPOSX1 port map( D => n1333, CLK => CLK, Q => 
                           address_0_port);
   currentPlainKey_reg_63_inst : DFFPOSX1 port map( D => n1269, CLK => CLK, Q 
                           => currentPlainKey_63_port);
   currentPlainKey_reg_62_inst : DFFPOSX1 port map( D => n1270, CLK => CLK, Q 
                           => currentPlainKey_62_port);
   currentPlainKey_reg_61_inst : DFFPOSX1 port map( D => n1271, CLK => CLK, Q 
                           => currentPlainKey_61_port);
   currentPlainKey_reg_60_inst : DFFPOSX1 port map( D => n1272, CLK => CLK, Q 
                           => currentPlainKey_60_port);
   currentPlainKey_reg_59_inst : DFFPOSX1 port map( D => n1273, CLK => CLK, Q 
                           => currentPlainKey_59_port);
   currentPlainKey_reg_58_inst : DFFPOSX1 port map( D => n1274, CLK => CLK, Q 
                           => currentPlainKey_58_port);
   currentPlainKey_reg_57_inst : DFFPOSX1 port map( D => n1275, CLK => CLK, Q 
                           => currentPlainKey_57_port);
   currentPlainKey_reg_56_inst : DFFPOSX1 port map( D => n1276, CLK => CLK, Q 
                           => currentPlainKey_56_port);
   currentPlainKey_reg_55_inst : DFFPOSX1 port map( D => n1277, CLK => CLK, Q 
                           => currentPlainKey_55_port);
   currentPlainKey_reg_54_inst : DFFPOSX1 port map( D => n1278, CLK => CLK, Q 
                           => currentPlainKey_54_port);
   currentPlainKey_reg_53_inst : DFFPOSX1 port map( D => n1279, CLK => CLK, Q 
                           => currentPlainKey_53_port);
   currentPlainKey_reg_52_inst : DFFPOSX1 port map( D => n1280, CLK => CLK, Q 
                           => currentPlainKey_52_port);
   currentPlainKey_reg_51_inst : DFFPOSX1 port map( D => n1281, CLK => CLK, Q 
                           => currentPlainKey_51_port);
   currentPlainKey_reg_50_inst : DFFPOSX1 port map( D => n1282, CLK => CLK, Q 
                           => currentPlainKey_50_port);
   currentPlainKey_reg_49_inst : DFFPOSX1 port map( D => n1283, CLK => CLK, Q 
                           => currentPlainKey_49_port);
   currentPlainKey_reg_48_inst : DFFPOSX1 port map( D => n1284, CLK => CLK, Q 
                           => currentPlainKey_48_port);
   currentPlainKey_reg_47_inst : DFFPOSX1 port map( D => n1285, CLK => CLK, Q 
                           => currentPlainKey_47_port);
   currentPlainKey_reg_46_inst : DFFPOSX1 port map( D => n1286, CLK => CLK, Q 
                           => currentPlainKey_46_port);
   currentPlainKey_reg_45_inst : DFFPOSX1 port map( D => n1287, CLK => CLK, Q 
                           => currentPlainKey_45_port);
   currentPlainKey_reg_44_inst : DFFPOSX1 port map( D => n1288, CLK => CLK, Q 
                           => currentPlainKey_44_port);
   currentPlainKey_reg_43_inst : DFFPOSX1 port map( D => n1289, CLK => CLK, Q 
                           => currentPlainKey_43_port);
   currentPlainKey_reg_42_inst : DFFPOSX1 port map( D => n1290, CLK => CLK, Q 
                           => currentPlainKey_42_port);
   currentPlainKey_reg_41_inst : DFFPOSX1 port map( D => n1291, CLK => CLK, Q 
                           => currentPlainKey_41_port);
   currentPlainKey_reg_40_inst : DFFPOSX1 port map( D => n1292, CLK => CLK, Q 
                           => currentPlainKey_40_port);
   currentPlainKey_reg_39_inst : DFFPOSX1 port map( D => n1293, CLK => CLK, Q 
                           => currentPlainKey_39_port);
   currentPlainKey_reg_38_inst : DFFPOSX1 port map( D => n1294, CLK => CLK, Q 
                           => currentPlainKey_38_port);
   currentPlainKey_reg_37_inst : DFFPOSX1 port map( D => n1295, CLK => CLK, Q 
                           => currentPlainKey_37_port);
   currentPlainKey_reg_36_inst : DFFPOSX1 port map( D => n1296, CLK => CLK, Q 
                           => currentPlainKey_36_port);
   currentPlainKey_reg_35_inst : DFFPOSX1 port map( D => n1297, CLK => CLK, Q 
                           => currentPlainKey_35_port);
   currentPlainKey_reg_34_inst : DFFPOSX1 port map( D => n1298, CLK => CLK, Q 
                           => currentPlainKey_34_port);
   currentPlainKey_reg_33_inst : DFFPOSX1 port map( D => n1299, CLK => CLK, Q 
                           => currentPlainKey_33_port);
   currentPlainKey_reg_32_inst : DFFPOSX1 port map( D => n1300, CLK => CLK, Q 
                           => currentPlainKey_32_port);
   currentPlainKey_reg_31_inst : DFFPOSX1 port map( D => n1301, CLK => CLK, Q 
                           => currentPlainKey_31_port);
   currentPlainKey_reg_30_inst : DFFPOSX1 port map( D => n1302, CLK => CLK, Q 
                           => currentPlainKey_30_port);
   currentPlainKey_reg_29_inst : DFFPOSX1 port map( D => n1303, CLK => CLK, Q 
                           => currentPlainKey_29_port);
   currentPlainKey_reg_28_inst : DFFPOSX1 port map( D => n1304, CLK => CLK, Q 
                           => currentPlainKey_28_port);
   currentPlainKey_reg_27_inst : DFFPOSX1 port map( D => n1305, CLK => CLK, Q 
                           => currentPlainKey_27_port);
   currentPlainKey_reg_26_inst : DFFPOSX1 port map( D => n1306, CLK => CLK, Q 
                           => currentPlainKey_26_port);
   currentPlainKey_reg_25_inst : DFFPOSX1 port map( D => n1307, CLK => CLK, Q 
                           => currentPlainKey_25_port);
   currentPlainKey_reg_24_inst : DFFPOSX1 port map( D => n1308, CLK => CLK, Q 
                           => currentPlainKey_24_port);
   currentPlainKey_reg_23_inst : DFFPOSX1 port map( D => n1309, CLK => CLK, Q 
                           => currentPlainKey_23_port);
   currentPlainKey_reg_22_inst : DFFPOSX1 port map( D => n1310, CLK => CLK, Q 
                           => currentPlainKey_22_port);
   currentPlainKey_reg_21_inst : DFFPOSX1 port map( D => n1311, CLK => CLK, Q 
                           => currentPlainKey_21_port);
   currentPlainKey_reg_20_inst : DFFPOSX1 port map( D => n1312, CLK => CLK, Q 
                           => currentPlainKey_20_port);
   currentPlainKey_reg_19_inst : DFFPOSX1 port map( D => n1313, CLK => CLK, Q 
                           => currentPlainKey_19_port);
   currentPlainKey_reg_18_inst : DFFPOSX1 port map( D => n1314, CLK => CLK, Q 
                           => currentPlainKey_18_port);
   currentPlainKey_reg_17_inst : DFFPOSX1 port map( D => n1315, CLK => CLK, Q 
                           => currentPlainKey_17_port);
   currentPlainKey_reg_16_inst : DFFPOSX1 port map( D => n1316, CLK => CLK, Q 
                           => currentPlainKey_16_port);
   currentPlainKey_reg_15_inst : DFFPOSX1 port map( D => n1317, CLK => CLK, Q 
                           => currentPlainKey_15_port);
   currentPlainKey_reg_14_inst : DFFPOSX1 port map( D => n1318, CLK => CLK, Q 
                           => currentPlainKey_14_port);
   currentPlainKey_reg_13_inst : DFFPOSX1 port map( D => n1319, CLK => CLK, Q 
                           => currentPlainKey_13_port);
   currentPlainKey_reg_12_inst : DFFPOSX1 port map( D => n1320, CLK => CLK, Q 
                           => currentPlainKey_12_port);
   currentPlainKey_reg_11_inst : DFFPOSX1 port map( D => n1321, CLK => CLK, Q 
                           => currentPlainKey_11_port);
   currentPlainKey_reg_10_inst : DFFPOSX1 port map( D => n1322, CLK => CLK, Q 
                           => currentPlainKey_10_port);
   currentPlainKey_reg_9_inst : DFFPOSX1 port map( D => n1323, CLK => CLK, Q =>
                           currentPlainKey_9_port);
   currentPlainKey_reg_8_inst : DFFPOSX1 port map( D => n1324, CLK => CLK, Q =>
                           currentPlainKey_8_port);
   currentPlainKey_reg_7_inst : DFFPOSX1 port map( D => n1325, CLK => CLK, Q =>
                           currentPlainKey_7_port);
   currentPlainKey_reg_6_inst : DFFPOSX1 port map( D => n1326, CLK => CLK, Q =>
                           currentPlainKey_6_port);
   currentPlainKey_reg_5_inst : DFFPOSX1 port map( D => n1327, CLK => CLK, Q =>
                           currentPlainKey_5_port);
   currentPlainKey_reg_4_inst : DFFPOSX1 port map( D => n1328, CLK => CLK, Q =>
                           currentPlainKey_4_port);
   currentPlainKey_reg_3_inst : DFFPOSX1 port map( D => n1329, CLK => CLK, Q =>
                           currentPlainKey_3_port);
   currentPlainKey_reg_2_inst : DFFPOSX1 port map( D => n1330, CLK => CLK, Q =>
                           currentPlainKey_2_port);
   currentPlainKey_reg_1_inst : DFFPOSX1 port map( D => n1331, CLK => CLK, Q =>
                           currentPlainKey_1_port);
   currentPlainKey_reg_0_inst : DFFPOSX1 port map( D => n1332, CLK => CLK, Q =>
                           currentPlainKey_0_port);
   PLAINKEY_reg_63_inst : DFFPOSX1 port map( D => n1260, CLK => CLK, Q => 
                           PLAINKEY_63_port);
   PLAINKEY_reg_62_inst : DFFPOSX1 port map( D => n1259, CLK => CLK, Q => 
                           PLAINKEY_62_port);
   PLAINKEY_reg_61_inst : DFFPOSX1 port map( D => n1258, CLK => CLK, Q => 
                           PLAINKEY_61_port);
   PLAINKEY_reg_60_inst : DFFPOSX1 port map( D => n1257, CLK => CLK, Q => 
                           PLAINKEY_60_port);
   PLAINKEY_reg_59_inst : DFFPOSX1 port map( D => n1256, CLK => CLK, Q => 
                           PLAINKEY_59_port);
   PLAINKEY_reg_58_inst : DFFPOSX1 port map( D => n1255, CLK => CLK, Q => 
                           PLAINKEY_58_port);
   PLAINKEY_reg_57_inst : DFFPOSX1 port map( D => n1254, CLK => CLK, Q => 
                           PLAINKEY_57_port);
   PLAINKEY_reg_56_inst : DFFPOSX1 port map( D => n1253, CLK => CLK, Q => 
                           PLAINKEY_56_port);
   PLAINKEY_reg_55_inst : DFFPOSX1 port map( D => n1252, CLK => CLK, Q => 
                           PLAINKEY_55_port);
   PLAINKEY_reg_54_inst : DFFPOSX1 port map( D => n1251, CLK => CLK, Q => 
                           PLAINKEY_54_port);
   PLAINKEY_reg_53_inst : DFFPOSX1 port map( D => n1250, CLK => CLK, Q => 
                           PLAINKEY_53_port);
   PLAINKEY_reg_52_inst : DFFPOSX1 port map( D => n1249, CLK => CLK, Q => 
                           PLAINKEY_52_port);
   PLAINKEY_reg_51_inst : DFFPOSX1 port map( D => n1248, CLK => CLK, Q => 
                           PLAINKEY_51_port);
   PLAINKEY_reg_50_inst : DFFPOSX1 port map( D => n1247, CLK => CLK, Q => 
                           PLAINKEY_50_port);
   PLAINKEY_reg_49_inst : DFFPOSX1 port map( D => n1246, CLK => CLK, Q => 
                           PLAINKEY_49_port);
   PLAINKEY_reg_48_inst : DFFPOSX1 port map( D => n1245, CLK => CLK, Q => 
                           PLAINKEY_48_port);
   PLAINKEY_reg_47_inst : DFFPOSX1 port map( D => n1244, CLK => CLK, Q => 
                           PLAINKEY_47_port);
   PLAINKEY_reg_46_inst : DFFPOSX1 port map( D => n1243, CLK => CLK, Q => 
                           PLAINKEY_46_port);
   PLAINKEY_reg_45_inst : DFFPOSX1 port map( D => n1242, CLK => CLK, Q => 
                           PLAINKEY_45_port);
   PLAINKEY_reg_44_inst : DFFPOSX1 port map( D => n1241, CLK => CLK, Q => 
                           PLAINKEY_44_port);
   PLAINKEY_reg_43_inst : DFFPOSX1 port map( D => n1240, CLK => CLK, Q => 
                           PLAINKEY_43_port);
   PLAINKEY_reg_42_inst : DFFPOSX1 port map( D => n1239, CLK => CLK, Q => 
                           PLAINKEY_42_port);
   PLAINKEY_reg_41_inst : DFFPOSX1 port map( D => n1238, CLK => CLK, Q => 
                           PLAINKEY_41_port);
   PLAINKEY_reg_40_inst : DFFPOSX1 port map( D => n1237, CLK => CLK, Q => 
                           PLAINKEY_40_port);
   PLAINKEY_reg_39_inst : DFFPOSX1 port map( D => n1236, CLK => CLK, Q => 
                           PLAINKEY_39_port);
   PLAINKEY_reg_38_inst : DFFPOSX1 port map( D => n1235, CLK => CLK, Q => 
                           PLAINKEY_38_port);
   PLAINKEY_reg_37_inst : DFFPOSX1 port map( D => n1234, CLK => CLK, Q => 
                           PLAINKEY_37_port);
   PLAINKEY_reg_36_inst : DFFPOSX1 port map( D => n1233, CLK => CLK, Q => 
                           PLAINKEY_36_port);
   PLAINKEY_reg_35_inst : DFFPOSX1 port map( D => n1232, CLK => CLK, Q => 
                           PLAINKEY_35_port);
   PLAINKEY_reg_34_inst : DFFPOSX1 port map( D => n1231, CLK => CLK, Q => 
                           PLAINKEY_34_port);
   PLAINKEY_reg_33_inst : DFFPOSX1 port map( D => n1230, CLK => CLK, Q => 
                           PLAINKEY_33_port);
   PLAINKEY_reg_32_inst : DFFPOSX1 port map( D => n1229, CLK => CLK, Q => 
                           PLAINKEY_32_port);
   PLAINKEY_reg_31_inst : DFFPOSX1 port map( D => n1228, CLK => CLK, Q => 
                           PLAINKEY_31_port);
   PLAINKEY_reg_30_inst : DFFPOSX1 port map( D => n1227, CLK => CLK, Q => 
                           PLAINKEY_30_port);
   PLAINKEY_reg_29_inst : DFFPOSX1 port map( D => n1226, CLK => CLK, Q => 
                           PLAINKEY_29_port);
   PLAINKEY_reg_28_inst : DFFPOSX1 port map( D => n1225, CLK => CLK, Q => 
                           PLAINKEY_28_port);
   PLAINKEY_reg_27_inst : DFFPOSX1 port map( D => n1224, CLK => CLK, Q => 
                           PLAINKEY_27_port);
   PLAINKEY_reg_26_inst : DFFPOSX1 port map( D => n1223, CLK => CLK, Q => 
                           PLAINKEY_26_port);
   PLAINKEY_reg_25_inst : DFFPOSX1 port map( D => n1222, CLK => CLK, Q => 
                           PLAINKEY_25_port);
   PLAINKEY_reg_24_inst : DFFPOSX1 port map( D => n1221, CLK => CLK, Q => 
                           PLAINKEY_24_port);
   PLAINKEY_reg_23_inst : DFFPOSX1 port map( D => n1220, CLK => CLK, Q => 
                           PLAINKEY_23_port);
   PLAINKEY_reg_22_inst : DFFPOSX1 port map( D => n1219, CLK => CLK, Q => 
                           PLAINKEY_22_port);
   PLAINKEY_reg_21_inst : DFFPOSX1 port map( D => n1218, CLK => CLK, Q => 
                           PLAINKEY_21_port);
   PLAINKEY_reg_20_inst : DFFPOSX1 port map( D => n1217, CLK => CLK, Q => 
                           PLAINKEY_20_port);
   PLAINKEY_reg_19_inst : DFFPOSX1 port map( D => n1216, CLK => CLK, Q => 
                           PLAINKEY_19_port);
   PLAINKEY_reg_18_inst : DFFPOSX1 port map( D => n1215, CLK => CLK, Q => 
                           PLAINKEY_18_port);
   PLAINKEY_reg_17_inst : DFFPOSX1 port map( D => n1214, CLK => CLK, Q => 
                           PLAINKEY_17_port);
   PLAINKEY_reg_16_inst : DFFPOSX1 port map( D => n1213, CLK => CLK, Q => 
                           PLAINKEY_16_port);
   PLAINKEY_reg_15_inst : DFFPOSX1 port map( D => n1212, CLK => CLK, Q => 
                           PLAINKEY_15_port);
   PLAINKEY_reg_14_inst : DFFPOSX1 port map( D => n1211, CLK => CLK, Q => 
                           PLAINKEY_14_port);
   PLAINKEY_reg_13_inst : DFFPOSX1 port map( D => n1210, CLK => CLK, Q => 
                           PLAINKEY_13_port);
   PLAINKEY_reg_12_inst : DFFPOSX1 port map( D => n1209, CLK => CLK, Q => 
                           PLAINKEY_12_port);
   PLAINKEY_reg_11_inst : DFFPOSX1 port map( D => n1208, CLK => CLK, Q => 
                           PLAINKEY_11_port);
   PLAINKEY_reg_10_inst : DFFPOSX1 port map( D => n1207, CLK => CLK, Q => 
                           PLAINKEY_10_port);
   PLAINKEY_reg_9_inst : DFFPOSX1 port map( D => n1206, CLK => CLK, Q => 
                           PLAINKEY_9_port);
   PLAINKEY_reg_8_inst : DFFPOSX1 port map( D => n1205, CLK => CLK, Q => 
                           PLAINKEY_8_port);
   PLAINKEY_reg_7_inst : DFFPOSX1 port map( D => n1204, CLK => CLK, Q => 
                           PLAINKEY_7_port);
   PLAINKEY_reg_6_inst : DFFPOSX1 port map( D => n1203, CLK => CLK, Q => 
                           PLAINKEY_6_port);
   PLAINKEY_reg_5_inst : DFFPOSX1 port map( D => n1202, CLK => CLK, Q => 
                           PLAINKEY_5_port);
   PLAINKEY_reg_4_inst : DFFPOSX1 port map( D => n1201, CLK => CLK, Q => 
                           PLAINKEY_4_port);
   PLAINKEY_reg_3_inst : DFFPOSX1 port map( D => n1200, CLK => CLK, Q => 
                           PLAINKEY_3_port);
   PLAINKEY_reg_2_inst : DFFPOSX1 port map( D => n1199, CLK => CLK, Q => 
                           PLAINKEY_2_port);
   PLAINKEY_reg_1_inst : DFFPOSX1 port map( D => n1198, CLK => CLK, Q => 
                           PLAINKEY_1_port);
   PLAINKEY_reg_0_inst : DFFPOSX1 port map( D => n1197, CLK => CLK, Q => 
                           PLAINKEY_0_port);
   U9 : NAND3X1 port map( A => parityAccumulator_7_port, B => 
                           parityAccumulator_6_port, C => n15, Y => n13);
   U10 : NOR2X1 port map( A => n1490, B => n1491, Y => n15);
   U11 : NAND3X1 port map( A => parityAccumulator_3_port, B => 
                           parityAccumulator_2_port, C => n18, Y => n12);
   U12 : NOR2X1 port map( A => n1486, B => n1487, Y => n18);
   U13 : OAI21X1 port map( A => n227, B => n1573, C => n22, Y => n1197);
   U14 : NAND2X1 port map( A => PLAINKEY_0_port, B => n231, Y => n22);
   U15 : OAI21X1 port map( A => n227, B => n1572, C => n24, Y => n1198);
   U16 : NAND2X1 port map( A => PLAINKEY_1_port, B => RST, Y => n24);
   U17 : OAI21X1 port map( A => n227, B => n1571, C => n26, Y => n1199);
   U18 : NAND2X1 port map( A => PLAINKEY_2_port, B => RST, Y => n26);
   U19 : OAI21X1 port map( A => n227, B => n1570, C => n28, Y => n1200);
   U20 : NAND2X1 port map( A => PLAINKEY_3_port, B => RST, Y => n28);
   U21 : OAI21X1 port map( A => n227, B => n1569, C => n30, Y => n1201);
   U22 : NAND2X1 port map( A => PLAINKEY_4_port, B => n231, Y => n30);
   U24 : OAI21X1 port map( A => n227, B => n1568, C => n32, Y => n1202);
   U25 : NAND2X1 port map( A => PLAINKEY_5_port, B => n232, Y => n32);
   U27 : OAI21X1 port map( A => n227, B => n1567, C => n34, Y => n1203);
   U28 : NAND2X1 port map( A => PLAINKEY_6_port, B => n233, Y => n34);
   U30 : OAI21X1 port map( A => n227, B => n1566, C => n36, Y => n1204);
   U31 : NAND2X1 port map( A => PLAINKEY_7_port, B => RST, Y => n36);
   U33 : OAI21X1 port map( A => n227, B => n1565, C => n38, Y => n1205);
   U34 : NAND2X1 port map( A => PLAINKEY_8_port, B => n231, Y => n38);
   U36 : OAI21X1 port map( A => n228, B => n1564, C => n40, Y => n1206);
   U37 : NAND2X1 port map( A => PLAINKEY_9_port, B => n232, Y => n40);
   U39 : OAI21X1 port map( A => n228, B => n1563, C => n42, Y => n1207);
   U40 : NAND2X1 port map( A => PLAINKEY_10_port, B => n233, Y => n42);
   U42 : OAI21X1 port map( A => n228, B => n1562, C => n44, Y => n1208);
   U43 : NAND2X1 port map( A => PLAINKEY_11_port, B => n233, Y => n44);
   U45 : OAI21X1 port map( A => n228, B => n1561, C => n46, Y => n1209);
   U46 : NAND2X1 port map( A => PLAINKEY_12_port, B => n233, Y => n46);
   U48 : OAI21X1 port map( A => n228, B => n1560, C => n48, Y => n1210);
   U49 : NAND2X1 port map( A => PLAINKEY_13_port, B => n233, Y => n48);
   U51 : OAI21X1 port map( A => n228, B => n1559, C => n50, Y => n1211);
   U52 : NAND2X1 port map( A => PLAINKEY_14_port, B => n233, Y => n50);
   U54 : OAI21X1 port map( A => n228, B => n1558, C => n52, Y => n1212);
   U55 : NAND2X1 port map( A => PLAINKEY_15_port, B => n233, Y => n52);
   U57 : OAI21X1 port map( A => n229, B => n1557, C => n54, Y => n1213);
   U58 : NAND2X1 port map( A => PLAINKEY_16_port, B => n233, Y => n54);
   U60 : OAI21X1 port map( A => n229, B => n1556, C => n56, Y => n1214);
   U61 : NAND2X1 port map( A => PLAINKEY_17_port, B => n233, Y => n56);
   U63 : OAI21X1 port map( A => n229, B => n1555, C => n58, Y => n1215);
   U64 : NAND2X1 port map( A => PLAINKEY_18_port, B => n233, Y => n58);
   U66 : OAI21X1 port map( A => n229, B => n1554, C => n60, Y => n1216);
   U67 : NAND2X1 port map( A => PLAINKEY_19_port, B => n233, Y => n60);
   U69 : OAI21X1 port map( A => n229, B => n1553, C => n62, Y => n1217);
   U70 : NAND2X1 port map( A => PLAINKEY_20_port, B => n233, Y => n62);
   U72 : OAI21X1 port map( A => n229, B => n1552, C => n64, Y => n1218);
   U73 : NAND2X1 port map( A => PLAINKEY_21_port, B => n233, Y => n64);
   U75 : OAI21X1 port map( A => n229, B => n1551, C => n66, Y => n1219);
   U76 : NAND2X1 port map( A => PLAINKEY_22_port, B => n233, Y => n66);
   U78 : OAI21X1 port map( A => n230, B => n1550, C => n68, Y => n1220);
   U79 : NAND2X1 port map( A => PLAINKEY_23_port, B => n233, Y => n68);
   U81 : OAI21X1 port map( A => n229, B => n1549, C => n70, Y => n1221);
   U82 : NAND2X1 port map( A => PLAINKEY_24_port, B => n233, Y => n70);
   U84 : OAI21X1 port map( A => n228, B => n1548, C => n72, Y => n1222);
   U85 : NAND2X1 port map( A => PLAINKEY_25_port, B => n233, Y => n72);
   U87 : OAI21X1 port map( A => n230, B => n1547, C => n74, Y => n1223);
   U88 : NAND2X1 port map( A => PLAINKEY_26_port, B => n233, Y => n74);
   U90 : OAI21X1 port map( A => n230, B => n1546, C => n76, Y => n1224);
   U91 : NAND2X1 port map( A => PLAINKEY_27_port, B => n233, Y => n76);
   U93 : OAI21X1 port map( A => n229, B => n1545, C => n78, Y => n1225);
   U94 : NAND2X1 port map( A => PLAINKEY_28_port, B => n233, Y => n78);
   U96 : OAI21X1 port map( A => n230, B => n1544, C => n80, Y => n1226);
   U97 : NAND2X1 port map( A => PLAINKEY_29_port, B => n232, Y => n80);
   U99 : OAI21X1 port map( A => n230, B => n1543, C => n82, Y => n1227);
   U100 : NAND2X1 port map( A => PLAINKEY_30_port, B => n232, Y => n82);
   U102 : OAI21X1 port map( A => n229, B => n1542, C => n84, Y => n1228);
   U103 : NAND2X1 port map( A => PLAINKEY_31_port, B => n232, Y => n84);
   U105 : OAI21X1 port map( A => RST, B => n1541, C => n86, Y => n1229);
   U106 : NAND2X1 port map( A => PLAINKEY_32_port, B => n232, Y => n86);
   U108 : OAI21X1 port map( A => n230, B => n1540, C => n88, Y => n1230);
   U109 : NAND2X1 port map( A => PLAINKEY_33_port, B => n232, Y => n88);
   U111 : OAI21X1 port map( A => n233, B => n1539, C => n90, Y => n1231);
   U112 : NAND2X1 port map( A => PLAINKEY_34_port, B => n232, Y => n90);
   U114 : OAI21X1 port map( A => n230, B => n1538, C => n92, Y => n1232);
   U115 : NAND2X1 port map( A => PLAINKEY_35_port, B => n232, Y => n92);
   U117 : OAI21X1 port map( A => n230, B => n1537, C => n94, Y => n1233);
   U118 : NAND2X1 port map( A => PLAINKEY_36_port, B => n232, Y => n94);
   U120 : OAI21X1 port map( A => n231, B => n1536, C => n96, Y => n1234);
   U121 : NAND2X1 port map( A => PLAINKEY_37_port, B => n232, Y => n96);
   U123 : OAI21X1 port map( A => n227, B => n1535, C => n98, Y => n1235);
   U124 : NAND2X1 port map( A => PLAINKEY_38_port, B => n232, Y => n98);
   U126 : OAI21X1 port map( A => n230, B => n1534, C => n100, Y => n1236);
   U127 : NAND2X1 port map( A => PLAINKEY_39_port, B => n232, Y => n100);
   U129 : OAI21X1 port map( A => n229, B => n1533, C => n102, Y => n1237);
   U130 : NAND2X1 port map( A => PLAINKEY_40_port, B => n232, Y => n102);
   U132 : OAI21X1 port map( A => n230, B => n1532, C => n104, Y => n1238);
   U133 : NAND2X1 port map( A => PLAINKEY_41_port, B => n232, Y => n104);
   U135 : OAI21X1 port map( A => n230, B => n1531, C => n106, Y => n1239);
   U136 : NAND2X1 port map( A => PLAINKEY_42_port, B => n232, Y => n106);
   U138 : OAI21X1 port map( A => RST, B => n1530, C => n108, Y => n1240);
   U139 : NAND2X1 port map( A => PLAINKEY_43_port, B => n232, Y => n108);
   U141 : OAI21X1 port map( A => n228, B => n1529, C => n110, Y => n1241);
   U142 : NAND2X1 port map( A => PLAINKEY_44_port, B => n231, Y => n110);
   U144 : OAI21X1 port map( A => n228, B => n1528, C => n112, Y => n1242);
   U145 : NAND2X1 port map( A => PLAINKEY_45_port, B => n231, Y => n112);
   U147 : OAI21X1 port map( A => n232, B => n1527, C => n114, Y => n1243);
   U148 : NAND2X1 port map( A => PLAINKEY_46_port, B => n232, Y => n114);
   U150 : OAI21X1 port map( A => n228, B => n1526, C => n116, Y => n1244);
   U151 : NAND2X1 port map( A => PLAINKEY_47_port, B => n231, Y => n116);
   U153 : OAI21X1 port map( A => n230, B => n1525, C => n118, Y => n1245);
   U154 : NAND2X1 port map( A => PLAINKEY_48_port, B => n231, Y => n118);
   U156 : OAI21X1 port map( A => n230, B => n1524, C => n120, Y => n1246);
   U157 : NAND2X1 port map( A => PLAINKEY_49_port, B => n231, Y => n120);
   U159 : OAI21X1 port map( A => n230, B => n1523, C => n122, Y => n1247);
   U160 : NAND2X1 port map( A => PLAINKEY_50_port, B => n231, Y => n122);
   U162 : OAI21X1 port map( A => n229, B => n1522, C => n124, Y => n1248);
   U163 : NAND2X1 port map( A => PLAINKEY_51_port, B => n231, Y => n124);
   U165 : OAI21X1 port map( A => n230, B => n1521, C => n126, Y => n1249);
   U166 : NAND2X1 port map( A => PLAINKEY_52_port, B => n231, Y => n126);
   U168 : OAI21X1 port map( A => n229, B => n1520, C => n128, Y => n1250);
   U169 : NAND2X1 port map( A => PLAINKEY_53_port, B => n231, Y => n128);
   U171 : OAI21X1 port map( A => n229, B => n1519, C => n130, Y => n1251);
   U172 : NAND2X1 port map( A => PLAINKEY_54_port, B => n231, Y => n130);
   U174 : OAI21X1 port map( A => n228, B => n1518, C => n132, Y => n1252);
   U175 : NAND2X1 port map( A => PLAINKEY_55_port, B => n232, Y => n132);
   U177 : OAI21X1 port map( A => n229, B => n1517, C => n134, Y => n1253);
   U178 : NAND2X1 port map( A => PLAINKEY_56_port, B => n231, Y => n134);
   U180 : OAI21X1 port map( A => n228, B => n1516, C => n136, Y => n1254);
   U181 : NAND2X1 port map( A => PLAINKEY_57_port, B => n231, Y => n136);
   U183 : OAI21X1 port map( A => n228, B => n1515, C => n138, Y => n1255);
   U184 : NAND2X1 port map( A => PLAINKEY_58_port, B => n231, Y => n138);
   U186 : OAI21X1 port map( A => n228, B => n1514, C => n140, Y => n1256);
   U187 : NAND2X1 port map( A => PLAINKEY_59_port, B => n231, Y => n140);
   U188 : OAI21X1 port map( A => n227, B => n1513, C => n142, Y => n1257);
   U189 : NAND2X1 port map( A => PLAINKEY_60_port, B => n231, Y => n142);
   U191 : OAI21X1 port map( A => n227, B => n1512, C => n144, Y => n1258);
   U192 : NAND2X1 port map( A => PLAINKEY_61_port, B => n231, Y => n144);
   U194 : OAI21X1 port map( A => n227, B => n1511, C => n146, Y => n1259);
   U195 : NAND2X1 port map( A => PLAINKEY_62_port, B => n231, Y => n146);
   U196 : OAI21X1 port map( A => n227, B => n1510, C => n148, Y => n1260);
   U197 : NAND2X1 port map( A => PLAINKEY_63_port, B => n232, Y => n148);
   U202 : OAI21X1 port map( A => n1449, B => n162, C => n157, Y => n155);
   U203 : AOI22X1 port map( A => n163, B => n164, C => n1498, D => n1576, Y => 
                           n162);
   U205 : OAI22X1 port map( A => RCV_DATA(3), B => n167, C => n1499, D => n169,
                           Y => n163);
   U206 : AOI22X1 port map( A => n170, B => n171, C => n1500, D => n1578, Y => 
                           n169);
   U208 : OAI22X1 port map( A => n174, B => n1501, C => RCV_DATA(1), D => n176,
                           Y => n170);
   U210 : NAND2X1 port map( A => n33, B => n14, Y => n176);
   U211 : AOI22X1 port map( A => n179, B => n156, C => n1507, D => n1510, Y => 
                           n174);
   U213 : NOR2X1 port map( A => n182, B => n149, Y => n179);
   U220 : OAI22X1 port map( A => n157, B => n1575, C => n159, D => n1576, Y => 
                           n191);
   U221 : OAI21X1 port map( A => n164, B => n1577, C => n194, Y => n190);
   U222 : AOI22X1 port map( A => RCV_DATA(2), B => n1499, C => n1496, D => n196
                           , Y => n194);
   U223 : OAI21X1 port map( A => n171, B => n226, C => n198, Y => n196);
   U224 : NAND2X1 port map( A => n199, B => n171, Y => n198);
   U225 : OAI21X1 port map( A => n182, B => n200, C => n201, Y => n199);
   U226 : OAI21X1 port map( A => n202, B => n182, C => currentPlainKey_62_port,
                           Y => n201);
   U227 : NAND2X1 port map( A => n31, B => n14, Y => n171);
   U233 : OAI21X1 port map( A => n212, B => n213, C => n152, Y => n211);
   U234 : OAI22X1 port map( A => n157, B => n1576, C => n164, D => n1578, Y => 
                           n213);
   U235 : OAI21X1 port map( A => n214, B => n204, C => n215, Y => n212);
   U236 : AOI22X1 port map( A => n225, B => n1499, C => RCV_DATA(3), D => n1449
                           , Y => n215);
   U238 : NAND2X1 port map( A => n216, B => n167, Y => n204);
   U239 : NAND2X1 port map( A => n29, B => n14, Y => n167);
   U240 : AOI22X1 port map( A => n218, B => n158, C => currentPlainKey_61_port,
                           D => n1506, Y => n214);
   U242 : NOR2X1 port map( A => n182, B => n220, Y => n218);
   U252 : OAI21X1 port map( A => n182, B => n236, C => n237, Y => n235);
   U253 : OAI21X1 port map( A => n238, B => n182, C => currentPlainKey_60_port,
                           Y => n237);
   U264 : OAI21X1 port map( A => n157, B => n1578, C => n252, Y => n251);
   U265 : AOI22X1 port map( A => n239, B => n253, C => n225, D => n1449, Y => 
                           n252);
   U266 : OAI22X1 port map( A => n254, B => n1514, C => n156, D => n1505, Y => 
                           n253);
   U270 : NOR2X1 port map( A => n182, B => n256, Y => n254);
   U271 : NOR2X1 port map( A => n1449, B => n1497, Y => n239);
   U284 : OAI22X1 port map( A => n157, B => n226, C => n1497, D => n273, Y => 
                           n272);
   U285 : AOI22X1 port map( A => n274, B => n158, C => currentPlainKey_58_port,
                           D => n1504, Y => n273);
   U287 : NOR2X1 port map( A => n182, B => n276, Y => n274);
   U300 : AOI22X1 port map( A => n290, B => n152, C => n225, D => n1450, Y => 
                           n288);
   U303 : OAI21X1 port map( A => n182, B => n292, C => n293, Y => n290);
   U304 : OAI21X1 port map( A => n294, B => n182, C => currentPlainKey_57_port,
                           Y => n293);
   U314 : OAI21X1 port map( A => n182, B => n307, C => n308, Y => n306);
   U315 : OAI21X1 port map( A => n309, B => n182, C => currentPlainKey_56_port,
                           Y => n308);
   U316 : NAND2X1 port map( A => address_3_port, B => n310, Y => n182);
   U330 : AOI22X1 port map( A => n325, B => n246, C => n1451, D => n225, Y => 
                           n323);
   U333 : OAI21X1 port map( A => n173, B => n328, C => n329, Y => n325);
   U334 : OAI21X1 port map( A => n149, B => n173, C => currentPlainKey_55_port,
                           Y => n329);
   U344 : OAI21X1 port map( A => n200, B => n173, C => n342, Y => n341);
   U345 : OAI21X1 port map( A => n202, B => n173, C => currentPlainKey_54_port,
                           Y => n342);
   U359 : AOI22X1 port map( A => n356, B => n283, C => n1452, D => RCV_DATA(1),
                           Y => n354);
   U362 : OAI21X1 port map( A => n173, B => n358, C => n359, Y => n356);
   U363 : OAI21X1 port map( A => n220, B => n173, C => currentPlainKey_53_port,
                           Y => n359);
   U373 : OAI21X1 port map( A => n236, B => n173, C => n372, Y => n371);
   U374 : OAI21X1 port map( A => n238, B => n173, C => currentPlainKey_52_port,
                           Y => n372);
   U388 : AOI22X1 port map( A => n386, B => n318, C => n1453, D => n225, Y => 
                           n384);
   U391 : OAI21X1 port map( A => n173, B => n388, C => n389, Y => n386);
   U392 : OAI21X1 port map( A => n256, B => n173, C => currentPlainKey_51_port,
                           Y => n389);
   U402 : OAI21X1 port map( A => n173, B => n402, C => n403, Y => n401);
   U403 : OAI21X1 port map( A => n276, B => n173, C => currentPlainKey_50_port,
                           Y => n403);
   U417 : AOI22X1 port map( A => n417, B => n349, C => n1454, D => RCV_DATA(1),
                           Y => n415);
   U422 : OAI21X1 port map( A => n292, B => n173, C => n421, Y => n417);
   U423 : OAI21X1 port map( A => n294, B => n173, C => currentPlainKey_49_port,
                           Y => n421);
   U433 : OAI21X1 port map( A => n307, B => n173, C => n434, Y => n433);
   U434 : OAI21X1 port map( A => n309, B => n173, C => currentPlainKey_48_port,
                           Y => n434);
   U449 : AOI22X1 port map( A => n449, B => n379, C => n1455, D => n225, Y => 
                           n447);
   U452 : OAI21X1 port map( A => n328, B => n172, C => n451, Y => n449);
   U453 : OAI21X1 port map( A => n149, B => n172, C => currentPlainKey_47_port,
                           Y => n451);
   U463 : OAI21X1 port map( A => n200, B => n172, C => n464, Y => n463);
   U464 : OAI21X1 port map( A => n202, B => n172, C => currentPlainKey_46_port,
                           Y => n464);
   U478 : AOI22X1 port map( A => n477, B => n410, C => n1456, D => RCV_DATA(1),
                           Y => n475);
   U481 : OAI21X1 port map( A => n358, B => n172, C => n478, Y => n477);
   U482 : OAI21X1 port map( A => n220, B => n172, C => currentPlainKey_45_port,
                           Y => n478);
   U492 : OAI21X1 port map( A => n236, B => n172, C => n491, Y => n490);
   U493 : OAI21X1 port map( A => n238, B => n172, C => currentPlainKey_44_port,
                           Y => n491);
   U507 : AOI22X1 port map( A => n504, B => n442, C => n1457, D => n225, Y => 
                           n502);
   U510 : OAI21X1 port map( A => n388, B => n172, C => n505, Y => n504);
   U511 : OAI21X1 port map( A => n256, B => n172, C => currentPlainKey_43_port,
                           Y => n505);
   U521 : OAI21X1 port map( A => n402, B => n172, C => n518, Y => n517);
   U522 : OAI21X1 port map( A => n276, B => n172, C => currentPlainKey_42_port,
                           Y => n518);
   U536 : AOI22X1 port map( A => n531, B => n470, C => n1458, D => n225, Y => 
                           n529);
   U539 : OAI21X1 port map( A => n292, B => n172, C => n532, Y => n531);
   U540 : OAI21X1 port map( A => n294, B => n172, C => currentPlainKey_41_port,
                           Y => n532);
   U550 : OAI21X1 port map( A => n307, B => n172, C => n545, Y => n544);
   U551 : OAI21X1 port map( A => n309, B => n172, C => currentPlainKey_40_port,
                           Y => n545);
   U566 : AOI22X1 port map( A => n560, B => n497, C => n1459, D => n225, Y => 
                           n558);
   U569 : OAI21X1 port map( A => n328, B => n168, C => n562, Y => n560);
   U570 : OAI21X1 port map( A => n149, B => n168, C => currentPlainKey_39_port,
                           Y => n562);
   U580 : OAI21X1 port map( A => n200, B => n168, C => n575, Y => n574);
   U581 : OAI21X1 port map( A => n202, B => n168, C => currentPlainKey_38_port,
                           Y => n575);
   U595 : AOI22X1 port map( A => n588, B => n524, C => n1460, D => RCV_DATA(1),
                           Y => n586);
   U598 : OAI21X1 port map( A => n358, B => n168, C => n589, Y => n588);
   U599 : OAI21X1 port map( A => n220, B => n168, C => currentPlainKey_37_port,
                           Y => n589);
   U609 : OAI21X1 port map( A => n236, B => n168, C => n602, Y => n601);
   U610 : OAI21X1 port map( A => n238, B => n168, C => currentPlainKey_36_port,
                           Y => n602);
   U624 : AOI22X1 port map( A => n615, B => n553, C => n1461, D => n225, Y => 
                           n613);
   U627 : OAI21X1 port map( A => n388, B => n168, C => n616, Y => n615);
   U628 : OAI21X1 port map( A => n256, B => n168, C => currentPlainKey_35_port,
                           Y => n616);
   U638 : OAI21X1 port map( A => n402, B => n168, C => n629, Y => n628);
   U639 : OAI21X1 port map( A => n276, B => n168, C => currentPlainKey_34_port,
                           Y => n629);
   U653 : AOI22X1 port map( A => n642, B => n581, C => n1462, D => n225, Y => 
                           n640);
   U658 : OAI21X1 port map( A => n292, B => n168, C => n643, Y => n642);
   U659 : OAI21X1 port map( A => n294, B => n168, C => currentPlainKey_33_port,
                           Y => n643);
   U669 : OAI21X1 port map( A => n307, B => n168, C => n656, Y => n655);
   U670 : OAI21X1 port map( A => n309, B => n168, C => currentPlainKey_32_port,
                           Y => n656);
   U672 : NOR2X1 port map( A => n1508, B => address_4_port, Y => n546);
   U686 : AOI22X1 port map( A => n671, B => n608, C => n1463, D => n225, Y => 
                           n669);
   U689 : OAI21X1 port map( A => n328, B => n166, C => n673, Y => n671);
   U690 : OAI21X1 port map( A => n149, B => n166, C => currentPlainKey_31_port,
                           Y => n673);
   U700 : OAI21X1 port map( A => n200, B => n166, C => n686, Y => n685);
   U701 : OAI21X1 port map( A => n202, B => n166, C => currentPlainKey_30_port,
                           Y => n686);
   U715 : AOI22X1 port map( A => n699, B => n635, C => n1464, D => n225, Y => 
                           n697);
   U718 : OAI21X1 port map( A => n358, B => n166, C => n700, Y => n699);
   U719 : OAI21X1 port map( A => n220, B => n166, C => currentPlainKey_29_port,
                           Y => n700);
   U729 : OAI21X1 port map( A => n236, B => n166, C => n713, Y => n712);
   U730 : OAI21X1 port map( A => n238, B => n166, C => currentPlainKey_28_port,
                           Y => n713);
   U744 : AOI22X1 port map( A => n726, B => n664, C => n1465, D => n225, Y => 
                           n724);
   U747 : OAI21X1 port map( A => n388, B => n166, C => n727, Y => n726);
   U748 : OAI21X1 port map( A => n256, B => n166, C => currentPlainKey_27_port,
                           Y => n727);
   U758 : OAI21X1 port map( A => n402, B => n166, C => n740, Y => n739);
   U759 : OAI21X1 port map( A => n276, B => n166, C => currentPlainKey_26_port,
                           Y => n740);
   U773 : AOI22X1 port map( A => n753, B => n692, C => n1466, D => n225, Y => 
                           n751);
   U776 : OAI21X1 port map( A => n292, B => n166, C => n754, Y => n753);
   U777 : OAI21X1 port map( A => n294, B => n166, C => currentPlainKey_25_port,
                           Y => n754);
   U787 : OAI21X1 port map( A => n307, B => n166, C => n767, Y => n766);
   U788 : OAI21X1 port map( A => n309, B => n166, C => currentPlainKey_24_port,
                           Y => n767);
   U803 : AOI22X1 port map( A => n782, B => n719, C => n1467, D => n225, Y => 
                           n780);
   U806 : OAI21X1 port map( A => n328, B => n165, C => n784, Y => n782);
   U807 : OAI21X1 port map( A => n149, B => n165, C => currentPlainKey_23_port,
                           Y => n784);
   U817 : OAI21X1 port map( A => n200, B => n165, C => n797, Y => n796);
   U818 : OAI21X1 port map( A => n202, B => n165, C => currentPlainKey_22_port,
                           Y => n797);
   U832 : AOI22X1 port map( A => n810, B => n746, C => n1468, D => n225, Y => 
                           n808);
   U835 : OAI21X1 port map( A => n358, B => n165, C => n811, Y => n810);
   U836 : OAI21X1 port map( A => n220, B => n165, C => currentPlainKey_21_port,
                           Y => n811);
   U846 : OAI21X1 port map( A => n236, B => n165, C => n824, Y => n823);
   U847 : OAI21X1 port map( A => n238, B => n165, C => currentPlainKey_20_port,
                           Y => n824);
   U861 : AOI22X1 port map( A => n837, B => n775, C => n1469, D => n225, Y => 
                           n835);
   U864 : OAI21X1 port map( A => n388, B => n165, C => n838, Y => n837);
   U865 : OAI21X1 port map( A => n256, B => n165, C => currentPlainKey_19_port,
                           Y => n838);
   U875 : OAI21X1 port map( A => n402, B => n165, C => n851, Y => n850);
   U876 : OAI21X1 port map( A => n276, B => n165, C => currentPlainKey_18_port,
                           Y => n851);
   U890 : AOI22X1 port map( A => n864, B => n803, C => n1470, D => n225, Y => 
                           n862);
   U895 : OAI21X1 port map( A => n292, B => n165, C => n865, Y => n864);
   U896 : OAI21X1 port map( A => n294, B => n165, C => currentPlainKey_17_port,
                           Y => n865);
   U906 : OAI21X1 port map( A => n307, B => n165, C => n878, Y => n877);
   U907 : OAI21X1 port map( A => n309, B => n165, C => currentPlainKey_16_port,
                           Y => n878);
   U909 : NOR2X1 port map( A => n1509, B => address_5_port, Y => n768);
   U923 : AOI22X1 port map( A => n893, B => n830, C => n1471, D => n225, Y => 
                           n891);
   U926 : OAI21X1 port map( A => n328, B => n161, C => n895, Y => n893);
   U927 : OAI21X1 port map( A => n149, B => n161, C => currentPlainKey_15_port,
                           Y => n895);
   U937 : OAI21X1 port map( A => n200, B => n161, C => n908, Y => n907);
   U938 : OAI21X1 port map( A => n202, B => n161, C => currentPlainKey_14_port,
                           Y => n908);
   U952 : AOI22X1 port map( A => n921, B => n857, C => n1472, D => n225, Y => 
                           n919);
   U955 : OAI21X1 port map( A => n358, B => n161, C => n922, Y => n921);
   U956 : OAI21X1 port map( A => n220, B => n161, C => currentPlainKey_13_port,
                           Y => n922);
   U966 : OAI21X1 port map( A => n236, B => n161, C => n935, Y => n934);
   U967 : OAI21X1 port map( A => n238, B => n161, C => currentPlainKey_12_port,
                           Y => n935);
   U981 : AOI22X1 port map( A => n948, B => n886, C => n1473, D => n225, Y => 
                           n946);
   U984 : OAI21X1 port map( A => n388, B => n161, C => n949, Y => n948);
   U985 : OAI21X1 port map( A => n256, B => n161, C => currentPlainKey_11_port,
                           Y => n949);
   U995 : OAI21X1 port map( A => n402, B => n161, C => n962, Y => n961);
   U996 : OAI21X1 port map( A => n276, B => n161, C => currentPlainKey_10_port,
                           Y => n962);
   U1010 : AOI22X1 port map( A => n975, B => n914, C => n1474, D => n225, Y => 
                           n973);
   U1014 : OAI21X1 port map( A => n292, B => n161, C => n976, Y => n975);
   U1015 : OAI21X1 port map( A => n294, B => n161, C => currentPlainKey_9_port,
                           Y => n976);
   U1025 : OAI21X1 port map( A => n307, B => n161, C => n989, Y => n988);
   U1026 : OAI21X1 port map( A => n309, B => n161, C => currentPlainKey_8_port,
                           Y => n989);
   U1041 : AOI22X1 port map( A => n1004, B => n941, C => n1475, D => n225, Y =>
                           n1002);
   U1044 : OAI21X1 port map( A => n328, B => n160, C => n1006, Y => n1004);
   U1045 : OAI21X1 port map( A => n149, B => n160, C => currentPlainKey_7_port,
                           Y => n1006);
   U1046 : NAND2X1 port map( A => n158, B => n16, Y => n328);
   U1057 : OAI21X1 port map( A => n200, B => n160, C => n1019, Y => n1018);
   U1058 : OAI21X1 port map( A => n202, B => n160, C => currentPlainKey_6_port,
                           Y => n1019);
   U1059 : NAND2X1 port map( A => n158, B => n147, Y => n200);
   U1074 : AOI22X1 port map( A => n1033, B => n968, C => n1476, D => n225, Y =>
                           n1031);
   U1077 : OAI21X1 port map( A => n358, B => n160, C => n1034, Y => n1033);
   U1078 : OAI21X1 port map( A => n220, B => n160, C => currentPlainKey_5_port,
                           Y => n1034);
   U1079 : NAND2X1 port map( A => n158, B => n1478, Y => n358);
   U1090 : OAI21X1 port map( A => n236, B => n160, C => n1047, Y => n1046);
   U1091 : OAI21X1 port map( A => n238, B => n160, C => currentPlainKey_4_port,
                           Y => n1047);
   U1092 : NAND2X1 port map( A => n158, B => n150, Y => n236);
   U1111 : OAI21X1 port map( A => n388, B => n160, C => n1063, Y => n1062);
   U1112 : OAI21X1 port map( A => n256, B => n160, C => currentPlainKey_3_port,
                           Y => n1063);
   U1113 : NAND2X1 port map( A => n158, B => n1481, Y => n388);
   U1126 : OAI21X1 port map( A => n402, B => n160, C => n1078, Y => n1077);
   U1127 : OAI21X1 port map( A => n276, B => n160, C => currentPlainKey_2_port,
                           Y => n1078);
   U1128 : NAND2X1 port map( A => n158, B => n151, Y => n402);
   U1154 : NOR2X1 port map( A => address_6_port, B => address_7_port, Y => n420
                           );
   U1155 : OAI21X1 port map( A => n292, B => n160, C => n1090, Y => n1089);
   U1156 : OAI21X1 port map( A => n294, B => n160, C => currentPlainKey_1_port,
                           Y => n1090);
   U1157 : NAND2X1 port map( A => n158, B => n143, Y => n292);
   U1182 : AOI22X1 port map( A => n21, B => n1576, C => n1103, D => n1104, Y =>
                           n1101);
   U1183 : AOI21X1 port map( A => n1105, B => n1038, C => n21, Y => n1104);
   U1184 : OAI21X1 port map( A => n226, B => n1011, C => n1106, Y => n1105);
   U1185 : NAND2X1 port map( A => n25, B => n1107, Y => n1106);
   U1186 : OAI21X1 port map( A => n307, B => n160, C => n1108, Y => n1107);
   U1187 : OAI21X1 port map( A => n309, B => n160, C => currentPlainKey_0_port,
                           Y => n1108);
   U1189 : NOR2X1 port map( A => address_4_port, B => address_5_port, Y => n990
                           );
   U1190 : NAND2X1 port map( A => n158, B => n1477, Y => n307);
   U1199 : AOI22X1 port map( A => n1479, B => RCV_DATA(2), C => n1502, D => 
                           RCV_DATA(3), Y => n1103);
   U1220 : NOR2X1 port map( A => n1508, B => n1509, Y => n310);
   U1273 : OAI21X1 port map( A => n1480, B => n1484, C => n1143, Y => n1349);
   U1274 : NAND3X1 port map( A => keyCount_0_port, B => n1484, C => n1144, Y =>
                           n1143);
   U1305 : NAND2X1 port map( A => n1579, B => n1574, Y => n1178);
   U1314 : NAND3X1 port map( A => keyCount_2_port, B => keyCount_1_port, C => 
                           n1186, Y => n1160);
   U1315 : NOR2X1 port map( A => keyCount_3_port, B => n1483, Y => n1186);
   U254 : AND2X2 port map( A => n239, B => n164, Y => n216);
   r577 : keyreg_1_DW01_add_0 port map( A(7) => parityAccumulator_7_port, A(6) 
                           => parityAccumulator_6_port, A(5) => 
                           parityAccumulator_5_port, A(4) => 
                           parityAccumulator_4_port, A(3) => 
                           parityAccumulator_3_port, A(2) => 
                           parityAccumulator_2_port, A(1) => 
                           parityAccumulator_1_port, A(0) => 
                           parityAccumulator_0_port, B(7) => RCV_DATA(7), B(6) 
                           => RCV_DATA(6), B(5) => RCV_DATA(5), B(4) => 
                           RCV_DATA(4), B(3) => RCV_DATA(3), B(2) => 
                           RCV_DATA(2), B(1) => RCV_DATA(1), B(0) => n158, CI 
                           => n3, SUM(7) => N1799, SUM(6) => N1798, SUM(5) => 
                           N1797, SUM(4) => N1796, SUM(3) => N1795, SUM(2) => 
                           N1794, SUM(1) => N1793, SUM(0) => N1792, CO => 
                           n_1025);
   state_reg_3_inst : DFFSR port map( D => n1354, CLK => CLK, R => n243, S => 
                           n81, Q => state_3_port);
   state_reg_2_inst : DFFSR port map( D => n1352, CLK => CLK, R => n243, S => 
                           n79, Q => state_2_port);
   state_reg_0_inst : DFFSR port map( D => n1353, CLK => CLK, R => n243, S => 
                           n77, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => n1351, CLK => CLK, R => n243, S => 
                           n75, Q => state_1_port);
   parityError_reg : DFFSR port map( D => nextParityError, CLK => CLK, R => 
                           n243, S => n73, Q => parityError);
   PARITY_ERROR_reg : DFFSR port map( D => nextParityError, CLK => CLK, R => 
                           n243, S => n71, Q => PARITY_ERROR);
   U3 : INVX4 port map( A => n327, Y => n1363);
   U4 : BUFX4 port map( A => n1363, Y => n210);
   U5 : BUFX4 port map( A => n1363, Y => n209);
   U7 : BUFX4 port map( A => n1363, Y => n217);
   U8 : INVX1 port map( A => n1367, Y => n1);
   U23 : INVX1 port map( A => n1367, Y => n2);
   U26 : INVX1 port map( A => n1367, Y => n4);
   U29 : INVX8 port map( A => n1174, Y => n1367);
   U32 : INVX2 port map( A => n1172, Y => n1184);
   U35 : BUFX2 port map( A => n1184, Y => n195);
   U38 : BUFX2 port map( A => n1417, Y => n89);
   U41 : BUFX2 port map( A => n1370, Y => n224);
   U44 : BUFX2 port map( A => n1370, Y => n219);
   U47 : INVX2 port map( A => n1409, Y => n5);
   U50 : INVX2 port map( A => n5, Y => n6);
   U53 : INVX1 port map( A => n5, Y => n7);
   U56 : AND2X2 port map( A => n105, B => n1482, Y => n8);
   U59 : AND2X2 port map( A => n107, B => n1482, Y => n9);
   U62 : AND2X2 port map( A => n109, B => n1482, Y => n10);
   U65 : AND2X2 port map( A => n14, B => n1482, Y => n11);
   U68 : INVX2 port map( A => n139, Y => n141);
   U71 : AND2X2 port map( A => n310, B => n420, Y => n14);
   U74 : AND2X2 port map( A => n65, B => address_0_port, Y => n16);
   U77 : INVX2 port map( A => n95, Y => n178);
   U80 : INVX2 port map( A => n178, Y => n177);
   U83 : NAND2X1 port map( A => n177, B => RCV_DATA(3), Y => n17);
   U86 : AND2X2 port map( A => n131, B => n141, Y => n19);
   U89 : AND2X2 port map( A => n1481, B => address_3_port, Y => n20);
   U92 : AND2X2 port map( A => n271, B => n29, Y => n21);
   U95 : AND2X2 port map( A => n271, B => n20, Y => n23);
   U98 : INVX2 port map( A => n189, Y => n185);
   U101 : INVX2 port map( A => n189, Y => n186);
   U104 : INVX2 port map( A => n131, Y => n133);
   U107 : AND2X2 port map( A => n300, B => n1011, Y => n25);
   U110 : AND2X2 port map( A => n151, B => address_3_port, Y => n27);
   U113 : AND2X2 port map( A => n150, B => address_3_port, Y => n29);
   U116 : AND2X2 port map( A => n1478, B => address_3_port, Y => n31);
   U119 : AND2X2 port map( A => n147, B => address_3_port, Y => n33);
   U122 : AND2X2 port map( A => n16, B => address_3_port, Y => n35);
   U125 : AND2X2 port map( A => n1477, B => address_3_port, Y => n37);
   U128 : AND2X2 port map( A => n319, B => n347, Y => n39);
   U131 : AND2X2 port map( A => n410, B => n1016, Y => n41);
   U134 : AND2X2 port map( A => n470, B => n955, Y => n43);
   U137 : AND2X2 port map( A => n914, B => n460, Y => n45);
   U140 : AND2X2 port map( A => n857, B => n522, Y => n47);
   U143 : AND2X2 port map( A => n692, B => n707, Y => n49);
   U146 : AND2X2 port map( A => n635, B => n770, Y => n51);
   U149 : AND2X2 port map( A => n968, B => n397, Y => n53);
   U152 : AND2X2 port map( A => n803, B => n584, Y => n55);
   U155 : AND2X2 port map( A => n746, B => n647, Y => n57);
   U158 : AND2X2 port map( A => n581, B => n831, Y => n59);
   U161 : AND2X2 port map( A => n524, B => n892, Y => n61);
   U164 : AND2X2 port map( A => n349, B => n1074, Y => n63);
   U167 : AND2X2 port map( A => address_1_port, B => address_2_port, Y => n65);
   U170 : AND2X2 port map( A => n216, B => n235, Y => n67);
   U173 : AND2X2 port map( A => n271, B => n27, Y => n69);
   n71 <= '1';
   n73 <= '1';
   n75 <= '1';
   n77 <= '1';
   n79 <= '1';
   n81 <= '1';
   U198 : INVX1 port map( A => n332, Y => n333);
   U199 : AND2X2 port map( A => n85, B => RCV_DATA(1), Y => n99);
   U200 : AND2X1 port map( A => n117, B => n19, Y => n83);
   U201 : INVX1 port map( A => n83, Y => n1432);
   U204 : BUFX2 port map( A => n177, Y => n85);
   U207 : BUFX4 port map( A => n177, Y => n87);
   U209 : AND2X2 port map( A => n91, B => n1263, Y => n1164);
   U212 : NOR2X1 port map( A => n1162, B => n1450, Y => n91);
   U214 : INVX2 port map( A => n226, Y => n225);
   U215 : BUFX2 port map( A => n17, Y => n97);
   U216 : INVX2 port map( A => n184, Y => n180);
   U217 : INVX2 port map( A => n1387, Y => n93);
   U218 : AND2X2 port map( A => n101, B => n1425, Y => n95);
   U219 : INVX1 port map( A => n95, Y => n1364);
   U228 : INVX2 port map( A => n178, Y => n175);
   U229 : INVX4 port map( A => n153, Y => n1136);
   U230 : INVX2 port map( A => n156, Y => n158);
   U231 : AND2X1 port map( A => n177, B => RCV_DATA(2), Y => n119);
   U232 : INVX2 port map( A => n240, Y => n230);
   U237 : INVX2 port map( A => n240, Y => n229);
   U241 : INVX2 port map( A => n234, Y => n228);
   U243 : INVX2 port map( A => n234, Y => n227);
   U244 : INVX2 port map( A => n241, Y => n231);
   U245 : INVX2 port map( A => n241, Y => n232);
   U246 : INVX2 port map( A => n242, Y => n233);
   U247 : INVX2 port map( A => n208, Y => n207);
   U248 : BUFX2 port map( A => n243, Y => n241);
   U249 : BUFX2 port map( A => n241, Y => n240);
   U250 : BUFX2 port map( A => n242, Y => n234);
   U251 : BUFX2 port map( A => n243, Y => n242);
   U255 : INVX2 port map( A => n99, Y => n154);
   U256 : INVX2 port map( A => n99, Y => n153);
   U257 : INVX2 port map( A => n208, Y => n206);
   U258 : INVX2 port map( A => n208, Y => n205);
   U259 : INVX2 port map( A => RST, Y => n243);
   U260 : BUFX2 port map( A => n1370, Y => n221);
   U261 : BUFX2 port map( A => n1370, Y => n222);
   U262 : BUFX2 port map( A => n1370, Y => n223);
   U263 : INVX2 port map( A => n184, Y => n181);
   U267 : BUFX2 port map( A => n1184, Y => n197);
   U268 : BUFX2 port map( A => n1184, Y => n193);
   U269 : BUFX2 port map( A => n1184, Y => n192);
   U272 : AND2X2 port map( A => n269, B => n1419, Y => n101);
   U273 : INVX2 port map( A => n184, Y => n183);
   U274 : INVX2 port map( A => n188, Y => n187);
   U275 : BUFX2 port map( A => n1184, Y => n203);
   U276 : INVX2 port map( A => n103, Y => n160);
   U277 : INVX2 port map( A => n111, Y => n173);
   U278 : INVX2 port map( A => n113, Y => n165);
   U279 : INVX2 port map( A => n115, Y => n168);
   U280 : INVX2 port map( A => n17, Y => n184);
   U281 : BUFX2 port map( A => n119, Y => n188);
   U282 : AND2X2 port map( A => n990, B => n1482, Y => n103);
   U283 : AND2X2 port map( A => n546, B => n420, Y => n105);
   U286 : AND2X2 port map( A => n990, B => n420, Y => n107);
   U288 : AND2X2 port map( A => n768, B => n420, Y => n109);
   U289 : INVX2 port map( A => n202, Y => n147);
   U290 : AND2X2 port map( A => n310, B => n1482, Y => n111);
   U291 : AND2X2 port map( A => n768, B => n1482, Y => n113);
   U292 : AND2X2 port map( A => n546, B => n1482, Y => n115);
   U293 : INVX2 port map( A => n121, Y => n161);
   U294 : INVX2 port map( A => n123, Y => n166);
   U295 : INVX2 port map( A => n125, Y => n172);
   U296 : INVX2 port map( A => RCV_DATA(1), Y => n226);
   U297 : AND2X2 port map( A => state_1_port, B => n1417, Y => n117);
   U298 : INVX2 port map( A => RCV_DATA(0), Y => n156);
   U299 : INVX2 port map( A => n294, Y => n143);
   U301 : INVX2 port map( A => n238, Y => n150);
   U302 : INVX2 port map( A => n276, Y => n151);
   U305 : INVX2 port map( A => n16, Y => n149);
   U306 : AND2X2 port map( A => n990, B => address_3_port, Y => n121);
   U307 : AND2X2 port map( A => n768, B => address_3_port, Y => n123);
   U308 : AND2X2 port map( A => n546, B => address_3_port, Y => n125);
   U309 : BUFX2 port map( A => n101, Y => n208);
   U310 : AND2X2 port map( A => n259, B => n129, Y => n127);
   U311 : BUFX2 port map( A => n1430, Y => n129);
   U312 : AND2X1 port map( A => n129, B => n93, Y => n1423);
   U313 : INVX2 port map( A => state_2_port, Y => n131);
   U317 : NOR2X1 port map( A => state_1_port, B => n141, Y => n135);
   U318 : INVX1 port map( A => n135, Y => n1413);
   U319 : INVX1 port map( A => state_1_port, Y => n250);
   U320 : INVX2 port map( A => n188, Y => n137);
   U321 : INVX2 port map( A => state_0_port, Y => n139);
   U322 : INVX1 port map( A => n7, Y => n1397);
   U323 : INVX1 port map( A => n7, Y => n1406);
   U324 : INVX1 port map( A => n7, Y => n1395);
   U325 : INVX1 port map( A => n7, Y => n1403);
   U326 : INVX1 port map( A => n7, Y => n1401);
   U327 : INVX1 port map( A => n7, Y => n1399);
   U328 : INVX1 port map( A => n7, Y => n1408);
   U329 : BUFX2 port map( A => n119, Y => n189);
   U331 : INVX1 port map( A => n1429, Y => n249);
   U332 : INVX1 port map( A => n1431, Y => n1387);
   U335 : INVX2 port map( A => n6, Y => n145);
   U336 : NAND2X1 port map( A => address_0_port, B => address_1_port, Y => n244
                           );
   U337 : OR2X2 port map( A => address_2_port, B => n244, Y => n256);
   U338 : INVX2 port map( A => n256, Y => n1481);
   U339 : NAND2X1 port map( A => n20, B => n14, Y => n164);
   U340 : INVX2 port map( A => address_2_port, Y => n267);
   U341 : INVX2 port map( A => address_1_port, Y => n266);
   U342 : NAND3X1 port map( A => address_0_port, B => n267, C => n266, Y => 
                           n294);
   U343 : NAND2X1 port map( A => n143, B => address_3_port, Y => n278);
   U346 : INVX2 port map( A => n278, Y => n925);
   U347 : NAND2X1 port map( A => n925, B => n14, Y => n157);
   U348 : INVX2 port map( A => state_3_port, Y => n1417);
   U349 : NAND3X1 port map( A => n117, B => n139, C => n131, Y => n1442);
   U350 : NAND3X1 port map( A => n133, B => n141, C => n117, Y => n1416);
   U351 : NAND2X1 port map( A => n1442, B => n1416, Y => CLR_RBUFF_port);
   U352 : NAND3X1 port map( A => n135, B => n133, C => n89, Y => n245);
   U353 : INVX2 port map( A => n245, Y => PROG_ERROR_port);
   U354 : NAND2X1 port map( A => n135, B => n131, Y => n1429);
   U355 : OAI21X1 port map( A => state_3_port, B => n1429, C => n1432, Y => 
                           n248);
   U356 : NAND3X1 port map( A => n117, B => n133, C => n139, Y => n1430);
   U357 : NAND2X1 port map( A => n1430, B => n245, Y => n247);
   U358 : NOR3X1 port map( A => CLR_RBUFF_port, B => n248, C => n247, Y => 
                           n1374);
   U360 : NAND2X1 port map( A => state_3_port, B => n249, Y => n1431);
   U361 : NAND3X1 port map( A => n141, B => n250, C => n1417, Y => n255);
   U364 : INVX2 port map( A => n255, Y => n257);
   U365 : NAND2X1 port map( A => n257, B => n133, Y => n1419);
   U366 : INVX2 port map( A => n1419, Y => n1439);
   U367 : NAND2X1 port map( A => n257, B => n131, Y => n259);
   U368 : INVX2 port map( A => n259, Y => n1386);
   U369 : AOI21X1 port map( A => n1439, B => parityError, C => n1386, Y => n258
                           );
   U370 : NAND3X1 port map( A => n1374, B => n1431, C => n258, Y => KEY_ERROR);
   U371 : NOR2X1 port map( A => PROG_ERROR_port, B => n227, Y => n261);
   U372 : NAND2X1 port map( A => n259, B => n1430, Y => n1424);
   U375 : NOR2X1 port map( A => n83, B => n1424, Y => n260);
   U376 : NAND3X1 port map( A => n261, B => n1431, C => n260, Y => n1409);
   U377 : NAND2X1 port map( A => n145, B => n1416, Y => n1446);
   U378 : INVX2 port map( A => n1446, Y => n269);
   U379 : INVX2 port map( A => n1442, Y => n1425);
   U380 : NAND2X1 port map( A => n269, B => n1425, Y => n1448);
   U381 : NOR2X1 port map( A => n1494, B => n1448, Y => n1144);
   U382 : NAND2X1 port map( A => keyCount_1_port, B => keyCount_0_port, Y => 
                           n262);
   U383 : NAND2X1 port map( A => n1425, B => n262, Y => n263);
   U384 : NAND2X1 port map( A => n269, B => n263, Y => n1443);
   U385 : INVX2 port map( A => n1443, Y => n1480);
   U386 : INVX2 port map( A => address_0_port, Y => n268);
   U387 : NAND2X1 port map( A => n65, B => n268, Y => n202);
   U389 : NAND3X1 port map( A => address_6_port, B => address_7_port, C => n310
                           , Y => n277);
   U390 : INVX2 port map( A => n277, Y => n271);
   U393 : NAND2X1 port map( A => n271, B => n33, Y => n300);
   U394 : INVX2 port map( A => n300, Y => n1479);
   U395 : NAND2X1 port map( A => address_0_port, B => address_2_port, Y => n264
                           );
   U396 : OR2X2 port map( A => address_1_port, B => n264, Y => n220);
   U397 : INVX2 port map( A => n220, Y => n1478);
   U398 : NAND2X1 port map( A => n271, B => n31, Y => n1038);
   U399 : INVX2 port map( A => n1038, Y => n1502);
   U400 : NOR2X1 port map( A => address_2_port, B => address_0_port, Y => n265)
                           ;
   U401 : NAND2X1 port map( A => n265, B => n266, Y => n309);
   U404 : INVX2 port map( A => n309, Y => n1477);
   U405 : INVX2 port map( A => address_3_port, Y => n1482);
   U406 : NAND2X1 port map( A => n271, B => n35, Y => n1011);
   U407 : NAND3X1 port map( A => address_2_port, B => n268, C => n266, Y => 
                           n238);
   U408 : INVX2 port map( A => RCV_DATA(4), Y => n1576);
   U409 : NAND3X1 port map( A => address_1_port, B => n268, C => n267, Y => 
                           n276);
   U410 : NAND2X1 port map( A => n9, B => n150, Y => n968);
   U411 : INVX2 port map( A => n968, Y => n1476);
   U412 : NAND2X1 port map( A => n9, B => n147, Y => n941);
   U413 : INVX2 port map( A => n941, Y => n1475);
   U414 : NAND2X1 port map( A => n107, B => n37, Y => n914);
   U415 : INVX2 port map( A => n914, Y => n1474);
   U416 : NAND2X1 port map( A => n107, B => n27, Y => n886);
   U418 : INVX2 port map( A => n886, Y => n1473);
   U419 : NAND2X1 port map( A => n107, B => n29, Y => n857);
   U420 : INVX2 port map( A => n857, Y => n1472);
   U421 : NAND2X1 port map( A => n107, B => n33, Y => n830);
   U424 : INVX2 port map( A => n830, Y => n1471);
   U425 : NAND2X1 port map( A => n10, B => n1477, Y => n803);
   U426 : INVX2 port map( A => n803, Y => n1470);
   U427 : NAND2X1 port map( A => n10, B => n151, Y => n775);
   U428 : INVX2 port map( A => n775, Y => n1469);
   U429 : NAND2X1 port map( A => n10, B => n150, Y => n746);
   U430 : INVX2 port map( A => n746, Y => n1468);
   U431 : NAND2X1 port map( A => n10, B => n147, Y => n719);
   U432 : INVX2 port map( A => n719, Y => n1467);
   U435 : NAND2X1 port map( A => n109, B => n37, Y => n692);
   U436 : INVX2 port map( A => n692, Y => n1466);
   U437 : NAND2X1 port map( A => n109, B => n27, Y => n664);
   U438 : INVX2 port map( A => n664, Y => n1465);
   U439 : NAND2X1 port map( A => n109, B => n29, Y => n635);
   U440 : INVX2 port map( A => n635, Y => n1464);
   U441 : NAND2X1 port map( A => n109, B => n33, Y => n608);
   U442 : INVX2 port map( A => n608, Y => n1463);
   U443 : NAND2X1 port map( A => n8, B => n1477, Y => n581);
   U444 : INVX2 port map( A => n581, Y => n1462);
   U445 : NAND2X1 port map( A => n8, B => n151, Y => n553);
   U446 : INVX2 port map( A => n553, Y => n1461);
   U447 : NAND2X1 port map( A => n8, B => n150, Y => n524);
   U448 : INVX2 port map( A => n524, Y => n1460);
   U450 : NAND2X1 port map( A => n8, B => n147, Y => n497);
   U451 : INVX2 port map( A => n497, Y => n1459);
   U454 : NAND2X1 port map( A => n105, B => n37, Y => n470);
   U455 : INVX2 port map( A => n470, Y => n1458);
   U456 : NAND2X1 port map( A => n105, B => n27, Y => n442);
   U457 : INVX2 port map( A => n442, Y => n1457);
   U458 : NAND2X1 port map( A => n29, B => n105, Y => n410);
   U459 : INVX2 port map( A => n410, Y => n1456);
   U460 : NAND2X1 port map( A => n33, B => n105, Y => n379);
   U461 : INVX2 port map( A => n379, Y => n1455);
   U462 : NAND2X1 port map( A => n11, B => n1477, Y => n349);
   U465 : INVX2 port map( A => n349, Y => n1454);
   U466 : NAND2X1 port map( A => n11, B => n151, Y => n318);
   U467 : INVX2 port map( A => n318, Y => n1453);
   U468 : NAND2X1 port map( A => n11, B => n150, Y => n283);
   U469 : INVX2 port map( A => n283, Y => n1452);
   U470 : NAND2X1 port map( A => n11, B => n147, Y => n246);
   U471 : INVX2 port map( A => n246, Y => n1451);
   U472 : NAND2X1 port map( A => n37, B => n14, Y => n152);
   U473 : INVX2 port map( A => n152, Y => n1450);
   U474 : NAND2X1 port map( A => n14, B => n27, Y => n159);
   U475 : INVX2 port map( A => n159, Y => n1449);
   U476 : INVX2 port map( A => RCV_DATA(2), Y => n1578);
   U477 : INVX2 port map( A => RCV_DATA(3), Y => n1577);
   U479 : INVX2 port map( A => RCV_DATA(5), Y => n1575);
   U480 : INVX2 port map( A => currentPlainKey_3_port, Y => n1570);
   U483 : INVX2 port map( A => currentPlainKey_2_port, Y => n1571);
   U484 : INVX2 port map( A => currentPlainKey_1_port, Y => n1572);
   U485 : NAND2X1 port map( A => n207, B => currentPlainKey_0_port, Y => n282);
   U486 : NAND2X1 port map( A => n175, B => RCV_DATA(5), Y => n1174);
   U487 : OAI21X1 port map( A => n23, B => n1364, C => n2, Y => n270);
   U488 : OAI21X1 port map( A => n1101, B => n23, C => n270, Y => n275);
   U489 : NAND2X1 port map( A => RCV_DATA(6), B => n85, Y => n327);
   U490 : MUX2X1 port map( B => n275, A => n327, S => n69, Y => n280);
   U491 : NAND2X1 port map( A => RCV_DATA(7), B => n175, Y => n1358);
   U494 : INVX2 port map( A => n1358, Y => n1370);
   U495 : NOR2X1 port map( A => n278, B => n277, Y => n279);
   U496 : MUX2X1 port map( B => n280, A => n222, S => n279, Y => n281);
   U497 : NAND2X1 port map( A => n282, B => n281, Y => n1332);
   U498 : NAND2X1 port map( A => n207, B => currentPlainKey_1_port, Y => n299);
   U499 : INVX2 port map( A => n1089, Y => n284);
   U500 : NAND2X1 port map( A => n9, B => n1477, Y => n319);
   U501 : INVX2 port map( A => n319, Y => n382);
   U502 : MUX2X1 port map( B => n284, A => n226, S => n382, Y => n286);
   U503 : NOR2X1 port map( A => n1578, B => n1011, Y => n285);
   U504 : AOI21X1 port map( A => n25, B => n286, C => n285, Y => n287);
   U505 : NOR2X1 port map( A => n287, B => n1364, Y => n289);
   U506 : AOI21X1 port map( A => n1479, B => n184, C => n289, Y => n291);
   U508 : NAND2X1 port map( A => n177, B => RCV_DATA(4), Y => n1172);
   U509 : MUX2X1 port map( B => n291, A => n1172, S => n1502, Y => n295);
   U512 : MUX2X1 port map( B => n295, A => n1367, S => n21, Y => n296);
   U513 : MUX2X1 port map( B => n296, A => n327, S => n23, Y => n297);
   U514 : MUX2X1 port map( B => n297, A => n224, S => n69, Y => n298);
   U515 : NAND2X1 port map( A => n299, B => n298, Y => n1331);
   U516 : NAND2X1 port map( A => n207, B => currentPlainKey_2_port, Y => n315);
   U517 : NOR2X1 port map( A => n1172, B => n300, Y => n311);
   U518 : NAND2X1 port map( A => n9, B => n143, Y => n347);
   U519 : NAND2X1 port map( A => n39, B => n87, Y => n336);
   U520 : INVX2 port map( A => n1077, Y => n301);
   U523 : OAI22X1 port map( A => n153, B => n347, C => n336, D => n301, Y => 
                           n303);
   U524 : OAI22X1 port map( A => n1011, B => n17, C => n137, D => n319, Y => 
                           n302);
   U525 : AOI21X1 port map( A => n25, B => n303, C => n302, Y => n304);
   U526 : MUX2X1 port map( B => n304, A => n1, S => n1502, Y => n305);
   U527 : NOR2X1 port map( A => n311, B => n305, Y => n312);
   U528 : MUX2X1 port map( B => n312, A => n327, S => n21, Y => n313);
   U529 : MUX2X1 port map( B => n313, A => n224, S => n23, Y => n314);
   U530 : NAND2X1 port map( A => n315, B => n314, Y => n1330);
   U531 : NAND2X1 port map( A => n207, B => currentPlainKey_3_port, Y => n334);
   U532 : NAND2X1 port map( A => n1479, B => n1367, Y => n326);
   U533 : INVX2 port map( A => n336, Y => n316);
   U534 : NAND2X1 port map( A => n1062, B => n316, Y => n317);
   U535 : NAND2X1 port map( A => n9, B => n151, Y => n348);
   U537 : INVX2 port map( A => n348, Y => n427);
   U538 : MUX2X1 port map( B => n317, A => n154, S => n427, Y => n321);
   U541 : OAI22X1 port map( A => n97, B => n319, C => n137, D => n347, Y => 
                           n320);
   U542 : OAI21X1 port map( A => n321, B => n320, C => n25, Y => n324);
   U543 : INVX2 port map( A => n1011, Y => n377);
   U544 : NAND2X1 port map( A => n195, B => n377, Y => n322);
   U545 : NAND3X1 port map( A => n326, B => n324, C => n322, Y => n330);
   U546 : MUX2X1 port map( B => n330, A => n217, S => n1502, Y => n331);
   U547 : MUX2X1 port map( B => n331, A => n1358, S => n21, Y => n332);
   U548 : NAND2X1 port map( A => n334, B => n333, Y => n1329);
   U549 : AOI22X1 port map( A => currentPlainKey_4_port, B => n207, C => n1479,
                           D => n209, Y => n346);
   U552 : NAND2X1 port map( A => n382, B => n192, Y => n343);
   U553 : OAI22X1 port map( A => n181, B => n347, C => n186, D => n348, Y => 
                           n338);
   U554 : NAND2X1 port map( A => n9, B => n1481, Y => n387);
   U555 : NAND2X1 port map( A => n348, B => n387, Y => n367);
   U556 : INVX2 port map( A => n367, Y => n425);
   U557 : NAND2X1 port map( A => n1046, B => n425, Y => n335);
   U558 : OAI22X1 port map( A => n153, B => n387, C => n336, D => n335, Y => 
                           n337);
   U559 : OAI21X1 port map( A => n338, B => n337, C => n25, Y => n340);
   U560 : NAND2X1 port map( A => n1367, B => n377, Y => n339);
   U561 : NAND3X1 port map( A => n343, B => n340, C => n339, Y => n344);
   U562 : MUX2X1 port map( B => n344, A => n224, S => n1502, Y => n345);
   U563 : NAND2X1 port map( A => n346, B => n345, Y => n1328);
   U564 : NAND2X1 port map( A => n1479, B => n224, Y => n365);
   U565 : INVX2 port map( A => n347, Y => n408);
   U567 : NAND2X1 port map( A => n408, B => n192, Y => n360);
   U568 : NOR2X1 port map( A => n180, B => n348, Y => n353);
   U571 : INVX2 port map( A => n1031, Y => n350);
   U572 : NAND3X1 port map( A => n425, B => n87, C => n350, Y => n351);
   U573 : OAI21X1 port map( A => n186, B => n387, C => n351, Y => n352);
   U574 : OAI21X1 port map( A => n353, B => n352, C => n39, Y => n357);
   U575 : NAND2X1 port map( A => n382, B => n1367, Y => n355);
   U576 : NAND3X1 port map( A => n360, B => n357, C => n355, Y => n361);
   U577 : NAND2X1 port map( A => n25, B => n361, Y => n364);
   U578 : AND2X2 port map( A => currentPlainKey_5_port, B => n207, Y => n362);
   U579 : AOI21X1 port map( A => n217, B => n377, C => n362, Y => n363);
   U582 : NAND3X1 port map( A => n365, B => n364, C => n363, Y => n1327);
   U583 : AOI22X1 port map( A => currentPlainKey_6_port, B => n206, C => n382, 
                           D => n209, Y => n381);
   U584 : NAND2X1 port map( A => n408, B => n1367, Y => n376);
   U585 : NAND2X1 port map( A => n9, B => n1478, Y => n397);
   U586 : INVX2 port map( A => n397, Y => n471);
   U587 : NAND2X1 port map( A => n471, B => n1136, Y => n369);
   U588 : NAND2X1 port map( A => n53, B => n87, Y => n399);
   U589 : INVX2 port map( A => n399, Y => n366);
   U590 : NAND2X1 port map( A => n1018, B => n366, Y => n368);
   U591 : AOI21X1 port map( A => n369, B => n368, C => n367, Y => n373);
   U592 : OAI22X1 port map( A => n181, B => n387, C => n968, D => n185, Y => 
                           n370);
   U593 : OAI21X1 port map( A => n373, B => n370, C => n39, Y => n375);
   U594 : NAND2X1 port map( A => n427, B => n192, Y => n374);
   U596 : NAND3X1 port map( A => n376, B => n375, C => n374, Y => n378);
   U597 : MUX2X1 port map( B => n378, A => n224, S => n377, Y => n380);
   U600 : NAND2X1 port map( A => n381, B => n380, Y => n1326);
   U601 : AOI22X1 port map( A => currentPlainKey_7_port, B => n206, C => n382, 
                           D => n219, Y => n396);
   U602 : NAND2X1 port map( A => n427, B => n1367, Y => n392);
   U603 : NOR2X1 port map( A => n968, B => n183, Y => n385);
   U604 : OAI22X1 port map( A => n187, B => n397, C => n1002, D => n399, Y => 
                           n383);
   U605 : OAI21X1 port map( A => n385, B => n383, C => n425, Y => n391);
   U606 : INVX2 port map( A => n387, Y => n443);
   U607 : NAND2X1 port map( A => n443, B => n192, Y => n390);
   U608 : NAND3X1 port map( A => n392, B => n391, C => n390, Y => n393);
   U611 : NAND2X1 port map( A => n39, B => n393, Y => n395);
   U612 : NAND2X1 port map( A => n408, B => n209, Y => n394);
   U613 : NAND3X1 port map( A => n396, B => n395, C => n394, Y => n1325);
   U614 : AOI22X1 port map( A => currentPlainKey_8_port, B => n207, C => n427, 
                           D => n209, Y => n412);
   U615 : NAND2X1 port map( A => n203, B => n1476, Y => n407);
   U616 : OAI22X1 port map( A => n181, B => n397, C => n941, D => n185, Y => 
                           n404);
   U617 : NAND2X1 port map( A => n9, B => n16, Y => n452);
   U618 : NAND2X1 port map( A => n941, B => n452, Y => n432);
   U619 : INVX2 port map( A => n432, Y => n486);
   U620 : NAND2X1 port map( A => n988, B => n486, Y => n398);
   U621 : OAI22X1 port map( A => n153, B => n452, C => n399, D => n398, Y => 
                           n400);
   U622 : OAI21X1 port map( A => n404, B => n400, C => n425, Y => n406);
   U623 : NAND2X1 port map( A => n443, B => n1367, Y => n405);
   U625 : NAND3X1 port map( A => n407, B => n406, C => n405, Y => n409);
   U626 : MUX2X1 port map( B => n409, A => n224, S => n408, Y => n411);
   U629 : NAND2X1 port map( A => n412, B => n411, Y => n1324);
   U630 : NAND2X1 port map( A => n443, B => n209, Y => n430);
   U631 : NAND2X1 port map( A => n471, B => n192, Y => n423);
   U632 : NOR2X1 port map( A => n941, B => n183, Y => n418);
   U633 : INVX2 port map( A => n973, Y => n413);
   U634 : NAND3X1 port map( A => n486, B => n87, C => n413, Y => n414);
   U635 : OAI21X1 port map( A => n187, B => n452, C => n414, Y => n416);
   U636 : OAI21X1 port map( A => n418, B => n416, C => n53, Y => n422);
   U637 : NAND2X1 port map( A => n1367, B => n1476, Y => n419);
   U640 : NAND3X1 port map( A => n423, B => n422, C => n419, Y => n424);
   U641 : NAND2X1 port map( A => n425, B => n424, Y => n429);
   U642 : AND2X2 port map( A => currentPlainKey_9_port, B => n205, Y => n426);
   U643 : AOI21X1 port map( A => n427, B => n221, C => n426, Y => n428);
   U644 : NAND3X1 port map( A => n430, B => n429, C => n428, Y => n1323);
   U645 : AOI22X1 port map( A => currentPlainKey_10_port, B => n207, C => n209,
                           D => n1476, Y => n446);
   U646 : NAND2X1 port map( A => n203, B => n1475, Y => n441);
   U647 : NAND2X1 port map( A => n107, B => n925, Y => n460);
   U648 : INVX2 port map( A => n460, Y => n534);
   U649 : NAND2X1 port map( A => n534, B => n1136, Y => n436);
   U650 : NAND2X1 port map( A => n45, B => n87, Y => n462);
   U651 : INVX2 port map( A => n462, Y => n431);
   U652 : NAND2X1 port map( A => n961, B => n431, Y => n435);
   U654 : AOI21X1 port map( A => n436, B => n435, C => n432, Y => n438);
   U655 : OAI22X1 port map( A => n181, B => n452, C => n914, D => n185, Y => 
                           n437);
   U656 : OAI21X1 port map( A => n438, B => n437, C => n53, Y => n440);
   U657 : NAND2X1 port map( A => n471, B => n1367, Y => n439);
   U660 : NAND3X1 port map( A => n441, B => n440, C => n439, Y => n444);
   U661 : MUX2X1 port map( B => n444, A => n224, S => n443, Y => n445);
   U662 : NAND2X1 port map( A => n446, B => n445, Y => n1322);
   U663 : AOI22X1 port map( A => currentPlainKey_11_port, B => n206, C => n219,
                           D => n1476, Y => n459);
   U664 : NAND2X1 port map( A => n1367, B => n1475, Y => n455);
   U665 : NOR2X1 port map( A => n914, B => n183, Y => n450);
   U666 : OAI22X1 port map( A => n187, B => n460, C => n946, D => n462, Y => 
                           n448);
   U667 : OAI21X1 port map( A => n450, B => n448, C => n486, Y => n454);
   U668 : INVX2 port map( A => n452, Y => n506);
   U671 : NAND2X1 port map( A => n506, B => n192, Y => n453);
   U673 : NAND3X1 port map( A => n455, B => n454, C => n453, Y => n456);
   U674 : NAND2X1 port map( A => n53, B => n456, Y => n458);
   U675 : NAND2X1 port map( A => n471, B => n209, Y => n457);
   U676 : NAND3X1 port map( A => n459, B => n458, C => n457, Y => n1321);
   U677 : AOI22X1 port map( A => currentPlainKey_12_port, B => n207, C => n209,
                           D => n1475, Y => n474);
   U678 : NAND2X1 port map( A => n203, B => n1474, Y => n469);
   U679 : OAI22X1 port map( A => n180, B => n460, C => n886, D => n185, Y => 
                           n466);
   U680 : NAND2X1 port map( A => n107, B => n20, Y => n512);
   U681 : NAND2X1 port map( A => n886, B => n512, Y => n494);
   U682 : INVX2 port map( A => n494, Y => n549);
   U683 : NAND2X1 port map( A => n934, B => n549, Y => n461);
   U684 : OAI22X1 port map( A => n153, B => n512, C => n462, D => n461, Y => 
                           n465);
   U685 : OAI21X1 port map( A => n466, B => n465, C => n486, Y => n468);
   U687 : NAND2X1 port map( A => n506, B => n1367, Y => n467);
   U688 : NAND3X1 port map( A => n469, B => n468, C => n467, Y => n472);
   U691 : MUX2X1 port map( B => n472, A => n224, S => n471, Y => n473);
   U692 : NAND2X1 port map( A => n474, B => n473, Y => n1320);
   U693 : NAND2X1 port map( A => n506, B => n209, Y => n492);
   U694 : NAND2X1 port map( A => n534, B => n192, Y => n484);
   U695 : NOR2X1 port map( A => n886, B => n183, Y => n481);
   U696 : INVX2 port map( A => n919, Y => n476);
   U697 : NAND3X1 port map( A => n549, B => n175, C => n476, Y => n479);
   U698 : OAI21X1 port map( A => n187, B => n512, C => n479, Y => n480);
   U699 : OAI21X1 port map( A => n481, B => n480, C => n45, Y => n483);
   U702 : NAND2X1 port map( A => n1367, B => n1474, Y => n482);
   U703 : NAND3X1 port map( A => n484, B => n483, C => n482, Y => n485);
   U704 : NAND2X1 port map( A => n486, B => n485, Y => n489);
   U705 : AND2X2 port map( A => currentPlainKey_13_port, B => n207, Y => n487);
   U706 : AOI21X1 port map( A => n221, B => n1475, C => n487, Y => n488);
   U707 : NAND3X1 port map( A => n492, B => n489, C => n488, Y => n1319);
   U708 : AOI22X1 port map( A => currentPlainKey_14_port, B => n207, C => n209,
                           D => n1474, Y => n509);
   U709 : NAND2X1 port map( A => n203, B => n1473, Y => n503);
   U710 : NAND2X1 port map( A => n107, B => n31, Y => n522);
   U711 : INVX2 port map( A => n522, Y => n595);
   U712 : NAND2X1 port map( A => n595, B => n1136, Y => n496);
   U713 : NAND2X1 port map( A => n47, B => n85, Y => n525);
   U714 : INVX2 port map( A => n525, Y => n493);
   U716 : NAND2X1 port map( A => n907, B => n493, Y => n495);
   U717 : AOI21X1 port map( A => n496, B => n495, C => n494, Y => n499);
   U720 : OAI22X1 port map( A => n97, B => n512, C => n857, D => n185, Y => 
                           n498);
   U721 : OAI21X1 port map( A => n499, B => n498, C => n45, Y => n501);
   U722 : NAND2X1 port map( A => n534, B => n1367, Y => n500);
   U723 : NAND3X1 port map( A => n503, B => n501, C => n500, Y => n507);
   U724 : MUX2X1 port map( B => n507, A => n224, S => n506, Y => n508);
   U725 : NAND2X1 port map( A => n509, B => n508, Y => n1318);
   U726 : AOI22X1 port map( A => currentPlainKey_15_port, B => n206, C => n219,
                           D => n1474, Y => n521);
   U727 : NAND2X1 port map( A => n1367, B => n1473, Y => n515);
   U728 : NOR2X1 port map( A => n857, B => n181, Y => n511);
   U731 : OAI22X1 port map( A => n187, B => n522, C => n891, D => n525, Y => 
                           n510);
   U732 : OAI21X1 port map( A => n511, B => n510, C => n549, Y => n514);
   U733 : INVX2 port map( A => n512, Y => n567);
   U734 : NAND2X1 port map( A => n567, B => n192, Y => n513);
   U735 : NAND3X1 port map( A => n515, B => n514, C => n513, Y => n516);
   U736 : NAND2X1 port map( A => n45, B => n516, Y => n520);
   U737 : NAND2X1 port map( A => n534, B => n209, Y => n519);
   U738 : NAND3X1 port map( A => n521, B => n520, C => n519, Y => n1317);
   U739 : AOI22X1 port map( A => currentPlainKey_16_port, B => n206, C => n210,
                           D => n1473, Y => n537);
   U740 : NAND2X1 port map( A => n203, B => n1472, Y => n533);
   U741 : OAI22X1 port map( A => n97, B => n522, C => n830, D => n186, Y => 
                           n527);
   U742 : NAND2X1 port map( A => n107, B => n35, Y => n573);
   U743 : NAND2X1 port map( A => n830, B => n573, Y => n556);
   U745 : INVX2 port map( A => n556, Y => n610);
   U746 : NAND2X1 port map( A => n877, B => n610, Y => n523);
   U749 : OAI22X1 port map( A => n154, B => n573, C => n525, D => n523, Y => 
                           n526);
   U750 : OAI21X1 port map( A => n527, B => n526, C => n549, Y => n530);
   U751 : NAND2X1 port map( A => n567, B => n1367, Y => n528);
   U752 : NAND3X1 port map( A => n533, B => n530, C => n528, Y => n535);
   U753 : MUX2X1 port map( B => n535, A => n224, S => n534, Y => n536);
   U754 : NAND2X1 port map( A => n537, B => n536, Y => n1316);
   U755 : NAND2X1 port map( A => n567, B => n209, Y => n554);
   U756 : NAND2X1 port map( A => n595, B => n192, Y => n547);
   U757 : NOR2X1 port map( A => n830, B => n181, Y => n541);
   U760 : INVX2 port map( A => n862, Y => n538);
   U761 : NAND3X1 port map( A => n610, B => n87, C => n538, Y => n539);
   U762 : OAI21X1 port map( A => n186, B => n573, C => n539, Y => n540);
   U763 : OAI21X1 port map( A => n541, B => n540, C => n47, Y => n543);
   U764 : NAND2X1 port map( A => n1367, B => n1472, Y => n542);
   U765 : NAND3X1 port map( A => n547, B => n543, C => n542, Y => n548);
   U766 : NAND2X1 port map( A => n549, B => n548, Y => n552);
   U767 : AND2X2 port map( A => currentPlainKey_17_port, B => n207, Y => n550);
   U768 : AOI21X1 port map( A => n221, B => n1473, C => n550, Y => n551);
   U769 : NAND3X1 port map( A => n554, B => n552, C => n551, Y => n1315);
   U770 : AOI22X1 port map( A => currentPlainKey_18_port, B => n206, C => n209,
                           D => n1472, Y => n570);
   U771 : NAND2X1 port map( A => n203, B => n1471, Y => n566);
   U772 : NAND2X1 port map( A => n10, B => n143, Y => n584);
   U774 : INVX2 port map( A => n584, Y => n657);
   U775 : NAND2X1 port map( A => n657, B => n1136, Y => n559);
   U778 : NAND2X1 port map( A => n55, B => n87, Y => n587);
   U779 : INVX2 port map( A => n587, Y => n555);
   U780 : NAND2X1 port map( A => n850, B => n555, Y => n557);
   U781 : AOI21X1 port map( A => n559, B => n557, C => n556, Y => n563);
   U782 : OAI22X1 port map( A => n180, B => n573, C => n803, D => n185, Y => 
                           n561);
   U783 : OAI21X1 port map( A => n563, B => n561, C => n47, Y => n565);
   U784 : NAND2X1 port map( A => n595, B => n1367, Y => n564);
   U785 : NAND3X1 port map( A => n566, B => n565, C => n564, Y => n568);
   U786 : MUX2X1 port map( B => n568, A => n223, S => n567, Y => n569);
   U789 : NAND2X1 port map( A => n570, B => n569, Y => n1314);
   U790 : AOI22X1 port map( A => currentPlainKey_19_port, B => n206, C => n219,
                           D => n1472, Y => n583);
   U791 : NAND2X1 port map( A => n1367, B => n1471, Y => n578);
   U792 : NOR2X1 port map( A => n803, B => n181, Y => n572);
   U793 : OAI22X1 port map( A => n187, B => n584, C => n835, D => n587, Y => 
                           n571);
   U794 : OAI21X1 port map( A => n572, B => n571, C => n610, Y => n577);
   U795 : INVX2 port map( A => n573, Y => n627);
   U796 : NAND2X1 port map( A => n627, B => n193, Y => n576);
   U797 : NAND3X1 port map( A => n578, B => n577, C => n576, Y => n579);
   U798 : NAND2X1 port map( A => n47, B => n579, Y => n582);
   U799 : NAND2X1 port map( A => n595, B => n210, Y => n580);
   U800 : NAND3X1 port map( A => n583, B => n582, C => n580, Y => n1313);
   U801 : AOI22X1 port map( A => currentPlainKey_20_port, B => n206, C => n210,
                           D => n1471, Y => n598);
   U802 : NAND2X1 port map( A => n203, B => n1470, Y => n594);
   U804 : OAI22X1 port map( A => n180, B => n584, C => n775, D => n186, Y => 
                           n591);
   U805 : NAND2X1 port map( A => n10, B => n1481, Y => n636);
   U808 : NAND2X1 port map( A => n775, B => n636, Y => n619);
   U809 : INVX2 port map( A => n619, Y => n672);
   U810 : NAND2X1 port map( A => n823, B => n672, Y => n585);
   U811 : OAI22X1 port map( A => n154, B => n636, C => n587, D => n585, Y => 
                           n590);
   U812 : OAI21X1 port map( A => n591, B => n590, C => n610, Y => n593);
   U813 : NAND2X1 port map( A => n627, B => n1367, Y => n592);
   U814 : NAND3X1 port map( A => n594, B => n593, C => n592, Y => n596);
   U815 : MUX2X1 port map( B => n596, A => n223, S => n595, Y => n597);
   U816 : NAND2X1 port map( A => n598, B => n597, Y => n1312);
   U819 : NAND2X1 port map( A => n627, B => n209, Y => n617);
   U820 : NAND2X1 port map( A => n657, B => n193, Y => n607);
   U821 : NOR2X1 port map( A => n775, B => n181, Y => n604);
   U822 : INVX2 port map( A => n808, Y => n599);
   U823 : NAND3X1 port map( A => n672, B => n87, C => n599, Y => n600);
   U824 : OAI21X1 port map( A => n187, B => n636, C => n600, Y => n603);
   U825 : OAI21X1 port map( A => n604, B => n603, C => n55, Y => n606);
   U826 : NAND2X1 port map( A => n1367, B => n1470, Y => n605);
   U827 : NAND3X1 port map( A => n607, B => n606, C => n605, Y => n609);
   U828 : NAND2X1 port map( A => n610, B => n609, Y => n614);
   U829 : AND2X2 port map( A => currentPlainKey_21_port, B => n207, Y => n611);
   U830 : AOI21X1 port map( A => n221, B => n1471, C => n611, Y => n612);
   U831 : NAND3X1 port map( A => n617, B => n614, C => n612, Y => n1311);
   U833 : AOI22X1 port map( A => currentPlainKey_22_port, B => n206, C => n210,
                           D => n1470, Y => n632);
   U834 : NAND2X1 port map( A => n197, B => n1469, Y => n626);
   U837 : NAND2X1 port map( A => n10, B => n1478, Y => n647);
   U838 : INVX2 port map( A => n647, Y => n717);
   U839 : NAND2X1 port map( A => n717, B => n1136, Y => n621);
   U840 : NAND2X1 port map( A => n57, B => n85, Y => n649);
   U841 : INVX2 port map( A => n649, Y => n618);
   U842 : NAND2X1 port map( A => n796, B => n618, Y => n620);
   U843 : AOI21X1 port map( A => n621, B => n620, C => n619, Y => n623);
   U844 : OAI22X1 port map( A => n180, B => n636, C => n746, D => n186, Y => 
                           n622);
   U845 : OAI21X1 port map( A => n623, B => n622, C => n55, Y => n625);
   U848 : NAND2X1 port map( A => n657, B => n1367, Y => n624);
   U849 : NAND3X1 port map( A => n626, B => n625, C => n624, Y => n630);
   U850 : MUX2X1 port map( B => n630, A => n223, S => n627, Y => n631);
   U851 : NAND2X1 port map( A => n632, B => n631, Y => n1310);
   U852 : AOI22X1 port map( A => currentPlainKey_23_port, B => n206, C => n219,
                           D => n1470, Y => n646);
   U853 : NAND2X1 port map( A => n1367, B => n1469, Y => n639);
   U854 : NOR2X1 port map( A => n746, B => n181, Y => n634);
   U855 : OAI22X1 port map( A => n187, B => n647, C => n780, D => n649, Y => 
                           n633);
   U856 : OAI21X1 port map( A => n634, B => n633, C => n672, Y => n638);
   U857 : INVX2 port map( A => n636, Y => n689);
   U858 : NAND2X1 port map( A => n689, B => n193, Y => n637);
   U859 : NAND3X1 port map( A => n639, B => n638, C => n637, Y => n641);
   U860 : NAND2X1 port map( A => n55, B => n641, Y => n645);
   U862 : NAND2X1 port map( A => n657, B => n1363, Y => n644);
   U863 : NAND3X1 port map( A => n646, B => n645, C => n644, Y => n1309);
   U866 : AOI22X1 port map( A => currentPlainKey_24_port, B => n206, C => n210,
                           D => n1469, Y => n660);
   U867 : NAND2X1 port map( A => n197, B => n1468, Y => n654);
   U868 : OAI22X1 port map( A => n97, B => n647, C => n719, D => n186, Y => 
                           n651);
   U869 : NAND2X1 port map( A => n10, B => n16, Y => n696);
   U870 : NAND2X1 port map( A => n719, B => n696, Y => n679);
   U871 : INVX2 port map( A => n679, Y => n733);
   U872 : NAND2X1 port map( A => n766, B => n733, Y => n648);
   U873 : OAI22X1 port map( A => n154, B => n696, C => n649, D => n648, Y => 
                           n650);
   U874 : OAI21X1 port map( A => n651, B => n650, C => n672, Y => n653);
   U877 : NAND2X1 port map( A => n689, B => n1367, Y => n652);
   U878 : NAND3X1 port map( A => n654, B => n653, C => n652, Y => n658);
   U879 : MUX2X1 port map( B => n658, A => n223, S => n657, Y => n659);
   U880 : NAND2X1 port map( A => n660, B => n659, Y => n1308);
   U881 : NAND2X1 port map( A => n689, B => n217, Y => n677);
   U882 : NAND2X1 port map( A => n717, B => n193, Y => n668);
   U883 : NOR2X1 port map( A => n719, B => n181, Y => n665);
   U884 : INVX2 port map( A => n751, Y => n661);
   U885 : NAND3X1 port map( A => n733, B => n175, C => n661, Y => n662);
   U886 : OAI21X1 port map( A => n187, B => n696, C => n662, Y => n663);
   U887 : OAI21X1 port map( A => n665, B => n663, C => n57, Y => n667);
   U888 : NAND2X1 port map( A => n1367, B => n1468, Y => n666);
   U889 : NAND3X1 port map( A => n668, B => n667, C => n666, Y => n670);
   U891 : NAND2X1 port map( A => n672, B => n670, Y => n676);
   U892 : AND2X2 port map( A => currentPlainKey_25_port, B => n206, Y => n674);
   U893 : AOI21X1 port map( A => n221, B => n1469, C => n674, Y => n675);
   U894 : NAND3X1 port map( A => n677, B => n676, C => n675, Y => n1307);
   U897 : AOI22X1 port map( A => currentPlainKey_26_port, B => n206, C => n210,
                           D => n1468, Y => n693);
   U898 : NAND2X1 port map( A => n197, B => n1467, Y => n688);
   U899 : NAND2X1 port map( A => n109, B => n925, Y => n707);
   U900 : INVX2 port map( A => n707, Y => n779);
   U901 : NAND2X1 port map( A => n779, B => n1136, Y => n681);
   U902 : NAND2X1 port map( A => n49, B => n87, Y => n709);
   U903 : INVX2 port map( A => n709, Y => n678);
   U904 : NAND2X1 port map( A => n739, B => n678, Y => n680);
   U905 : AOI21X1 port map( A => n681, B => n680, C => n679, Y => n683);
   U908 : OAI22X1 port map( A => n97, B => n696, C => n692, D => n186, Y => 
                           n682);
   U910 : OAI21X1 port map( A => n683, B => n682, C => n57, Y => n687);
   U911 : NAND2X1 port map( A => n717, B => n1367, Y => n684);
   U912 : NAND3X1 port map( A => n688, B => n687, C => n684, Y => n690);
   U913 : MUX2X1 port map( B => n690, A => n223, S => n689, Y => n691);
   U914 : NAND2X1 port map( A => n693, B => n691, Y => n1306);
   U915 : AOI22X1 port map( A => currentPlainKey_27_port, B => n206, C => n219,
                           D => n1468, Y => n706);
   U916 : NAND2X1 port map( A => n1367, B => n1467, Y => n702);
   U917 : NOR2X1 port map( A => n692, B => n183, Y => n695);
   U918 : OAI22X1 port map( A => n137, B => n707, C => n724, D => n709, Y => 
                           n694_port);
   U919 : OAI21X1 port map( A => n695, B => n694_port, C => n733, Y => n701);
   U920 : INVX2 port map( A => n696, Y => n750);
   U921 : NAND2X1 port map( A => n750, B => n192, Y => n698);
   U922 : NAND3X1 port map( A => n702, B => n701, C => n698, Y => n703);
   U924 : NAND2X1 port map( A => n57, B => n703, Y => n705);
   U925 : NAND2X1 port map( A => n717, B => n217, Y => n704);
   U928 : NAND3X1 port map( A => n706, B => n705, C => n704, Y => n1305);
   U929 : AOI22X1 port map( A => currentPlainKey_28_port, B => n205, C => n210,
                           D => n1467, Y => n721);
   U930 : NAND2X1 port map( A => n197, B => n1466, Y => n716);
   U931 : OAI22X1 port map( A => n180, B => n707, C => n664, D => n186, Y => 
                           n711);
   U932 : NAND2X1 port map( A => n109, B => n20, Y => n759);
   U933 : NAND2X1 port map( A => n664, B => n759, Y => n741);
   U934 : INVX2 port map( A => n741, Y => n794);
   U935 : NAND2X1 port map( A => n712, B => n794, Y => n708);
   U936 : OAI22X1 port map( A => n154, B => n759, C => n709, D => n708, Y => 
                           n710);
   U939 : OAI21X1 port map( A => n711, B => n710, C => n733, Y => n715);
   U940 : NAND2X1 port map( A => n750, B => n1367, Y => n714);
   U941 : NAND3X1 port map( A => n716, B => n715, C => n714, Y => n718);
   U942 : MUX2X1 port map( B => n718, A => n223, S => n717, Y => n720);
   U943 : NAND2X1 port map( A => n721, B => n720, Y => n1304);
   U944 : NAND2X1 port map( A => n750, B => n217, Y => n737);
   U945 : NAND2X1 port map( A => n779, B => n193, Y => n731);
   U946 : NOR2X1 port map( A => n664, B => n181, Y => n728);
   U947 : INVX2 port map( A => n697, Y => n722);
   U948 : NAND3X1 port map( A => n794, B => n85, C => n722, Y => n723);
   U949 : OAI21X1 port map( A => n187, B => n759, C => n723, Y => n725);
   U950 : OAI21X1 port map( A => n728, B => n725, C => n49, Y => n730);
   U951 : NAND2X1 port map( A => n1367, B => n1466, Y => n729);
   U953 : NAND3X1 port map( A => n731, B => n730, C => n729, Y => n732);
   U954 : NAND2X1 port map( A => n733, B => n732, Y => n736);
   U957 : AND2X2 port map( A => currentPlainKey_29_port, B => n207, Y => n734);
   U958 : AOI21X1 port map( A => n221, B => n1467, C => n734, Y => n735);
   U959 : NAND3X1 port map( A => n737, B => n736, C => n735, Y => n1303);
   U960 : AOI22X1 port map( A => currentPlainKey_30_port, B => n205, C => n217,
                           D => n1466, Y => n756);
   U961 : NAND2X1 port map( A => n197, B => n1465, Y => n749);
   U962 : NAND2X1 port map( A => n109, B => n31, Y => n770);
   U963 : INVX2 port map( A => n770, Y => n842);
   U964 : NAND2X1 port map( A => n842, B => n1136, Y => n743);
   U965 : NAND2X1 port map( A => n51, B => n87, Y => n772);
   U968 : INVX2 port map( A => n772, Y => n738);
   U969 : NAND2X1 port map( A => n685, B => n738, Y => n742);
   U970 : AOI21X1 port map( A => n743, B => n742, C => n741, Y => n745);
   U971 : OAI22X1 port map( A => n180, B => n759, C => n635, D => n185, Y => 
                           n744);
   U972 : OAI21X1 port map( A => n745, B => n744, C => n49, Y => n748);
   U973 : NAND2X1 port map( A => n779, B => n1367, Y => n747);
   U974 : NAND3X1 port map( A => n749, B => n748, C => n747, Y => n752);
   U975 : MUX2X1 port map( B => n752, A => n223, S => n750, Y => n755);
   U976 : NAND2X1 port map( A => n756, B => n755, Y => n1302);
   U977 : AOI22X1 port map( A => currentPlainKey_31_port, B => n205, C => n219,
                           D => n1466, Y => n769);
   U978 : NAND2X1 port map( A => n1367, B => n1465, Y => n762);
   U979 : NOR2X1 port map( A => n635, B => n181, Y => n758);
   U980 : OAI22X1 port map( A => n137, B => n770, C => n669, D => n772, Y => 
                           n757);
   U982 : OAI21X1 port map( A => n758, B => n757, C => n794, Y => n761);
   U983 : INVX2 port map( A => n759, Y => n814);
   U986 : NAND2X1 port map( A => n814, B => n195, Y => n760);
   U987 : NAND3X1 port map( A => n762, B => n761, C => n760, Y => n763);
   U988 : NAND2X1 port map( A => n49, B => n763, Y => n765);
   U989 : NAND2X1 port map( A => n779, B => n217, Y => n764);
   U990 : NAND3X1 port map( A => n769, B => n765, C => n764, Y => n1301);
   U991 : AOI22X1 port map( A => currentPlainKey_32_port, B => n205, C => n217,
                           D => n1465, Y => n785);
   U992 : NAND2X1 port map( A => n197, B => n1464, Y => n778);
   U993 : OAI22X1 port map( A => n97, B => n770, C => n608, D => n186, Y => 
                           n774);
   U994 : NAND2X1 port map( A => n109, B => n35, Y => n820);
   U997 : NAND2X1 port map( A => n608, B => n820, Y => n802);
   U998 : INVX2 port map( A => n802, Y => n856);
   U999 : NAND2X1 port map( A => n655, B => n856, Y => n771);
   U1000 : OAI22X1 port map( A => n154, B => n820, C => n772, D => n771, Y => 
                           n773);
   U1001 : OAI21X1 port map( A => n774, B => n773, C => n794, Y => n777);
   U1002 : NAND2X1 port map( A => n814, B => n1367, Y => n776);
   U1003 : NAND3X1 port map( A => n778, B => n777, C => n776, Y => n781);
   U1004 : MUX2X1 port map( B => n781, A => n223, S => n779, Y => n783);
   U1005 : NAND2X1 port map( A => n785, B => n783, Y => n1300);
   U1006 : NAND2X1 port map( A => n814, B => n217, Y => n800);
   U1007 : NAND2X1 port map( A => n842, B => n195, Y => n792);
   U1008 : NOR2X1 port map( A => n608, B => n181, Y => n789);
   U1009 : INVX2 port map( A => n640, Y => n786);
   U1011 : NAND3X1 port map( A => n856, B => n87, C => n786, Y => n787);
   U1012 : OAI21X1 port map( A => n187, B => n820, C => n787, Y => n788);
   U1013 : OAI21X1 port map( A => n789, B => n788, C => n51, Y => n791);
   U1016 : NAND2X1 port map( A => n1367, B => n1464, Y => n790);
   U1017 : NAND3X1 port map( A => n792, B => n791, C => n790, Y => n793);
   U1018 : NAND2X1 port map( A => n794, B => n793, Y => n799);
   U1019 : AND2X2 port map( A => currentPlainKey_33_port, B => n207, Y => n795)
                           ;
   U1020 : AOI21X1 port map( A => n221, B => n1465, C => n795, Y => n798);
   U1021 : NAND3X1 port map( A => n800, B => n799, C => n798, Y => n1299);
   U1022 : AOI22X1 port map( A => currentPlainKey_34_port, B => n205, C => n210
                           , D => n1464, Y => n817);
   U1023 : NAND2X1 port map( A => n197, B => n1463, Y => n813);
   U1024 : NAND2X1 port map( A => n8, B => n143, Y => n831);
   U1027 : INVX2 port map( A => n831, Y => n902);
   U1028 : NAND2X1 port map( A => n902, B => n1136, Y => n805);
   U1029 : NAND2X1 port map( A => n59, B => n175, Y => n833);
   U1030 : INVX2 port map( A => n833, Y => n801);
   U1031 : NAND2X1 port map( A => n628, B => n801, Y => n804);
   U1032 : AOI21X1 port map( A => n805, B => n804, C => n802, Y => n807);
   U1033 : OAI22X1 port map( A => n97, B => n820, C => n581, D => n186, Y => 
                           n806);
   U1034 : OAI21X1 port map( A => n807, B => n806, C => n51, Y => n812);
   U1035 : NAND2X1 port map( A => n842, B => n1367, Y => n809);
   U1036 : NAND3X1 port map( A => n813, B => n812, C => n809, Y => n815);
   U1037 : MUX2X1 port map( B => n815, A => n223, S => n814, Y => n816);
   U1038 : NAND2X1 port map( A => n817, B => n816, Y => n1298);
   U1039 : AOI22X1 port map( A => currentPlainKey_35_port, B => n205, C => n221
                           , D => n1464, Y => n829);
   U1040 : NAND2X1 port map( A => n1367, B => n1463, Y => n825);
   U1042 : NOR2X1 port map( A => n581, B => n181, Y => n819);
   U1043 : OAI22X1 port map( A => n137, B => n831, C => n613, D => n833, Y => 
                           n818);
   U1047 : OAI21X1 port map( A => n819, B => n818, C => n856, Y => n822);
   U1048 : INVX2 port map( A => n820, Y => n874);
   U1049 : NAND2X1 port map( A => n874, B => n193, Y => n821);
   U1050 : NAND3X1 port map( A => n825, B => n822, C => n821, Y => n826);
   U1051 : NAND2X1 port map( A => n51, B => n826, Y => n828);
   U1052 : NAND2X1 port map( A => n842, B => n217, Y => n827);
   U1053 : NAND3X1 port map( A => n829, B => n828, C => n827, Y => n1297);
   U1054 : AOI22X1 port map( A => currentPlainKey_36_port, B => n205, C => n217
                           , D => n1463, Y => n845);
   U1055 : NAND2X1 port map( A => n197, B => n1462, Y => n841);
   U1056 : OAI22X1 port map( A => n97, B => n831, C => n553, D => n186, Y => 
                           n836);
   U1060 : NAND2X1 port map( A => n8, B => n1481, Y => n882);
   U1061 : NAND2X1 port map( A => n553, B => n882, Y => n866);
   U1062 : INVX2 port map( A => n866, Y => n917);
   U1063 : NAND2X1 port map( A => n601, B => n917, Y => n832);
   U1064 : OAI22X1 port map( A => n154, B => n882, C => n833, D => n832, Y => 
                           n834);
   U1065 : OAI21X1 port map( A => n836, B => n834, C => n856, Y => n840);
   U1066 : NAND2X1 port map( A => n874, B => n1367, Y => n839);
   U1067 : NAND3X1 port map( A => n841, B => n840, C => n839, Y => n843);
   U1068 : MUX2X1 port map( B => n843, A => n223, S => n842, Y => n844);
   U1069 : NAND2X1 port map( A => n845, B => n844, Y => n1296);
   U1070 : NAND2X1 port map( A => n874, B => n217, Y => n861);
   U1071 : NAND2X1 port map( A => n902, B => n195, Y => n854);
   U1072 : NOR2X1 port map( A => n553, B => n183, Y => n849);
   U1073 : INVX2 port map( A => n586, Y => n846);
   U1075 : NAND3X1 port map( A => n917, B => n87, C => n846, Y => n847);
   U1076 : OAI21X1 port map( A => n185, B => n882, C => n847, Y => n848);
   U1080 : OAI21X1 port map( A => n849, B => n848, C => n59, Y => n853);
   U1081 : NAND2X1 port map( A => n1367, B => n1462, Y => n852);
   U1082 : NAND3X1 port map( A => n854, B => n853, C => n852, Y => n855);
   U1083 : NAND2X1 port map( A => n856, B => n855, Y => n860);
   U1084 : AND2X2 port map( A => currentPlainKey_37_port, B => n207, Y => n858)
                           ;
   U1085 : AOI21X1 port map( A => n222, B => n1463, C => n858, Y => n859);
   U1086 : NAND3X1 port map( A => n861, B => n860, C => n859, Y => n1295);
   U1087 : AOI22X1 port map( A => currentPlainKey_38_port, B => n205, C => n210
                           , D => n1462, Y => n879);
   U1088 : NAND2X1 port map( A => n197, B => n1461, Y => n873);
   U1089 : NAND2X1 port map( A => n8, B => n1478, Y => n892);
   U1093 : INVX2 port map( A => n892, Y => n965);
   U1094 : NAND2X1 port map( A => n965, B => n1136, Y => n868);
   U1095 : NAND2X1 port map( A => n61, B => n175, Y => n896);
   U1096 : INVX2 port map( A => n896, Y => n863);
   U1097 : NAND2X1 port map( A => n574, B => n863, Y => n867);
   U1098 : AOI21X1 port map( A => n868, B => n867, C => n866, Y => n870);
   U1099 : OAI22X1 port map( A => n180, B => n882, C => n524, D => n186, Y => 
                           n869);
   U1100 : OAI21X1 port map( A => n870, B => n869, C => n59, Y => n872);
   U1101 : NAND2X1 port map( A => n902, B => n1367, Y => n871);
   U1102 : NAND3X1 port map( A => n873, B => n872, C => n871, Y => n875);
   U1103 : MUX2X1 port map( B => n875, A => n223, S => n874, Y => n876);
   U1104 : NAND2X1 port map( A => n879, B => n876, Y => n1294);
   U1105 : AOI22X1 port map( A => currentPlainKey_39_port, B => n205, C => n219
                           , D => n1462, Y => n890);
   U1106 : NAND2X1 port map( A => n1367, B => n1461, Y => n885);
   U1107 : NOR2X1 port map( A => n524, B => n183, Y => n881);
   U1108 : OAI22X1 port map( A => n187, B => n892, C => n558, D => n896, Y => 
                           n880);
   U1109 : OAI21X1 port map( A => n881, B => n880, C => n917, Y => n884);
   U1110 : INVX2 port map( A => n882, Y => n937);
   U1114 : NAND2X1 port map( A => n937, B => n195, Y => n883);
   U1115 : NAND3X1 port map( A => n885, B => n884, C => n883, Y => n887);
   U1116 : NAND2X1 port map( A => n59, B => n887, Y => n889);
   U1117 : NAND2X1 port map( A => n902, B => n217, Y => n888);
   U1118 : NAND3X1 port map( A => n890, B => n889, C => n888, Y => n1293);
   U1119 : AOI22X1 port map( A => currentPlainKey_40_port, B => n205, C => n210
                           , D => n1461, Y => n905);
   U1120 : NAND2X1 port map( A => n197, B => n1460, Y => n901);
   U1121 : OAI22X1 port map( A => n180, B => n892, C => n497, D => n186, Y => 
                           n898);
   U1122 : NAND2X1 port map( A => n8, B => n16, Y => n944);
   U1123 : NAND2X1 port map( A => n497, B => n944, Y => n927);
   U1124 : INVX2 port map( A => n927, Y => n981);
   U1125 : NAND2X1 port map( A => n544, B => n981, Y => n894);
   U1129 : OAI22X1 port map( A => n154, B => n944, C => n896, D => n894, Y => 
                           n897);
   U1130 : OAI21X1 port map( A => n898, B => n897, C => n917, Y => n900);
   U1131 : NAND2X1 port map( A => n937, B => n1367, Y => n899);
   U1132 : NAND3X1 port map( A => n901, B => n900, C => n899, Y => n903);
   U1133 : MUX2X1 port map( B => n903, A => n223, S => n902, Y => n904);
   U1134 : NAND2X1 port map( A => n905, B => n904, Y => n1292);
   U1135 : NAND2X1 port map( A => n937, B => n217, Y => n924);
   U1136 : NAND2X1 port map( A => n965, B => n193, Y => n915);
   U1137 : NOR2X1 port map( A => n497, B => n183, Y => n911);
   U1138 : INVX2 port map( A => n529, Y => n906);
   U1139 : NAND3X1 port map( A => n981, B => n87, C => n906, Y => n909);
   U1140 : OAI21X1 port map( A => n187, B => n944, C => n909, Y => n910);
   U1141 : OAI21X1 port map( A => n911, B => n910, C => n61, Y => n913);
   U1142 : NAND2X1 port map( A => n1367, B => n1460, Y => n912);
   U1143 : NAND3X1 port map( A => n915, B => n913, C => n912, Y => n916);
   U1144 : NAND2X1 port map( A => n917, B => n916, Y => n923);
   U1145 : AND2X2 port map( A => currentPlainKey_41_port, B => n207, Y => n918)
                           ;
   U1146 : AOI21X1 port map( A => n222, B => n1461, C => n918, Y => n920);
   U1147 : NAND3X1 port map( A => n924, B => n923, C => n920, Y => n1291);
   U1148 : AOI22X1 port map( A => currentPlainKey_42_port, B => n205, C => n210
                           , D => n1460, Y => n940);
   U1149 : NAND2X1 port map( A => n197, B => n1459, Y => n936);
   U1150 : NAND2X1 port map( A => n105, B => n925, Y => n955);
   U1151 : INVX2 port map( A => n955, Y => n1026);
   U1152 : NAND2X1 port map( A => n1026, B => n1136, Y => n929);
   U1153 : NAND2X1 port map( A => n43, B => n87, Y => n957);
   U1158 : INVX2 port map( A => n957, Y => n926);
   U1159 : NAND2X1 port map( A => n517, B => n926, Y => n928);
   U1160 : AOI21X1 port map( A => n929, B => n928, C => n927, Y => n931);
   U1161 : OAI22X1 port map( A => n97, B => n944, C => n470, D => n186, Y => 
                           n930);
   U1162 : OAI21X1 port map( A => n931, B => n930, C => n61, Y => n933);
   U1163 : NAND2X1 port map( A => n965, B => n1367, Y => n932);
   U1164 : NAND3X1 port map( A => n936, B => n933, C => n932, Y => n938);
   U1165 : MUX2X1 port map( B => n938, A => n222, S => n937, Y => n939);
   U1166 : NAND2X1 port map( A => n940, B => n939, Y => n1290);
   U1167 : AOI22X1 port map( A => currentPlainKey_43_port, B => n205, C => n221
                           , D => n1460, Y => n954);
   U1168 : NAND2X1 port map( A => n1367, B => n1459, Y => n950);
   U1169 : NOR2X1 port map( A => n470, B => n183, Y => n943);
   U1170 : OAI22X1 port map( A => n187, B => n955, C => n502, D => n957, Y => 
                           n942);
   U1171 : OAI21X1 port map( A => n943, B => n942, C => n981, Y => n947);
   U1172 : INVX2 port map( A => n944, Y => n998);
   U1173 : NAND2X1 port map( A => n998, B => n195, Y => n945);
   U1174 : NAND3X1 port map( A => n950, B => n947, C => n945, Y => n951);
   U1175 : NAND2X1 port map( A => n61, B => n951, Y => n953);
   U1176 : NAND2X1 port map( A => n965, B => n217, Y => n952);
   U1177 : NAND3X1 port map( A => n954, B => n953, C => n952, Y => n1289);
   U1178 : AOI22X1 port map( A => currentPlainKey_44_port, B => n205, C => n210
                           , D => n1459, Y => n969);
   U1179 : NAND2X1 port map( A => n195, B => n1458, Y => n964);
   U1180 : OAI22X1 port map( A => n97, B => n955, C => n442, D => n185, Y => 
                           n959);
   U1181 : NAND2X1 port map( A => n105, B => n20, Y => n1007);
   U1188 : NAND2X1 port map( A => n442, B => n1007, Y => n987);
   U1191 : INVX2 port map( A => n987, Y => n1042);
   U1192 : NAND2X1 port map( A => n490, B => n1042, Y => n956);
   U1193 : OAI22X1 port map( A => n154, B => n1007, C => n957, D => n956, Y => 
                           n958);
   U1194 : OAI21X1 port map( A => n959, B => n958, C => n981, Y => n963);
   U1195 : NAND2X1 port map( A => n998, B => n1367, Y => n960);
   U1196 : NAND3X1 port map( A => n964, B => n963, C => n960, Y => n966);
   U1197 : MUX2X1 port map( B => n966, A => n222, S => n965, Y => n967);
   U1198 : NAND2X1 port map( A => n969, B => n967, Y => n1288);
   U1200 : NAND2X1 port map( A => n998, B => n210, Y => n985);
   U1201 : NAND2X1 port map( A => n1026, B => n193, Y => n979);
   U1202 : NOR2X1 port map( A => n442, B => n183, Y => n974);
   U1203 : INVX2 port map( A => n475, Y => n970);
   U1204 : NAND3X1 port map( A => n1042, B => n87, C => n970, Y => n971);
   U1205 : OAI21X1 port map( A => n185, B => n1007, C => n971, Y => n972);
   U1206 : OAI21X1 port map( A => n974, B => n972, C => n43, Y => n978);
   U1207 : NAND2X1 port map( A => n1367, B => n1458, Y => n977);
   U1208 : NAND3X1 port map( A => n979, B => n978, C => n977, Y => n980);
   U1209 : NAND2X1 port map( A => n981, B => n980, Y => n984);
   U1210 : AND2X2 port map( A => currentPlainKey_45_port, B => n206, Y => n982)
                           ;
   U1211 : AOI21X1 port map( A => n221, B => n1459, C => n982, Y => n983);
   U1212 : NAND3X1 port map( A => n985, B => n984, C => n983, Y => n1287);
   U1213 : AOI22X1 port map( A => currentPlainKey_46_port, B => n206, C => n210
                           , D => n1458, Y => n1001);
   U1214 : NAND2X1 port map( A => n195, B => n1457, Y => n997);
   U1215 : NAND2X1 port map( A => n31, B => n105, Y => n1016);
   U1216 : INVX2 port map( A => n1016, Y => n1084);
   U1217 : NAND2X1 port map( A => n1084, B => n1136, Y => n992);
   U1218 : NAND2X1 port map( A => n41, B => n87, Y => n1020);
   U1219 : INVX2 port map( A => n1020, Y => n986);
   U1221 : NAND2X1 port map( A => n463, B => n986, Y => n991);
   U1222 : AOI21X1 port map( A => n992, B => n991, C => n987, Y => n994);
   U1223 : OAI22X1 port map( A => n180, B => n1007, C => n410, D => n185, Y => 
                           n993);
   U1224 : OAI21X1 port map( A => n994, B => n993, C => n43, Y => n996);
   U1225 : NAND2X1 port map( A => n1026, B => n1367, Y => n995);
   U1226 : NAND3X1 port map( A => n997, B => n996, C => n995, Y => n999);
   U1227 : MUX2X1 port map( B => n999, A => n222, S => n998, Y => n1000);
   U1228 : NAND2X1 port map( A => n1001, B => n1000, Y => n1286);
   U1229 : AOI22X1 port map( A => currentPlainKey_47_port, B => n206, C => n219
                           , D => n1458, Y => n1015);
   U1230 : NAND2X1 port map( A => n1367, B => n1457, Y => n1010);
   U1231 : NOR2X1 port map( A => n410, B => n183, Y => n1005);
   U1232 : OAI22X1 port map( A => n187, B => n1016, C => n447, D => n1020, Y =>
                           n1003);
   U1233 : OAI21X1 port map( A => n1005, B => n1003, C => n1042, Y => n1009);
   U1234 : INVX2 port map( A => n1007, Y => n1058);
   U1235 : NAND2X1 port map( A => n1058, B => n193, Y => n1008);
   U1236 : NAND3X1 port map( A => n1010, B => n1009, C => n1008, Y => n1012);
   U1237 : NAND2X1 port map( A => n43, B => n1012, Y => n1014);
   U1238 : NAND2X1 port map( A => n1026, B => n1363, Y => n1013);
   U1239 : NAND3X1 port map( A => n1015, B => n1014, C => n1013, Y => n1285);
   U1240 : AOI22X1 port map( A => currentPlainKey_48_port, B => n205, C => n210
                           , D => n1457, Y => n1029);
   U1241 : NAND2X1 port map( A => n195, B => n1456, Y => n1025);
   U1242 : OAI22X1 port map( A => n180, B => n1016, C => n379, D => n185, Y => 
                           n1022);
   U1243 : NAND2X1 port map( A => n105, B => n35, Y => n1066);
   U1244 : NAND2X1 port map( A => n379, B => n1066, Y => n1050);
   U1245 : INVX2 port map( A => n1050, Y => n1098);
   U1246 : NAND2X1 port map( A => n433, B => n1098, Y => n1017);
   U1247 : OAI22X1 port map( A => n154, B => n1066, C => n1020, D => n1017, Y 
                           => n1021);
   U1248 : OAI21X1 port map( A => n1022, B => n1021, C => n1042, Y => n1024);
   U1249 : NAND2X1 port map( A => n1058, B => n1367, Y => n1023);
   U1250 : NAND3X1 port map( A => n1025, B => n1024, C => n1023, Y => n1027);
   U1251 : MUX2X1 port map( B => n1027, A => n222, S => n1026, Y => n1028);
   U1252 : NAND2X1 port map( A => n1029, B => n1028, Y => n1284);
   U1253 : NAND2X1 port map( A => n1058, B => n210, Y => n1048);
   U1254 : NAND2X1 port map( A => n1084, B => n193, Y => n1040);
   U1255 : NOR2X1 port map( A => n379, B => n183, Y => n1036);
   U1256 : INVX2 port map( A => n415, Y => n1030);
   U1257 : NAND3X1 port map( A => n1098, B => n87, C => n1030, Y => n1032);
   U1258 : OAI21X1 port map( A => n186, B => n1066, C => n1032, Y => n1035);
   U1259 : OAI21X1 port map( A => n1036, B => n1035, C => n41, Y => n1039);
   U1260 : NAND2X1 port map( A => n1367, B => n1456, Y => n1037);
   U1261 : NAND3X1 port map( A => n1040, B => n1039, C => n1037, Y => n1041);
   U1262 : NAND2X1 port map( A => n1042, B => n1041, Y => n1045);
   U1263 : AND2X2 port map( A => currentPlainKey_49_port, B => n207, Y => n1043
                           );
   U1264 : AOI21X1 port map( A => n221, B => n1457, C => n1043, Y => n1044);
   U1265 : NAND3X1 port map( A => n1048, B => n1045, C => n1044, Y => n1283);
   U1266 : AOI22X1 port map( A => currentPlainKey_50_port, B => n206, C => n209
                           , D => n1456, Y => n1061);
   U1267 : NAND2X1 port map( A => n197, B => n1455, Y => n1057);
   U1268 : NAND2X1 port map( A => n11, B => n143, Y => n1074);
   U1269 : INVX2 port map( A => n1074, Y => n1146);
   U1270 : NAND2X1 port map( A => n1146, B => n1136, Y => n1052);
   U1271 : NAND2X1 port map( A => n63, B => n87, Y => n1076);
   U1272 : INVX2 port map( A => n1076, Y => n1049);
   U1275 : NAND2X1 port map( A => n401, B => n1049, Y => n1051);
   U1276 : AOI21X1 port map( A => n1052, B => n1051, C => n1050, Y => n1054);
   U1277 : OAI22X1 port map( A => n97, B => n1066, C => n349, D => n185, Y => 
                           n1053);
   U1278 : OAI21X1 port map( A => n1054, B => n1053, C => n41, Y => n1056);
   U1279 : NAND2X1 port map( A => n1084, B => n1367, Y => n1055);
   U1280 : NAND3X1 port map( A => n1057, B => n1056, C => n1055, Y => n1059);
   U1281 : MUX2X1 port map( B => n1059, A => n222, S => n1058, Y => n1060);
   U1282 : NAND2X1 port map( A => n1061, B => n1060, Y => n1282);
   U1283 : AOI22X1 port map( A => currentPlainKey_51_port, B => n205, C => n219
                           , D => n1456, Y => n1073);
   U1284 : NAND2X1 port map( A => n1367, B => n1455, Y => n1069);
   U1285 : NOR2X1 port map( A => n349, B => n183, Y => n1065);
   U1286 : OAI22X1 port map( A => n187, B => n1074, C => n384, D => n1076, Y =>
                           n1064);
   U1287 : OAI21X1 port map( A => n1065, B => n1064, C => n1098, Y => n1068);
   U1288 : INVX2 port map( A => n1066, Y => n1118);
   U1289 : NAND2X1 port map( A => n1118, B => n193, Y => n1067);
   U1290 : NAND3X1 port map( A => n1069, B => n1068, C => n1067, Y => n1070);
   U1291 : NAND2X1 port map( A => n41, B => n1070, Y => n1072);
   U1292 : NAND2X1 port map( A => n1084, B => n217, Y => n1071);
   U1293 : NAND3X1 port map( A => n1073, B => n1072, C => n1071, Y => n1281);
   U1294 : AOI22X1 port map( A => currentPlainKey_52_port, B => n205, C => n209
                           , D => n1455, Y => n1087);
   U1295 : NAND2X1 port map( A => n195, B => n1454, Y => n1083);
   U1296 : OAI22X1 port map( A => n180, B => n1074, C => n318, D => n185, Y => 
                           n1080);
   U1297 : NAND2X1 port map( A => n11, B => n1481, Y => n1122);
   U1298 : NAND2X1 port map( A => n318, B => n1122, Y => n1110);
   U1299 : INVX2 port map( A => n1110, Y => n1157);
   U1300 : NAND2X1 port map( A => n371, B => n1157, Y => n1075);
   U1301 : OAI22X1 port map( A => n1122, B => n153, C => n1076, D => n1075, Y 
                           => n1079);
   U1302 : OAI21X1 port map( A => n1080, B => n1079, C => n1098, Y => n1082);
   U1303 : NAND2X1 port map( A => n1118, B => n1367, Y => n1081);
   U1304 : NAND3X1 port map( A => n1083, B => n1082, C => n1081, Y => n1085);
   U1306 : MUX2X1 port map( B => n1085, A => n222, S => n1084, Y => n1086);
   U1307 : NAND2X1 port map( A => n1087, B => n1086, Y => n1280);
   U1308 : NAND2X1 port map( A => n1118, B => n209, Y => n1109);
   U1309 : NAND2X1 port map( A => n1146, B => n193, Y => n1096);
   U1310 : NOR2X1 port map( A => n318, B => n183, Y => n1093);
   U1311 : INVX2 port map( A => n354, Y => n1088);
   U1312 : NAND3X1 port map( A => n1157, B => n175, C => n1088, Y => n1091);
   U1313 : OAI21X1 port map( A => n185, B => n1122, C => n1091, Y => n1092);
   U1316 : OAI21X1 port map( A => n1093, B => n1092, C => n63, Y => n1095);
   U1317 : NAND2X1 port map( A => n1367, B => n1454, Y => n1094);
   U1318 : NAND3X1 port map( A => n1096, B => n1095, C => n1094, Y => n1097);
   U1319 : NAND2X1 port map( A => n1098, B => n1097, Y => n1102);
   U1320 : AND2X2 port map( A => currentPlainKey_53_port, B => n205, Y => n1099
                           );
   U1321 : AOI21X1 port map( A => n221, B => n1455, C => n1099, Y => n1100);
   U1322 : NAND3X1 port map( A => n1109, B => n1102, C => n1100, Y => n1279);
   U1323 : AOI22X1 port map( A => currentPlainKey_54_port, B => n207, C => n209
                           , D => n1454, Y => n1121);
   U1324 : NAND2X1 port map( A => n195, B => n1453, Y => n1117);
   U1325 : NAND2X1 port map( A => n11, B => n1478, Y => n1125);
   U1326 : NAND2X1 port map( A => n283, B => n1125, Y => n1138);
   U1327 : INVX2 port map( A => n1138, Y => n1177);
   U1328 : NAND3X1 port map( A => n341, B => n87, C => n1177, Y => n1112);
   U1329 : INVX2 port map( A => n1125, Y => n1193);
   U1330 : NAND2X1 port map( A => n1136, B => n1193, Y => n1111);
   U1331 : AOI21X1 port map( A => n1112, B => n1111, C => n1110, Y => n1114);
   U1332 : OAI22X1 port map( A => n283, B => n137, C => n97, D => n1122, Y => 
                           n1113);
   U1333 : OAI21X1 port map( A => n1114, B => n1113, C => n63, Y => n1116);
   U1334 : NAND2X1 port map( A => n1146, B => n1367, Y => n1115);
   U1335 : NAND3X1 port map( A => n1117, B => n1116, C => n1115, Y => n1119);
   U1336 : MUX2X1 port map( B => n1119, A => n222, S => n1118, Y => n1120);
   U1337 : NAND2X1 port map( A => n1121, B => n1120, Y => n1278);
   U1338 : NAND2X1 port map( A => n1146, B => n209, Y => n1135);
   U1339 : INVX2 port map( A => n1122, Y => n1168);
   U1340 : NAND2X1 port map( A => n1168, B => n192, Y => n1130);
   U1341 : NOR2X1 port map( A => n283, B => n183, Y => n1127);
   U1342 : INVX2 port map( A => n323, Y => n1123);
   U1343 : NAND3X1 port map( A => n1177, B => n175, C => n1123, Y => n1124);
   U1344 : OAI21X1 port map( A => n1125, B => n137, C => n1124, Y => n1126);
   U1345 : OAI21X1 port map( A => n1127, B => n1126, C => n1157, Y => n1129);
   U1346 : NAND2X1 port map( A => n1367, B => n1453, Y => n1128);
   U1347 : NAND3X1 port map( A => n1130, B => n1129, C => n1128, Y => n1131);
   U1348 : NAND2X1 port map( A => n63, B => n1131, Y => n1134);
   U1349 : AND2X2 port map( A => currentPlainKey_55_port, B => n207, Y => n1132
                           );
   U1350 : AOI21X1 port map( A => n221, B => n1454, C => n1132, Y => n1133);
   U1351 : NAND3X1 port map( A => n1135, B => n1134, C => n1133, Y => n1277);
   U1352 : AOI22X1 port map( A => currentPlainKey_56_port, B => n206, C => n209
                           , D => n1453, Y => n1149);
   U1353 : NAND2X1 port map( A => n195, B => n1452, Y => n1145);
   U1354 : NAND2X1 port map( A => n11, B => n16, Y => n1173);
   U1355 : NAND3X1 port map( A => n87, B => n1173, C => n246, Y => n1150);
   U1356 : INVX2 port map( A => n1150, Y => n1263);
   U1357 : INVX2 port map( A => n1173, Y => n1357);
   U1358 : AOI22X1 port map( A => n306, B => n1263, C => n1136, D => n1357, Y 
                           => n1139);
   U1359 : AOI22X1 port map( A => n184, B => n1193, C => n188, D => n1451, Y =>
                           n1137);
   U1360 : OAI21X1 port map( A => n1139, B => n1138, C => n1137, Y => n1140);
   U1361 : NAND2X1 port map( A => n1157, B => n1140, Y => n1142);
   U1362 : NAND2X1 port map( A => n1168, B => n1367, Y => n1141);
   U1363 : NAND3X1 port map( A => n1145, B => n1142, C => n1141, Y => n1147);
   U1364 : MUX2X1 port map( B => n1147, A => n222, S => n1146, Y => n1148);
   U1365 : NAND2X1 port map( A => n1149, B => n1148, Y => n1276);
   U1366 : AOI22X1 port map( A => currentPlainKey_57_port, B => n206, C => n219
                           , D => n1453, Y => n1161);
   U1367 : NAND2X1 port map( A => n1367, B => n1452, Y => n1155);
   U1368 : NOR2X1 port map( A => n288, B => n1150, Y => n1152);
   U1369 : OAI22X1 port map( A => n246, B => n97, C => n1173, D => n185, Y => 
                           n1151);
   U1370 : OAI21X1 port map( A => n1152, B => n1151, C => n1177, Y => n1154);
   U1371 : NAND2X1 port map( A => n1193, B => n192, Y => n1153);
   U1372 : NAND3X1 port map( A => n1155, B => n1154, C => n1153, Y => n1156);
   U1373 : NAND2X1 port map( A => n1157, B => n1156, Y => n1159);
   U1374 : NAND2X1 port map( A => n1168, B => n210, Y => n1158);
   U1375 : NAND3X1 port map( A => n1161, B => n1159, C => n1158, Y => n1275);
   U1376 : AOI22X1 port map( A => currentPlainKey_58_port, B => n205, C => n209
                           , D => n1452, Y => n1171);
   U1377 : NAND2X1 port map( A => n195, B => n1451, Y => n1167);
   U1378 : NAND2X1 port map( A => n1263, B => n152, Y => n1187);
   U1379 : INVX2 port map( A => n272, Y => n1162);
   U1380 : OAI22X1 port map( A => n152, B => n137, C => n1173, D => n180, Y => 
                           n1163);
   U1381 : OAI21X1 port map( A => n1164, B => n1163, C => n1177, Y => n1166);
   U1382 : NAND2X1 port map( A => n1193, B => n1367, Y => n1165);
   U1383 : NAND3X1 port map( A => n1167, B => n1166, C => n1165, Y => n1169);
   U1384 : MUX2X1 port map( B => n1169, A => n222, S => n1168, Y => n1170);
   U1385 : NAND2X1 port map( A => n1171, B => n1170, Y => n1274);
   U1386 : AOI22X1 port map( A => currentPlainKey_59_port, B => n205, C => n219
                           , D => n1452, Y => n1183);
   U1387 : OAI22X1 port map( A => n246, B => n4, C => n1173, D => n1172, Y => 
                           n1180);
   U1388 : INVX2 port map( A => n251, Y => n1176);
   U1389 : NAND3X1 port map( A => RCV_DATA(3), B => n1450, C => n1263, Y => 
                           n1175);
   U1390 : OAI21X1 port map( A => n1187, B => n1176, C => n1175, Y => n1179);
   U1391 : OAI21X1 port map( A => n1180, B => n1179, C => n1177, Y => n1182);
   U1392 : NAND2X1 port map( A => n1193, B => n210, Y => n1181);
   U1393 : NAND3X1 port map( A => n1183, B => n1182, C => n1181, Y => n1273);
   U1394 : AOI22X1 port map( A => currentPlainKey_60_port, B => n207, C => n209
                           , D => n1451, Y => n1196);
   U1395 : NAND2X1 port map( A => n197, B => n1450, Y => n1192);
   U1396 : AOI22X1 port map( A => n1497, B => RCV_DATA(3), C => n1449, D => 
                           RCV_DATA(2), Y => n1185);
   U1397 : OAI21X1 port map( A => n226, B => n164, C => n1185, Y => n1189);
   U1398 : INVX2 port map( A => n1187, Y => n1188);
   U1399 : OAI21X1 port map( A => n67, B => n1189, C => n1188, Y => n1191);
   U1400 : NAND2X1 port map( A => n1367, B => n1357, Y => n1190);
   U1401 : NAND3X1 port map( A => n1192, B => n1191, C => n1190, Y => n1194);
   U1402 : MUX2X1 port map( B => n1194, A => n222, S => n1193, Y => n1195);
   U1403 : NAND2X1 port map( A => n1196, B => n1195, Y => n1272);
   U1404 : AOI22X1 port map( A => currentPlainKey_61_port, B => n207, C => n219
                           , D => n1451, Y => n1266);
   U1405 : NAND2X1 port map( A => n1450, B => RCV_DATA(5), Y => n1261);
   U1406 : NAND2X1 port map( A => n211, B => n1261, Y => n1262);
   U1407 : NAND2X1 port map( A => n1263, B => n1262, Y => n1265);
   U1408 : NAND2X1 port map( A => n1357, B => n1363, Y => n1264);
   U1409 : NAND3X1 port map( A => n1266, B => n1265, C => n1264, Y => n1271);
   U1410 : AND2X2 port map( A => n207, B => currentPlainKey_62_port, Y => n1267
                           );
   U1411 : AOI21X1 port map( A => n217, B => n1450, C => n1267, Y => n1362);
   U1412 : NOR2X1 port map( A => n1450, B => n1364, Y => n1268);
   U1413 : OAI21X1 port map( A => n190, B => n191, C => n1268, Y => n1359);
   U1414 : MUX2X1 port map( B => n1359, A => n1358, S => n1357, Y => n1360);
   U1415 : INVX2 port map( A => n1360, Y => n1361);
   U1416 : NAND2X1 port map( A => n1362, B => n1361, Y => n1270);
   U1417 : NAND2X1 port map( A => n207, B => currentPlainKey_63_port, Y => 
                           n1373);
   U1418 : NAND2X1 port map( A => n210, B => n1497, Y => n1369);
   U1419 : NOR2X1 port map( A => n1449, B => n1364, Y => n1366);
   U1420 : INVX2 port map( A => n155, Y => n1365);
   U1421 : OAI21X1 port map( A => n1367, B => n1366, C => n1365, Y => n1368);
   U1422 : NAND2X1 port map( A => n1369, B => n1368, Y => n1371);
   U1423 : MUX2X1 port map( B => n1371, A => n223, S => n1450, Y => n1372);
   U1424 : NAND2X1 port map( A => n1373, B => n1372, Y => n1269);
   U1425 : NAND2X1 port map( A => n1374, B => n1419, Y => n1385);
   U1426 : INVX2 port map( A => n1385, Y => n1375);
   U1427 : NAND3X1 port map( A => n1375, B => n242, C => n1431, Y => n1383);
   U1428 : INVX2 port map( A => n1383, Y => n1381);
   U1429 : NAND2X1 port map( A => n1381, B => keyCount_3_port, Y => n1384);
   U1430 : NAND2X1 port map( A => address_0_port, B => n1383, Y => n1376);
   U1431 : NAND2X1 port map( A => n1384, B => n1376, Y => n1333);
   U1432 : NAND2X1 port map( A => address_1_port, B => n1383, Y => n1377);
   U1433 : NAND2X1 port map( A => n1384, B => n1377, Y => n1334);
   U1434 : NAND2X1 port map( A => address_2_port, B => n1383, Y => n1378);
   U1435 : NAND2X1 port map( A => n1384, B => n1378, Y => n1335);
   U1436 : MUX2X1 port map( B => address_3_port, A => keyCount_0_port, S => 
                           n1381, Y => n1379);
   U1437 : NAND2X1 port map( A => n1384, B => n1379, Y => n1336);
   U1438 : MUX2X1 port map( B => address_4_port, A => keyCount_1_port, S => 
                           n1381, Y => n1380);
   U1439 : NAND2X1 port map( A => n1384, B => n1380, Y => n1337);
   U1440 : MUX2X1 port map( B => address_5_port, A => keyCount_2_port, S => 
                           n1381, Y => n1382);
   U1441 : NAND2X1 port map( A => n1384, B => n1382, Y => n1338);
   U1442 : OAI21X1 port map( A => n1503, B => n1381, C => n1384, Y => n1339);
   U1443 : OAI21X1 port map( A => n1495, B => n1381, C => n1384, Y => n1340);
   U1444 : OAI21X1 port map( A => n1386, B => n1385, C => parityError, Y => 
                           n1389);
   U1445 : OAI21X1 port map( A => n12, B => n13, C => n1387, Y => n1388);
   U1446 : NAND2X1 port map( A => n1389, B => n1388, Y => nextParityError);
   U1447 : NOR2X1 port map( A => keyCount_0_port, B => n1442, Y => n1390);
   U1448 : NOR2X1 port map( A => n1390, B => n1446, Y => n1393);
   U1449 : INVX2 port map( A => n1448, Y => n1391);
   U1450 : NAND2X1 port map( A => keyCount_0_port, B => n1391, Y => n1392);
   U1451 : MUX2X1 port map( B => n1393, A => n1392, S => n1494, Y => n1350);
   U1452 : NAND2X1 port map( A => n1399, B => CLR_RBUFF_port, Y => n1411);
   U1453 : INVX2 port map( A => n1411, Y => n1404);
   U1454 : NAND2X1 port map( A => N1799, B => n1404, Y => n1394);
   U1455 : OAI21X1 port map( A => n1493, B => n1395, C => n1394, Y => n1341);
   U1456 : NAND2X1 port map( A => N1798, B => n1404, Y => n1396);
   U1457 : OAI21X1 port map( A => n1492, B => n1397, C => n1396, Y => n1342);
   U1458 : NAND2X1 port map( A => N1797, B => n1404, Y => n1398);
   U1459 : OAI21X1 port map( A => n1491, B => n1399, C => n1398, Y => n1343);
   U1460 : NAND2X1 port map( A => N1796, B => n1404, Y => n1400);
   U1461 : OAI21X1 port map( A => n1490, B => n1401, C => n1400, Y => n1344);
   U1462 : NAND2X1 port map( A => N1795, B => n1404, Y => n1402);
   U1463 : OAI21X1 port map( A => n1489, B => n1403, C => n1402, Y => n1345);
   U1464 : NAND2X1 port map( A => N1794, B => n1404, Y => n1405);
   U1465 : OAI21X1 port map( A => n1488, B => n1406, C => n1405, Y => n1346);
   U1466 : INVX2 port map( A => N1793, Y => n1407);
   U1467 : OAI22X1 port map( A => n1487, B => n1408, C => n1411, D => n1407, Y 
                           => n1347);
   U1468 : INVX2 port map( A => N1792, Y => n1410);
   U1469 : OAI22X1 port map( A => n1486, B => n1408, C => n1411, D => n1410, Y 
                           => n1348);
   U1470 : AOI21X1 port map( A => N694, B => RBUF_FULL, C => n1178, Y => n1412)
                           ;
   U1471 : NAND2X1 port map( A => n1412, B => n83, Y => n1415);
   U1472 : NAND2X1 port map( A => n1413, B => n89, Y => n1414);
   U1473 : NAND2X1 port map( A => n1414, B => n1429, Y => n1436);
   U1474 : NAND2X1 port map( A => n1415, B => n1436, Y => n1426);
   U1475 : INVX2 port map( A => n1426, Y => n1418);
   U1476 : OAI21X1 port map( A => n1418, B => n89, C => n1416, Y => n1354);
   U1477 : OAI21X1 port map( A => OE, B => SBE, C => n83, Y => n1422);
   U1478 : OAI22X1 port map( A => RBUF_FULL, B => n1419, C => n131, D => n1436,
                           Y => n1420);
   U1479 : AOI21X1 port map( A => n1425, B => n1437, C => n1420, Y => n1421);
   U1480 : NAND3X1 port map( A => n1423, B => n1422, C => n1421, Y => n1352);
   U1481 : AOI21X1 port map( A => state_1_port, B => n1426, C => n1425, Y => 
                           n1427);
   U1482 : NAND2X1 port map( A => n127, B => n1427, Y => n1351);
   U1483 : INVX2 port map( A => RBUF_FULL, Y => n1428);
   U1484 : AOI21X1 port map( A => n1430, B => n1429, C => n1428, Y => n1435);
   U1485 : NAND2X1 port map( A => n1574, B => n1579, Y => n1433);
   U1486 : OAI21X1 port map( A => n1433, B => n1432, C => n93, Y => n1434);
   U1487 : NOR2X1 port map( A => n1435, B => n1434, Y => n1441);
   U1488 : INVX2 port map( A => n1160, Y => n1437);
   U1489 : OAI22X1 port map( A => n1442, B => n1437, C => n139, D => n1436, Y 
                           => n1438);
   U1490 : NOR2X1 port map( A => n1439, B => n1438, Y => n1440);
   U1491 : NAND2X1 port map( A => n1441, B => n1440, Y => n1353);
   U1492 : NOR2X1 port map( A => keyCount_2_port, B => n1442, Y => n1444);
   U1493 : OAI21X1 port map( A => n1444, B => n1443, C => keyCount_3_port, Y =>
                           n1445);
   U1494 : OAI21X1 port map( A => n1160, B => n1448, C => n1445, Y => n1355);
   U1495 : NAND2X1 port map( A => n1446, B => keyCount_0_port, Y => n1447);
   U1496 : OAI21X1 port map( A => keyCount_0_port, B => n1448, C => n1447, Y =>
                           n1356);
   U1497 : INVX2 port map( A => keyCount_3_port, Y => N694);
   U1498 : INVX2 port map( A => keyCount_0_port, Y => n1483);
   U1499 : INVX2 port map( A => keyCount_2_port, Y => n1484);
   U1500 : INVX2 port map( A => parityAccumulator_0_port, Y => n1486);
   U1501 : INVX2 port map( A => parityAccumulator_1_port, Y => n1487);
   U1502 : INVX2 port map( A => parityAccumulator_2_port, Y => n1488);
   U1503 : INVX2 port map( A => parityAccumulator_3_port, Y => n1489);
   U1504 : INVX2 port map( A => parityAccumulator_4_port, Y => n1490);
   U1505 : INVX2 port map( A => parityAccumulator_5_port, Y => n1491);
   U1506 : INVX2 port map( A => parityAccumulator_6_port, Y => n1492);
   U1507 : INVX2 port map( A => parityAccumulator_7_port, Y => n1493);
   U1508 : INVX2 port map( A => keyCount_1_port, Y => n1494);
   U1509 : INVX2 port map( A => address_7_port, Y => n1495);
   U1510 : INVX2 port map( A => n204, Y => n1496);
   U1511 : INVX2 port map( A => n157, Y => n1497);
   U1512 : INVX2 port map( A => n164, Y => n1498);
   U1513 : INVX2 port map( A => n167, Y => n1499);
   U1514 : INVX2 port map( A => n171, Y => n1500);
   U1515 : INVX2 port map( A => n176, Y => n1501);
   U1516 : INVX2 port map( A => address_6_port, Y => n1503);
   U1517 : INVX2 port map( A => n274, Y => n1504);
   U1518 : INVX2 port map( A => n254, Y => n1505);
   U1519 : INVX2 port map( A => n218, Y => n1506);
   U1520 : INVX2 port map( A => n179, Y => n1507);
   U1521 : INVX2 port map( A => address_5_port, Y => n1508);
   U1522 : INVX2 port map( A => address_4_port, Y => n1509);
   U1523 : INVX2 port map( A => currentPlainKey_63_port, Y => n1510);
   U1524 : INVX2 port map( A => currentPlainKey_62_port, Y => n1511);
   U1525 : INVX2 port map( A => currentPlainKey_61_port, Y => n1512);
   U1526 : INVX2 port map( A => currentPlainKey_60_port, Y => n1513);
   U1527 : INVX2 port map( A => currentPlainKey_59_port, Y => n1514);
   U1528 : INVX2 port map( A => currentPlainKey_58_port, Y => n1515);
   U1529 : INVX2 port map( A => currentPlainKey_57_port, Y => n1516);
   U1530 : INVX2 port map( A => currentPlainKey_56_port, Y => n1517);
   U1531 : INVX2 port map( A => currentPlainKey_55_port, Y => n1518);
   U1532 : INVX2 port map( A => currentPlainKey_54_port, Y => n1519);
   U1533 : INVX2 port map( A => currentPlainKey_53_port, Y => n1520);
   U1534 : INVX2 port map( A => currentPlainKey_52_port, Y => n1521);
   U1535 : INVX2 port map( A => currentPlainKey_51_port, Y => n1522);
   U1536 : INVX2 port map( A => currentPlainKey_50_port, Y => n1523);
   U1537 : INVX2 port map( A => currentPlainKey_49_port, Y => n1524);
   U1538 : INVX2 port map( A => currentPlainKey_48_port, Y => n1525);
   U1539 : INVX2 port map( A => currentPlainKey_47_port, Y => n1526);
   U1540 : INVX2 port map( A => currentPlainKey_46_port, Y => n1527);
   U1541 : INVX2 port map( A => currentPlainKey_45_port, Y => n1528);
   U1542 : INVX2 port map( A => currentPlainKey_44_port, Y => n1529);
   U1543 : INVX2 port map( A => currentPlainKey_43_port, Y => n1530);
   U1544 : INVX2 port map( A => currentPlainKey_42_port, Y => n1531);
   U1545 : INVX2 port map( A => currentPlainKey_41_port, Y => n1532);
   U1546 : INVX2 port map( A => currentPlainKey_40_port, Y => n1533);
   U1547 : INVX2 port map( A => currentPlainKey_39_port, Y => n1534);
   U1548 : INVX2 port map( A => currentPlainKey_38_port, Y => n1535);
   U1549 : INVX2 port map( A => currentPlainKey_37_port, Y => n1536);
   U1550 : INVX2 port map( A => currentPlainKey_36_port, Y => n1537);
   U1551 : INVX2 port map( A => currentPlainKey_35_port, Y => n1538);
   U1552 : INVX2 port map( A => currentPlainKey_34_port, Y => n1539);
   U1553 : INVX2 port map( A => currentPlainKey_33_port, Y => n1540);
   U1554 : INVX2 port map( A => currentPlainKey_32_port, Y => n1541);
   U1555 : INVX2 port map( A => currentPlainKey_31_port, Y => n1542);
   U1556 : INVX2 port map( A => currentPlainKey_30_port, Y => n1543);
   U1557 : INVX2 port map( A => currentPlainKey_29_port, Y => n1544);
   U1558 : INVX2 port map( A => currentPlainKey_28_port, Y => n1545);
   U1559 : INVX2 port map( A => currentPlainKey_27_port, Y => n1546);
   U1560 : INVX2 port map( A => currentPlainKey_26_port, Y => n1547);
   U1561 : INVX2 port map( A => currentPlainKey_25_port, Y => n1548);
   U1562 : INVX2 port map( A => currentPlainKey_24_port, Y => n1549);
   U1563 : INVX2 port map( A => currentPlainKey_23_port, Y => n1550);
   U1564 : INVX2 port map( A => currentPlainKey_22_port, Y => n1551);
   U1565 : INVX2 port map( A => currentPlainKey_21_port, Y => n1552);
   U1566 : INVX2 port map( A => currentPlainKey_20_port, Y => n1553);
   U1567 : INVX2 port map( A => currentPlainKey_19_port, Y => n1554);
   U1568 : INVX2 port map( A => currentPlainKey_18_port, Y => n1555);
   U1569 : INVX2 port map( A => currentPlainKey_17_port, Y => n1556);
   U1570 : INVX2 port map( A => currentPlainKey_16_port, Y => n1557);
   U1571 : INVX2 port map( A => currentPlainKey_15_port, Y => n1558);
   U1572 : INVX2 port map( A => currentPlainKey_14_port, Y => n1559);
   U1573 : INVX2 port map( A => currentPlainKey_13_port, Y => n1560);
   U1574 : INVX2 port map( A => currentPlainKey_12_port, Y => n1561);
   U1575 : INVX2 port map( A => currentPlainKey_11_port, Y => n1562);
   U1576 : INVX2 port map( A => currentPlainKey_10_port, Y => n1563);
   U1577 : INVX2 port map( A => currentPlainKey_9_port, Y => n1564);
   U1578 : INVX2 port map( A => currentPlainKey_8_port, Y => n1565);
   U1579 : INVX2 port map( A => currentPlainKey_7_port, Y => n1566);
   U1580 : INVX2 port map( A => currentPlainKey_6_port, Y => n1567);
   U1581 : INVX2 port map( A => currentPlainKey_5_port, Y => n1568);
   U1582 : INVX2 port map( A => currentPlainKey_4_port, Y => n1569);
   U1583 : INVX2 port map( A => currentPlainKey_0_port, Y => n1573);
   U1584 : INVX2 port map( A => SBE, Y => n1574);
   U1585 : INVX2 port map( A => OE, Y => n1579);

end SYN_keyb;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_sr_10bit_1 is

   port( CLK, RST, SHIFT_STROBE, SERIAL_IN : in std_logic;  LOAD_DATA : out 
         std_logic_vector (7 downto 0);  STOP_DATA : out std_logic_vector (1 
         downto 0));

end uart_sr_10bit_1;

architecture SYN_dataflow of uart_sr_10bit_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal LOAD_DATA_7_port, LOAD_DATA_6_port, LOAD_DATA_5_port, 
      LOAD_DATA_4_port, LOAD_DATA_3_port, LOAD_DATA_2_port, LOAD_DATA_1_port, 
      LOAD_DATA_0_port, STOP_DATA_1_port, STOP_DATA_0_port, n3, n12, n14, n16, 
      n18, n20, n22, n24, n26, n28, n30, n33, n1, n2, n4, n5, n6, n7, n8, n9, 
      n10, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, n32 : 
      std_logic;

begin
   LOAD_DATA <= ( LOAD_DATA_7_port, LOAD_DATA_6_port, LOAD_DATA_5_port, 
      LOAD_DATA_4_port, LOAD_DATA_3_port, LOAD_DATA_2_port, LOAD_DATA_1_port, 
      LOAD_DATA_0_port );
   STOP_DATA <= ( STOP_DATA_1_port, STOP_DATA_0_port );
   
   U2 : OAI21X1 port map( A => n32, B => n13, C => n3, Y => n14);
   U3 : NAND2X1 port map( A => LOAD_DATA_0_port, B => n13, Y => n3);
   U4 : OAI22X1 port map( A => n13, B => n31, C => SHIFT_STROBE, D => n32, Y =>
                           n16);
   U6 : OAI22X1 port map( A => n13, B => n29, C => SHIFT_STROBE, D => n31, Y =>
                           n18);
   U8 : OAI22X1 port map( A => n13, B => n27, C => SHIFT_STROBE, D => n29, Y =>
                           n20);
   U10 : OAI22X1 port map( A => n13, B => n25, C => SHIFT_STROBE, D => n27, Y 
                           => n22);
   U12 : OAI22X1 port map( A => n13, B => n23, C => SHIFT_STROBE, D => n25, Y 
                           => n24);
   U14 : OAI22X1 port map( A => n13, B => n21, C => SHIFT_STROBE, D => n23, Y 
                           => n26);
   U16 : OAI22X1 port map( A => n13, B => n19, C => SHIFT_STROBE, D => n21, Y 
                           => n28);
   U18 : OAI22X1 port map( A => n13, B => n17, C => SHIFT_STROBE, D => n19, Y 
                           => n30);
   U22 : OAI21X1 port map( A => SHIFT_STROBE, B => n17, C => n12, Y => n33);
   U23 : NAND2X1 port map( A => SERIAL_IN, B => SHIFT_STROBE, Y => n12);
   present_val_reg_9_inst : DFFSR port map( D => n33, CLK => CLK, R => n15, S 
                           => n11, Q => STOP_DATA_1_port);
   present_val_reg_8_inst : DFFSR port map( D => n30, CLK => CLK, R => n15, S 
                           => n10, Q => STOP_DATA_0_port);
   present_val_reg_7_inst : DFFSR port map( D => n28, CLK => CLK, R => n15, S 
                           => n9, Q => LOAD_DATA_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n26, CLK => CLK, R => n15, S 
                           => n8, Q => LOAD_DATA_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n24, CLK => CLK, R => n15, S 
                           => n7, Q => LOAD_DATA_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n22, CLK => CLK, R => n15, S 
                           => n6, Q => LOAD_DATA_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n20, CLK => CLK, R => n15, S 
                           => n5, Q => LOAD_DATA_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n18, CLK => CLK, R => n15, S 
                           => n4, Q => LOAD_DATA_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n16, CLK => CLK, R => n15, S 
                           => n2, Q => LOAD_DATA_1_port);
   present_val_reg_0_inst : DFFSR port map( D => n14, CLK => CLK, R => n15, S 
                           => n1, Q => LOAD_DATA_0_port);
   n1 <= '1';
   n2 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   U24 : INVX2 port map( A => RST, Y => n15);
   U25 : INVX2 port map( A => SHIFT_STROBE, Y => n13);
   U26 : INVX2 port map( A => STOP_DATA_1_port, Y => n17);
   U27 : INVX2 port map( A => STOP_DATA_0_port, Y => n19);
   U28 : INVX2 port map( A => LOAD_DATA_7_port, Y => n21);
   U29 : INVX2 port map( A => LOAD_DATA_6_port, Y => n23);
   U30 : INVX2 port map( A => LOAD_DATA_5_port, Y => n25);
   U31 : INVX2 port map( A => LOAD_DATA_4_port, Y => n27);
   U32 : INVX2 port map( A => LOAD_DATA_3_port, Y => n29);
   U33 : INVX2 port map( A => LOAD_DATA_2_port, Y => n31);
   U34 : INVX2 port map( A => LOAD_DATA_1_port, Y => n32);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_sb_check_1 is

   port( RST, CLK, SBC_CLR, SBC_EN : in std_logic;  STOP_DATA : in 
         std_logic_vector (1 downto 0);  SB_DETECT, SBE : out std_logic);

end uart_sb_check_1;

architecture SYN_behavioral of uart_sb_check_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal SBE_prime, sb_detect_flag, n7, n8, n9, n1, n2, n3, n4, n5, n6 : 
      std_logic;

begin
   
   U6 : OR2X2 port map( A => SBC_CLR, B => STOP_DATA(0), Y => n7);
   U10 : NOR2X1 port map( A => n7, B => n8, Y => sb_detect_flag);
   U11 : NAND2X1 port map( A => STOP_DATA(1), B => SBC_EN, Y => n8);
   U12 : NOR2X1 port map( A => n6, B => n9, Y => SBE_prime);
   U13 : OAI21X1 port map( A => STOP_DATA(0), B => n4, C => n5, Y => n9);
   SBE_reg : DFFSR port map( D => SBE_prime, CLK => CLK, R => n3, S => n2, Q =>
                           SBE);
   SB_DETECT_reg : DFFSR port map( D => sb_detect_flag, CLK => CLK, R => n3, S 
                           => n1, Q => SB_DETECT);
   n1 <= '1';
   n2 <= '1';
   U5 : INVX2 port map( A => RST, Y => n3);
   U7 : INVX2 port map( A => STOP_DATA(1), Y => n4);
   U8 : INVX2 port map( A => SBC_CLR, Y => n5);
   U9 : INVX2 port map( A => SBC_EN, Y => n6);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_buf_full_1 is

   port( CLK, RST, CLR_RBUF, SET_RBUF_FULL : in std_logic;  RBUF_FULL : out 
         std_logic);

end uart_rcv_buf_full_1;

architecture SYN_Behavioral of uart_rcv_buf_full_1 is

   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal RBUF_FULL_port, n1, n3, n2 : std_logic;

begin
   RBUF_FULL <= RBUF_FULL_port;
   
   U3 : NOR2X1 port map( A => RST, B => CLR_RBUF, Y => n1);
   U4 : OR2X2 port map( A => RBUF_FULL_port, B => SET_RBUF_FULL, Y => n3);
   Q_int_reg : DFFSR port map( D => n3, CLK => CLK, R => n1, S => n2, Q => 
                           RBUF_FULL_port);
   n2 <= '1';

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_buf_1 is

   port( CLK, RST, LOAD_RBUF : in std_logic;  LOAD_DATA : in std_logic_vector 
         (7 downto 0);  RCV_DATA : out std_logic_vector (7 downto 0));

end uart_rcv_buf_1;

architecture SYN_Behavioral of uart_rcv_buf_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, n1, 
      n3, n4, n5, n6, n7, n8, n9, n2, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27 : std_logic;

begin
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   U3 : AOI22X1 port map( A => n17, B => LOAD_DATA(0), C => RCV_DATA_0_port, D 
                           => n27, Y => n1);
   U5 : AOI22X1 port map( A => LOAD_DATA(1), B => n17, C => RCV_DATA_1_port, D 
                           => n27, Y => n3);
   U7 : AOI22X1 port map( A => LOAD_DATA(2), B => n17, C => RCV_DATA_2_port, D 
                           => n27, Y => n4);
   U9 : AOI22X1 port map( A => LOAD_DATA(3), B => n17, C => RCV_DATA_3_port, D 
                           => n27, Y => n5);
   U11 : AOI22X1 port map( A => LOAD_DATA(4), B => n17, C => RCV_DATA_4_port, D
                           => n27, Y => n6);
   U13 : AOI22X1 port map( A => LOAD_DATA(5), B => n17, C => RCV_DATA_5_port, D
                           => n27, Y => n7);
   U15 : AOI22X1 port map( A => LOAD_DATA(6), B => n17, C => RCV_DATA_6_port, D
                           => n27, Y => n8);
   U18 : AOI22X1 port map( A => LOAD_DATA(7), B => n17, C => RCV_DATA_7_port, D
                           => n27, Y => n9);
   Q_int_reg_0_inst : DFFSR port map( D => n26, CLK => CLK, R => n18, S => n16,
                           Q => RCV_DATA_0_port);
   Q_int_reg_7_inst : DFFSR port map( D => n19, CLK => CLK, R => n18, S => n15,
                           Q => RCV_DATA_7_port);
   Q_int_reg_6_inst : DFFSR port map( D => n20, CLK => CLK, R => n18, S => n14,
                           Q => RCV_DATA_6_port);
   Q_int_reg_5_inst : DFFSR port map( D => n21, CLK => CLK, R => n18, S => n13,
                           Q => RCV_DATA_5_port);
   Q_int_reg_4_inst : DFFSR port map( D => n22, CLK => CLK, R => n18, S => n12,
                           Q => RCV_DATA_4_port);
   Q_int_reg_2_inst : DFFSR port map( D => n24, CLK => CLK, R => n18, S => n11,
                           Q => RCV_DATA_2_port);
   Q_int_reg_3_inst : DFFSR port map( D => n23, CLK => CLK, R => n18, S => n10,
                           Q => RCV_DATA_3_port);
   Q_int_reg_1_inst : DFFSR port map( D => n25, CLK => CLK, R => n18, S => n2, 
                           Q => RCV_DATA_1_port);
   n2 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   U17 : INVX2 port map( A => RST, Y => n18);
   U19 : BUFX2 port map( A => LOAD_RBUF, Y => n17);
   U20 : INVX2 port map( A => n9, Y => n19);
   U21 : INVX2 port map( A => n8, Y => n20);
   U22 : INVX2 port map( A => n7, Y => n21);
   U23 : INVX2 port map( A => n6, Y => n22);
   U24 : INVX2 port map( A => n5, Y => n23);
   U25 : INVX2 port map( A => n4, Y => n24);
   U26 : INVX2 port map( A => n3, Y => n25);
   U27 : INVX2 port map( A => n1, Y => n26);
   U28 : INVX2 port map( A => n17, Y => n27);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcu_1 is

   port( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT : in std_logic;  RBUF_LOAD
         , TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR : out 
         std_logic);

end uart_rcu_1;

architecture SYN_rcub of uart_rcu_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal RBUF_LOAD_port, TIMER_TRIG_port, CHK_ERROR_port, SET_RBUF_FULL_port, 
      SBC_EN_port, SBC_CLR_port, state_2_port, state_1_port, state_0_port, 
      timerRunning, count_7_port, count_6_port, count_5_port, count_4_port, 
      count_3_port, count_2_port, count_1_port, count_0_port, nextCount_7_port,
      nextCount_6_port, nextCount_5_port, nextCount_4_port, nextCount_3_port, 
      nextCount_2_port, nextCount_1_port, nextCount_0_port, nextState_1_port, 
      nextState_0_port, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, 
      N35, N36, N37, N38, N99, n21, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, add_46_carry_3_port, 
      add_46_carry_4_port, add_46_carry_5_port, add_46_carry_6_port, 
      add_46_carry_7_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n22, n23, n24_port, n25_port, 
      n26_port, n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, 
      n33_port, n34_port, n35_port, n36_port, n37_port, n38_port, n39, n40, n41
      , n42, n43, n44, n45, n46, n47 : std_logic;

begin
   RBUF_LOAD <= RBUF_LOAD_port;
   TIMER_TRIG <= TIMER_TRIG_port;
   CHK_ERROR <= CHK_ERROR_port;
   SET_RBUF_FULL <= SET_RBUF_FULL_port;
   SBC_EN <= SBC_EN_port;
   SBC_CLR <= SBC_CLR_port;
   
   nextCount_reg_0_inst : DFFSR port map( D => N31, CLK => CLK, R => n21, S => 
                           n27_port, Q => nextCount_0_port);
   n21 <= '1';
   U33 : AND2X2 port map( A => N30, B => timerRunning, Y => N38);
   U34 : AND2X2 port map( A => N29, B => timerRunning, Y => N37);
   U35 : AND2X2 port map( A => N28, B => timerRunning, Y => N36);
   U36 : AND2X2 port map( A => N27, B => timerRunning, Y => N35);
   U37 : AND2X2 port map( A => N26, B => timerRunning, Y => N34);
   U38 : AND2X2 port map( A => N25, B => timerRunning, Y => N33);
   U39 : AND2X2 port map( A => N24, B => timerRunning, Y => N32);
   U54 : OAI21X1 port map( A => n49, B => n43, C => n50, Y => n48);
   U55 : OAI21X1 port map( A => n44, B => n42, C => n43, Y => n50);
   U56 : NAND2X1 port map( A => n51, B => n52, Y => n74);
   U57 : OAI21X1 port map( A => n53, B => n54, C => timerRunning, Y => n52);
   U58 : NAND2X1 port map( A => n55, B => n56, Y => n54);
   U59 : NAND2X1 port map( A => n57, B => n56, Y => n75);
   U60 : NAND3X1 port map( A => n35_port, B => n51, C => CHK_ERROR_port, Y => 
                           n57);
   U61 : OAI21X1 port map( A => n58, B => n47, C => n59, Y => n76);
   U62 : NAND2X1 port map( A => n56, B => n60, Y => n58);
   U63 : NAND2X1 port map( A => n61, B => n38_port, Y => n56);
   U64 : NAND3X1 port map( A => n62, B => n63, C => n64, Y => n77);
   U65 : NAND3X1 port map( A => n34_port, B => n51, C => SET_RBUF_FULL_port, Y 
                           => n64);
   U66 : NAND2X1 port map( A => n60, B => n63, Y => n53);
   U67 : NAND3X1 port map( A => nextState_0_port, B => nextState_1_port, C => 
                           n61, Y => n63);
   U68 : NAND3X1 port map( A => n36_port, B => n38_port, C => n61, Y => n62);
   U69 : OAI21X1 port map( A => n65, B => n45, C => n51, Y => n78);
   U70 : OAI21X1 port map( A => n65, B => n46, C => n51, Y => n79);
   U71 : NAND2X1 port map( A => n60, B => n59, Y => n65);
   U72 : NAND3X1 port map( A => nextState_1_port, B => n36_port, C => n39, Y =>
                           n59);
   U73 : NAND2X1 port map( A => n66, B => n55, Y => n80);
   U74 : NAND3X1 port map( A => nextState_1_port, B => n36_port, C => n61, Y =>
                           n55);
   U75 : NAND3X1 port map( A => n60, B => n51, C => RBUF_LOAD_port, Y => n66);
   U76 : NAND3X1 port map( A => nextState_0_port, B => n38_port, C => n39, Y =>
                           n51);
   U77 : NAND3X1 port map( A => n36_port, B => n38_port, C => n39, Y => n60);
   U78 : OAI21X1 port map( A => n40, B => n43, C => n67, Y => n61);
   U79 : NAND3X1 port map( A => state_0_port, B => n43, C => state_1_port, Y =>
                           n67);
   U80 : NAND2X1 port map( A => n68, B => n69, Y => n49);
   U81 : OAI21X1 port map( A => n70, B => n69, C => n68, Y => nextState_1_port)
                           ;
   U82 : NOR2X1 port map( A => N99, B => state_2_port, Y => n70);
   U83 : OAI21X1 port map( A => state_2_port, B => n71, C => n68, Y => 
                           nextState_0_port);
   U84 : NAND2X1 port map( A => state_1_port, B => n44, Y => n68);
   U85 : AOI21X1 port map( A => START_BIT, B => n44, C => n72, Y => n71);
   U86 : OAI21X1 port map( A => N99, B => n69, C => n73, Y => n72);
   U87 : NAND2X1 port map( A => SB_DETECT, B => state_1_port, Y => n73);
   U88 : NAND2X1 port map( A => state_0_port, B => n42, Y => n69);
   U89 : NAND2X1 port map( A => n37_port, B => timerRunning, Y => N31);
   count_reg_7_inst : DFFSR port map( D => nextCount_7_port, CLK => CLK, R => 
                           n27_port, S => n26_port, Q => count_7_port);
   count_reg_6_inst : DFFSR port map( D => nextCount_6_port, CLK => CLK, R => 
                           n27_port, S => n25_port, Q => count_6_port);
   count_reg_5_inst : DFFSR port map( D => nextCount_5_port, CLK => CLK, R => 
                           n27_port, S => n24_port, Q => count_5_port);
   count_reg_4_inst : DFFSR port map( D => nextCount_4_port, CLK => CLK, R => 
                           n27_port, S => n23, Q => count_4_port);
   count_reg_3_inst : DFFSR port map( D => nextCount_3_port, CLK => CLK, R => 
                           n27_port, S => n22, Q => count_3_port);
   count_reg_2_inst : DFFSR port map( D => nextCount_2_port, CLK => CLK, R => 
                           n27_port, S => n20, Q => count_2_port);
   count_reg_1_inst : DFFSR port map( D => nextCount_1_port, CLK => CLK, R => 
                           n27_port, S => n19, Q => count_1_port);
   count_reg_0_inst : DFFSR port map( D => nextCount_0_port, CLK => CLK, R => 
                           n27_port, S => n18, Q => count_0_port);
   nextCount_reg_2_inst : DFFSR port map( D => N33, CLK => CLK, R => n27_port, 
                           S => n17, Q => nextCount_2_port);
   nextCount_reg_1_inst : DFFSR port map( D => N32, CLK => CLK, R => n27_port, 
                           S => n16, Q => nextCount_1_port);
   state_reg_2_inst : DFFSR port map( D => n41, CLK => CLK, R => n27_port, S =>
                           n15, Q => state_2_port);
   nextCount_reg_3_inst : DFFSR port map( D => N34, CLK => CLK, R => n27_port, 
                           S => n14, Q => nextCount_3_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n27_port, S => n13, Q => state_1_port);
   nextCount_reg_4_inst : DFFSR port map( D => N35, CLK => CLK, R => n27_port, 
                           S => n12, Q => nextCount_4_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n27_port, S => n11, Q => state_0_port);
   nextCount_reg_5_inst : DFFSR port map( D => N36, CLK => CLK, R => n27_port, 
                           S => n10, Q => nextCount_5_port);
   nextCount_reg_6_inst : DFFSR port map( D => N37, CLK => CLK, R => n27_port, 
                           S => n9, Q => nextCount_6_port);
   RBUF_LOAD_reg : DFFSR port map( D => n80, CLK => CLK, R => n27_port, S => n8
                           , Q => RBUF_LOAD_port);
   timerRunning_reg : DFFSR port map( D => n74, CLK => CLK, R => n27_port, S =>
                           n7, Q => timerRunning);
   TIMER_TRIG_reg : DFFSR port map( D => n79, CLK => CLK, R => n27_port, S => 
                           n6, Q => TIMER_TRIG_port);
   SBC_CLR_reg : DFFSR port map( D => n78, CLK => CLK, R => n27_port, S => n5, 
                           Q => SBC_CLR_port);
   SBC_EN_reg : DFFSR port map( D => n76, CLK => CLK, R => n27_port, S => n4, Q
                           => SBC_EN_port);
   nextCount_reg_7_inst : DFFSR port map( D => N38, CLK => CLK, R => n27_port, 
                           S => n3, Q => nextCount_7_port);
   SET_RBUF_FULL_reg : DFFSR port map( D => n77, CLK => CLK, R => n27_port, S 
                           => n2, Q => SET_RBUF_FULL_port);
   CHK_ERROR_reg : DFFSR port map( D => n75, CLK => CLK, R => n27_port, S => n1
                           , Q => CHK_ERROR_port);
   U3 : INVX4 port map( A => RST, Y => n27_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   n18 <= '1';
   n19 <= '1';
   n20 <= '1';
   n22 <= '1';
   n23 <= '1';
   n24_port <= '1';
   n25_port <= '1';
   n26_port <= '1';
   U30 : XOR2X1 port map( A => count_7_port, B => add_46_carry_7_port, Y => N30
                           );
   U31 : AND2X1 port map( A => count_6_port, B => add_46_carry_6_port, Y => 
                           add_46_carry_7_port);
   U32 : XOR2X1 port map( A => add_46_carry_6_port, B => count_6_port, Y => N29
                           );
   U40 : AND2X1 port map( A => count_5_port, B => add_46_carry_5_port, Y => 
                           add_46_carry_6_port);
   U41 : XOR2X1 port map( A => add_46_carry_5_port, B => count_5_port, Y => N28
                           );
   U42 : AND2X1 port map( A => count_4_port, B => add_46_carry_4_port, Y => 
                           add_46_carry_5_port);
   U43 : XOR2X1 port map( A => add_46_carry_4_port, B => count_4_port, Y => N27
                           );
   U44 : AND2X1 port map( A => count_3_port, B => add_46_carry_3_port, Y => 
                           add_46_carry_4_port);
   U45 : XOR2X1 port map( A => add_46_carry_3_port, B => count_3_port, Y => N26
                           );
   U46 : AND2X1 port map( A => count_2_port, B => count_1_port, Y => 
                           add_46_carry_3_port);
   U47 : XOR2X1 port map( A => count_1_port, B => count_2_port, Y => N25);
   U48 : INVX2 port map( A => count_1_port, Y => N24);
   U49 : OAI21X1 port map( A => count_0_port, B => count_1_port, C => 
                           count_2_port, Y => n28_port);
   U50 : NOR2X1 port map( A => n33_port, B => n28_port, Y => n29_port);
   U51 : OAI21X1 port map( A => n29_port, B => count_4_port, C => count_6_port,
                           Y => n30_port);
   U52 : OAI21X1 port map( A => n32_port, B => n30_port, C => n31_port, Y => 
                           N99);
   U53 : INVX2 port map( A => count_7_port, Y => n31_port);
   U90 : INVX2 port map( A => count_5_port, Y => n32_port);
   U91 : INVX2 port map( A => count_3_port, Y => n33_port);
   U92 : INVX2 port map( A => n53, Y => n34_port);
   U93 : INVX2 port map( A => n58, Y => n35_port);
   U94 : INVX2 port map( A => nextState_0_port, Y => n36_port);
   U95 : INVX2 port map( A => count_0_port, Y => n37_port);
   U96 : INVX2 port map( A => nextState_1_port, Y => n38_port);
   U97 : INVX2 port map( A => n61, Y => n39);
   U98 : INVX2 port map( A => n49, Y => n40);
   U99 : INVX2 port map( A => n48, Y => n41);
   U100 : INVX2 port map( A => state_1_port, Y => n42);
   U101 : INVX2 port map( A => state_2_port, Y => n43);
   U102 : INVX2 port map( A => state_0_port, Y => n44);
   U103 : INVX2 port map( A => SBC_CLR_port, Y => n45);
   U104 : INVX2 port map( A => TIMER_TRIG_port, Y => n46);
   U105 : INVX2 port map( A => SBC_EN_port, Y => n47);

end SYN_rcub;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_error_1 is

   port( RST, CLK, RBUF_FULL, CHK_ERROR : in std_logic;  OE : out std_logic);

end uart_error_1;

architecture SYN_behavioral of uart_error_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal OE_prime, n1, n2 : std_logic;

begin
   
   U5 : AND2X2 port map( A => RBUF_FULL, B => CHK_ERROR, Y => OE_prime);
   OE_reg : DFFSR port map( D => OE_prime, CLK => CLK, R => n2, S => n1, Q => 
                           OE);
   n1 <= '1';
   U4 : INVX2 port map( A => RST, Y => n2);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_edge_detector_1 is

   port( CLK, RST, SERIAL_IN : in std_logic;  START_BIT : out std_logic);

end uart_edge_detector_1;

architecture SYN_Behavioral of uart_edge_detector_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal Q_int, Q_int2, n3, n1, n2, n4 : std_logic;

begin
   
   Q_int_reg : DFFSR port map( D => SERIAL_IN, CLK => CLK, R => n2, S => n3, Q 
                           => Q_int);
   n3 <= '1';
   U7 : NOR2X1 port map( A => Q_int, B => n4, Y => START_BIT);
   Q_int2_reg : DFFSR port map( D => Q_int, CLK => CLK, R => n2, S => n1, Q => 
                           Q_int2);
   n1 <= '1';
   U4 : INVX2 port map( A => RST, Y => n2);
   U6 : INVX2 port map( A => Q_int2, Y => n4);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_timer_1 is

   port( CLK, RST, SENDING : in std_logic;  SHIFT_ENABLE_R, SHIFT_ENABLE_E : 
         out std_logic);

end tx_timer_1;

architecture SYN_moore of tx_timer_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_3_port, count_2_port, count_1_port, count_0_port, state, 
      nextcount_3_port, nextcount_2_port, nextcount_1_port, nextcount_0_port, 
      nxt_SHIFT_ENABLE_E, n12, n13, n14, n15, n16, n17, n18, n19, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   SHIFT_ENABLE_R <= nxt_SHIFT_ENABLE_E;
   
   U14 : NOR2X1 port map( A => n12, B => n13, Y => nextcount_3_port);
   U15 : XNOR2X1 port map( A => count_3_port, B => n14, Y => n12);
   U16 : NOR2X1 port map( A => n15, B => n9, Y => n14);
   U17 : AOI21X1 port map( A => n16, B => state, C => n11, Y => 
                           nextcount_2_port);
   U18 : XNOR2X1 port map( A => n15, B => n9, Y => n16);
   U19 : NAND2X1 port map( A => count_1_port, B => count_0_port, Y => n15);
   U20 : NOR2X1 port map( A => n17, B => n13, Y => nextcount_1_port);
   U21 : NAND3X1 port map( A => SENDING, B => n18, C => state, Y => n13);
   U22 : XNOR2X1 port map( A => count_0_port, B => count_1_port, Y => n17);
   U23 : OAI21X1 port map( A => count_0_port, B => n11, C => state, Y => 
                           nextcount_0_port);
   U24 : NOR2X1 port map( A => n18, B => n19, Y => nxt_SHIFT_ENABLE_E);
   U25 : NAND3X1 port map( A => count_3_port, B => SENDING, C => state, Y => 
                           n19);
   U26 : NAND3X1 port map( A => n10, B => n9, C => n8, Y => n18);
   state_reg : DFFSR port map( D => SENDING, CLK => CLK, R => n7, S => n6, Q =>
                           state);
   count_reg_2_inst : DFFSR port map( D => nextcount_2_port, CLK => CLK, R => 
                           n7, S => n5, Q => count_2_port);
   count_reg_0_inst : DFFSR port map( D => nextcount_0_port, CLK => CLK, R => 
                           n7, S => n4, Q => count_0_port);
   count_reg_3_inst : DFFSR port map( D => nextcount_3_port, CLK => CLK, R => 
                           n7, S => n3, Q => count_3_port);
   count_reg_1_inst : DFFSR port map( D => nextcount_1_port, CLK => CLK, R => 
                           n7, S => n2, Q => count_1_port);
   SHIFT_ENABLE_E_reg : DFFSR port map( D => nxt_SHIFT_ENABLE_E, CLK => CLK, R 
                           => n7, S => n1, Q => SHIFT_ENABLE_E);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   U9 : INVX2 port map( A => RST, Y => n7);
   U10 : INVX2 port map( A => count_0_port, Y => n8);
   U11 : INVX2 port map( A => count_2_port, Y => n9);
   U12 : INVX2 port map( A => count_1_port, Y => n10);
   U13 : INVX2 port map( A => SENDING, Y => n11);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_tcu_1 is

   port( clk, rst, p_ready, t_bitstuff : in std_logic;  PRGA_OUT : in 
         std_logic_vector (7 downto 0);  prga_opcode : in std_logic_vector (1 
         downto 0);  t_crc : in std_logic_vector (15 downto 0);  sending, EOP, 
         next_byte : out std_logic;  send_data : out std_logic_vector (7 downto
         0);  t_strobe : out std_logic);

end tx_tcu_1;

architecture SYN_behavioral of tx_tcu_1 is

   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component tx_tcu_1_DW01_inc_0
      port( A : in std_logic_vector (6 downto 0);  SUM : out std_logic_vector 
            (6 downto 0));
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal send_data_7_port, send_data_6_port, send_data_5_port, 
      send_data_4_port, send_data_3_port, send_data_2_port, send_data_1_port, 
      send_data_0_port, state_2_port, state_1_port, state_0_port, count_5_port,
      count_4_port, count_3_port, count_2_port, count_1_port, count_0_port, 
      nextstate_2_port, nextstate_1_port, nextstate_0_port, flop_data_7_port, 
      flop_data_6_port, flop_data_5_port, flop_data_4_port, flop_data_3_port, 
      flop_data_2_port, flop_data_1_port, flop_data_0_port, 
      current_send_data_7_port, current_send_data_6_port, 
      current_send_data_5_port, current_send_data_4_port, 
      current_send_data_3_port, current_send_data_2_port, 
      current_send_data_1_port, current_send_data_0_port, N59, N60, N61, N62, 
      N63, N64, N65, N84, N85, N86, N87, N88, N89, N90, N188, n158, n159, n160,
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n194, n195, n196, n197, n198, n199, n200, r81_carry_1_port, 
      r81_carry_2_port, r81_carry_3_port, r81_carry_4_port, r81_carry_5_port, 
      r81_carry_6_port, r81_B_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59_port, n60_port, n61_port, n62_port, n63_port, 
      n64_port, n65_port, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83, n84_port, n85_port, n86_port, 
      n87_port, n88_port, n89_port, n90_port, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n174, n175 : std_logic;

begin
   send_data <= ( send_data_7_port, send_data_6_port, send_data_5_port, 
      send_data_4_port, send_data_3_port, send_data_2_port, send_data_1_port, 
      send_data_0_port );
   
   flop_data_reg_7_inst : DFFPOSX1 port map( D => n152, CLK => clk, Q => 
                           flop_data_7_port);
   current_send_data_reg_7_inst : DFFPOSX1 port map( D => n173, CLK => clk, Q 
                           => current_send_data_7_port);
   flop_data_reg_6_inst : DFFPOSX1 port map( D => n153, CLK => clk, Q => 
                           flop_data_6_port);
   current_send_data_reg_6_inst : DFFPOSX1 port map( D => n172, CLK => clk, Q 
                           => current_send_data_6_port);
   flop_data_reg_5_inst : DFFPOSX1 port map( D => n154, CLK => clk, Q => 
                           flop_data_5_port);
   current_send_data_reg_5_inst : DFFPOSX1 port map( D => n171, CLK => clk, Q 
                           => current_send_data_5_port);
   flop_data_reg_4_inst : DFFPOSX1 port map( D => n155, CLK => clk, Q => 
                           flop_data_4_port);
   current_send_data_reg_4_inst : DFFPOSX1 port map( D => n170, CLK => clk, Q 
                           => current_send_data_4_port);
   flop_data_reg_3_inst : DFFPOSX1 port map( D => n156, CLK => clk, Q => 
                           flop_data_3_port);
   current_send_data_reg_3_inst : DFFPOSX1 port map( D => n169, CLK => clk, Q 
                           => current_send_data_3_port);
   flop_data_reg_2_inst : DFFPOSX1 port map( D => n157, CLK => clk, Q => 
                           flop_data_2_port);
   current_send_data_reg_2_inst : DFFPOSX1 port map( D => n168, CLK => clk, Q 
                           => current_send_data_2_port);
   flop_data_reg_1_inst : DFFPOSX1 port map( D => n174, CLK => clk, Q => 
                           flop_data_1_port);
   current_send_data_reg_1_inst : DFFPOSX1 port map( D => n167, CLK => clk, Q 
                           => current_send_data_1_port);
   flop_data_reg_0_inst : DFFPOSX1 port map( D => n175, CLK => clk, Q => 
                           flop_data_0_port);
   current_send_data_reg_0_inst : DFFPOSX1 port map( D => n166, CLK => clk, Q 
                           => current_send_data_0_port);
   send_data_reg_7_inst : DFFPOSX1 port map( D => n165, CLK => clk, Q => 
                           send_data_7_port);
   send_data_reg_6_inst : DFFPOSX1 port map( D => n164, CLK => clk, Q => 
                           send_data_6_port);
   send_data_reg_5_inst : DFFPOSX1 port map( D => n163, CLK => clk, Q => 
                           send_data_5_port);
   send_data_reg_4_inst : DFFPOSX1 port map( D => n162, CLK => clk, Q => 
                           send_data_4_port);
   send_data_reg_3_inst : DFFPOSX1 port map( D => n161, CLK => clk, Q => 
                           send_data_3_port);
   send_data_reg_2_inst : DFFPOSX1 port map( D => n160, CLK => clk, Q => 
                           send_data_2_port);
   send_data_reg_1_inst : DFFPOSX1 port map( D => n159, CLK => clk, Q => 
                           send_data_1_port);
   send_data_reg_0_inst : DFFPOSX1 port map( D => n158, CLK => clk, Q => 
                           send_data_0_port);
   r80 : tx_tcu_1_DW01_inc_0 port map( A(6) => N188, A(5) => count_5_port, A(4)
                           => count_4_port, A(3) => count_3_port, A(2) => 
                           count_2_port, A(1) => count_1_port, A(0) => 
                           count_0_port, SUM(6) => N65, SUM(5) => N64, SUM(4) 
                           => N63, SUM(3) => N62, SUM(2) => N61, SUM(1) => N60,
                           SUM(0) => N59);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n15, S => n10, Q => state_2_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n15, S => n9, Q => state_1_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n15, S => n8, Q => state_0_port);
   count_reg_3_inst : DFFSR port map( D => n196, CLK => clk, R => n15, S => n7,
                           Q => count_3_port);
   count_reg_2_inst : DFFSR port map( D => n195, CLK => clk, R => n15, S => n6,
                           Q => count_2_port);
   count_reg_1_inst : DFFSR port map( D => n194, CLK => clk, R => n15, S => n5,
                           Q => count_1_port);
   count_reg_0_inst : DFFSR port map( D => n200, CLK => clk, R => n15, S => n4,
                           Q => count_0_port);
   count_reg_4_inst : DFFSR port map( D => n197, CLK => clk, R => n15, S => n3,
                           Q => count_4_port);
   count_reg_5_inst : DFFSR port map( D => n198, CLK => clk, R => n15, S => n2,
                           Q => count_5_port);
   count_reg_6_inst : DFFSR port map( D => n199, CLK => clk, R => n15, S => n1,
                           Q => N188);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   U13 : INVX2 port map( A => n12, Y => n15);
   U14 : BUFX2 port map( A => rst, Y => n13);
   U15 : BUFX2 port map( A => rst, Y => n12);
   U16 : BUFX2 port map( A => rst, Y => n14);
   U17 : INVX2 port map( A => N188, Y => n11);
   U18 : XOR2X1 port map( A => N188, B => r81_carry_6_port, Y => N90);
   U19 : AND2X1 port map( A => count_5_port, B => r81_carry_5_port, Y => 
                           r81_carry_6_port);
   U20 : XOR2X1 port map( A => r81_carry_5_port, B => count_5_port, Y => N89);
   U21 : AND2X1 port map( A => count_4_port, B => r81_carry_4_port, Y => 
                           r81_carry_5_port);
   U22 : XOR2X1 port map( A => r81_carry_4_port, B => count_4_port, Y => N88);
   U23 : AND2X1 port map( A => count_3_port, B => r81_carry_3_port, Y => 
                           r81_carry_4_port);
   U24 : XOR2X1 port map( A => r81_carry_3_port, B => count_3_port, Y => N87);
   U25 : AND2X1 port map( A => count_2_port, B => r81_carry_2_port, Y => 
                           r81_carry_3_port);
   U26 : XOR2X1 port map( A => r81_carry_2_port, B => count_2_port, Y => N86);
   U27 : AND2X1 port map( A => count_1_port, B => r81_carry_1_port, Y => 
                           r81_carry_2_port);
   U28 : XOR2X1 port map( A => r81_carry_1_port, B => count_1_port, Y => N85);
   U29 : AND2X1 port map( A => count_0_port, B => r81_B_0_port, Y => 
                           r81_carry_1_port);
   U30 : XOR2X1 port map( A => r81_B_0_port, B => count_0_port, Y => N84);
   U31 : NOR2X1 port map( A => n16, B => n17, Y => t_strobe);
   U32 : NAND2X1 port map( A => n18, B => n19, Y => n17);
   U33 : NAND2X1 port map( A => n11, B => n20, Y => n16);
   U34 : OR2X1 port map( A => n21, B => n22, Y => sending);
   U35 : OAI21X1 port map( A => N188, B => n23, C => n24, Y => n22);
   U36 : NAND3X1 port map( A => n25, B => n26, C => n27, Y => n21);
   U37 : NAND3X1 port map( A => n28, B => n27, C => n29, Y => nextstate_2_port)
                           ;
   U38 : AOI22X1 port map( A => n30, B => p_ready, C => n31, D => n32, Y => n29
                           );
   U39 : NOR2X1 port map( A => state_1_port, B => state_0_port, Y => n30);
   U40 : NAND3X1 port map( A => n33, B => n34, C => n35, Y => nextstate_1_port)
                           ;
   U41 : AOI22X1 port map( A => n36, B => n18, C => n31, D => n37, Y => n35);
   U42 : INVX1 port map( A => n38, Y => n36);
   U43 : NAND3X1 port map( A => n39, B => n40, C => p_ready, Y => n33);
   U44 : NAND3X1 port map( A => n41, B => n28, C => n42, Y => nextstate_0_port)
                           ;
   U45 : AOI21X1 port map( A => n18, B => n38, C => n43, Y => n42);
   U46 : OAI21X1 port map( A => n44, B => n27, C => n45, Y => n43);
   U47 : NAND3X1 port map( A => p_ready, B => n37, C => n31, Y => n45);
   U48 : AND2X1 port map( A => n46, B => n47, Y => n31);
   U49 : INVX1 port map( A => n48, Y => n44);
   U50 : NAND3X1 port map( A => n19, B => n11, C => count_0_port, Y => n38);
   U51 : INVX1 port map( A => n49, Y => n28);
   U52 : AND2X1 port map( A => n26, B => n25, Y => n41);
   U53 : OAI21X1 port map( A => n50, B => n51, C => n52, Y => next_byte);
   U54 : MUX2X1 port map( B => n53, A => n54, S => n55, Y => n152);
   U55 : INVX1 port map( A => n56, Y => n153);
   U56 : MUX2X1 port map( B => PRGA_OUT(6), A => flop_data_6_port, S => n55, Y 
                           => n56);
   U57 : INVX1 port map( A => n57, Y => n154);
   U58 : MUX2X1 port map( B => PRGA_OUT(5), A => flop_data_5_port, S => n55, Y 
                           => n57);
   U59 : INVX1 port map( A => n58, Y => n155);
   U60 : MUX2X1 port map( B => PRGA_OUT(4), A => flop_data_4_port, S => n55, Y 
                           => n58);
   U61 : INVX1 port map( A => n59_port, Y => n156);
   U62 : MUX2X1 port map( B => PRGA_OUT(3), A => flop_data_3_port, S => n55, Y 
                           => n59_port);
   U63 : INVX1 port map( A => n60_port, Y => n157);
   U64 : MUX2X1 port map( B => PRGA_OUT(2), A => flop_data_2_port, S => n55, Y 
                           => n60_port);
   U65 : INVX1 port map( A => n61_port, Y => n174);
   U66 : MUX2X1 port map( B => PRGA_OUT(1), A => flop_data_1_port, S => n55, Y 
                           => n61_port);
   U67 : INVX1 port map( A => n62_port, Y => n175);
   U68 : MUX2X1 port map( B => PRGA_OUT(0), A => flop_data_0_port, S => n55, Y 
                           => n62_port);
   U69 : NAND3X1 port map( A => n63_port, B => n23, C => n64_port, Y => n55);
   U70 : AND2X1 port map( A => n24, B => n52, Y => n64_port);
   U71 : MUX2X1 port map( B => n65_port, A => n66, S => n40, Y => n52);
   U72 : NOR2X1 port map( A => p_ready, B => n67, Y => n66);
   U73 : NOR2X1 port map( A => n14, B => n65_port, Y => n63_port);
   U74 : INVX1 port map( A => t_bitstuff, Y => r81_B_0_port);
   U75 : OAI21X1 port map( A => n20, B => n68, C => n69, Y => n200);
   U76 : AOI22X1 port map( A => N59, B => n70, C => N84, D => n71, Y => n69);
   U77 : OAI21X1 port map( A => n11, B => n68, C => n72, Y => n199);
   U78 : AOI22X1 port map( A => N65, B => n70, C => N90, D => n71, Y => n72);
   U79 : OAI21X1 port map( A => n73, B => n68, C => n74, Y => n198);
   U80 : AOI22X1 port map( A => N64, B => n70, C => N89, D => n71, Y => n74);
   U81 : OAI21X1 port map( A => n75, B => n68, C => n76, Y => n197);
   U82 : AOI22X1 port map( A => N63, B => n70, C => N88, D => n71, Y => n76);
   U83 : OAI21X1 port map( A => n77, B => n68, C => n78, Y => n196);
   U84 : AOI22X1 port map( A => N62, B => n70, C => N87, D => n71, Y => n78);
   U85 : OAI21X1 port map( A => n79, B => n68, C => n80, Y => n195);
   U86 : AOI22X1 port map( A => N61, B => n70, C => N86, D => n71, Y => n80);
   U87 : OAI21X1 port map( A => n81, B => n68, C => n82, Y => n194);
   U88 : AOI22X1 port map( A => N60, B => n70, C => N85, D => n71, Y => n82);
   U89 : OAI21X1 port map( A => n32, B => n51, C => n34, Y => n71);
   U90 : OR2X1 port map( A => n25, B => n48, Y => n34);
   U91 : NAND3X1 port map( A => state_0_port, B => n83, C => state_1_port, Y =>
                           n25);
   U92 : INVX1 port map( A => n37, Y => n32);
   U93 : NAND2X1 port map( A => n48, B => n50, Y => n37);
   U94 : AND2X1 port map( A => prga_opcode(1), B => prga_opcode(0), Y => n50);
   U95 : AND2X1 port map( A => n68, B => n84_port, Y => n70);
   U96 : OAI21X1 port map( A => n48, B => n27, C => n85_port, Y => n84_port);
   U97 : NOR2X1 port map( A => n18, B => n49, Y => n85_port);
   U98 : NOR2X1 port map( A => n86_port, B => n87_port, Y => n48);
   U99 : NAND3X1 port map( A => count_4_port, B => count_1_port, C => 
                           count_5_port, Y => n87_port);
   U100 : NAND3X1 port map( A => count_0_port, B => count_3_port, C => n88_port
                           , Y => n86_port);
   U101 : NOR2X1 port map( A => N188, B => n79, Y => n88_port);
   U102 : NAND2X1 port map( A => n18, B => t_bitstuff, Y => n68);
   U103 : INVX1 port map( A => count_1_port, Y => n81);
   U104 : OAI21X1 port map( A => n89_port, B => n90_port, C => n91, Y => n173);
   U105 : INVX1 port map( A => current_send_data_7_port, Y => n90_port);
   U106 : OAI21X1 port map( A => n89_port, B => n92, C => n93, Y => n172);
   U107 : INVX1 port map( A => current_send_data_6_port, Y => n92);
   U108 : OAI21X1 port map( A => n89_port, B => n94, C => n95, Y => n171);
   U109 : INVX1 port map( A => current_send_data_5_port, Y => n94);
   U110 : OAI21X1 port map( A => n89_port, B => n96, C => n97, Y => n170);
   U111 : INVX1 port map( A => current_send_data_4_port, Y => n96);
   U112 : OAI21X1 port map( A => n89_port, B => n98, C => n99, Y => n169);
   U113 : INVX1 port map( A => current_send_data_3_port, Y => n98);
   U114 : OAI21X1 port map( A => n89_port, B => n100, C => n101, Y => n168);
   U115 : INVX1 port map( A => current_send_data_2_port, Y => n100);
   U116 : OAI21X1 port map( A => n89_port, B => n102, C => n103, Y => n167);
   U117 : INVX1 port map( A => current_send_data_1_port, Y => n102);
   U118 : OAI21X1 port map( A => n89_port, B => n104, C => n105, Y => n166);
   U119 : INVX1 port map( A => current_send_data_0_port, Y => n104);
   U120 : AOI21X1 port map( A => state_0_port, B => state_1_port, C => n13, Y 
                           => n89_port);
   U121 : NAND2X1 port map( A => n106, B => n91, Y => n165);
   U122 : NOR2X1 port map( A => n107, B => n108, Y => n91);
   U123 : OAI21X1 port map( A => n53, B => n109, C => n110, Y => n108);
   U124 : NAND2X1 port map( A => t_crc(15), B => n111, Y => n110);
   U125 : INVX1 port map( A => n112, Y => n109);
   U126 : INVX1 port map( A => PRGA_OUT(7), Y => n53);
   U127 : OAI22X1 port map( A => n54, B => n113, C => n114, D => n115, Y => 
                           n107);
   U128 : NAND2X1 port map( A => n116, B => state_0_port, Y => n115);
   U129 : OAI21X1 port map( A => N188, B => t_crc(7), C => n15, Y => n114);
   U130 : INVX1 port map( A => n117, Y => n113);
   U131 : INVX1 port map( A => flop_data_7_port, Y => n54);
   U132 : AOI22X1 port map( A => n118, B => current_send_data_7_port, C => 
                           send_data_7_port, D => n12, Y => n106);
   U133 : NAND2X1 port map( A => n119, B => n93, Y => n164);
   U134 : AND2X1 port map( A => n120, B => n121, Y => n93);
   U135 : AOI22X1 port map( A => t_crc(6), B => n122, C => n117, D => 
                           flop_data_6_port, Y => n121);
   U136 : AOI22X1 port map( A => t_crc(14), B => n111, C => n112, D => 
                           PRGA_OUT(6), Y => n120);
   U137 : AOI22X1 port map( A => n118, B => current_send_data_6_port, C => 
                           send_data_6_port, D => n12, Y => n119);
   U138 : NAND2X1 port map( A => n123, B => n95, Y => n163);
   U139 : AND2X1 port map( A => n124, B => n125, Y => n95);
   U140 : AOI22X1 port map( A => t_crc(5), B => n122, C => n117, D => 
                           flop_data_5_port, Y => n125);
   U141 : AOI22X1 port map( A => t_crc(13), B => n111, C => n112, D => 
                           PRGA_OUT(5), Y => n124);
   U142 : AOI22X1 port map( A => n118, B => current_send_data_5_port, C => 
                           send_data_5_port, D => n13, Y => n123);
   U143 : NAND2X1 port map( A => n126, B => n97, Y => n162);
   U144 : AND2X1 port map( A => n127, B => n128, Y => n97);
   U145 : AOI22X1 port map( A => t_crc(4), B => n122, C => n117, D => 
                           flop_data_4_port, Y => n128);
   U146 : AOI22X1 port map( A => t_crc(12), B => n111, C => n112, D => 
                           PRGA_OUT(4), Y => n127);
   U147 : AOI22X1 port map( A => n118, B => current_send_data_4_port, C => 
                           send_data_4_port, D => n13, Y => n126);
   U148 : NAND2X1 port map( A => n129, B => n99, Y => n161);
   U149 : AND2X1 port map( A => n130, B => n131, Y => n99);
   U150 : AOI22X1 port map( A => t_crc(3), B => n122, C => n117, D => 
                           flop_data_3_port, Y => n131);
   U151 : AOI22X1 port map( A => t_crc(11), B => n111, C => n112, D => 
                           PRGA_OUT(3), Y => n130);
   U152 : AOI22X1 port map( A => n118, B => current_send_data_3_port, C => 
                           send_data_3_port, D => n13, Y => n129);
   U153 : NAND2X1 port map( A => n132, B => n101, Y => n160);
   U154 : AND2X1 port map( A => n133, B => n134, Y => n101);
   U155 : AOI22X1 port map( A => t_crc(2), B => n122, C => n117, D => 
                           flop_data_2_port, Y => n134);
   U156 : AOI22X1 port map( A => t_crc(10), B => n111, C => n112, D => 
                           PRGA_OUT(2), Y => n133);
   U157 : AOI22X1 port map( A => n118, B => current_send_data_2_port, C => 
                           send_data_2_port, D => n13, Y => n132);
   U158 : NAND2X1 port map( A => n135, B => n103, Y => n159);
   U159 : AND2X1 port map( A => n136, B => n137, Y => n103);
   U160 : AOI22X1 port map( A => t_crc(1), B => n122, C => n117, D => 
                           flop_data_1_port, Y => n137);
   U161 : AOI22X1 port map( A => t_crc(9), B => n111, C => n112, D => 
                           PRGA_OUT(1), Y => n136);
   U162 : AOI22X1 port map( A => n118, B => current_send_data_1_port, C => 
                           send_data_1_port, D => n13, Y => n135);
   U163 : NAND2X1 port map( A => n138, B => n105, Y => n158);
   U164 : AND2X1 port map( A => n139, B => n140, Y => n105);
   U165 : AOI22X1 port map( A => t_crc(0), B => n122, C => n117, D => 
                           flop_data_0_port, Y => n140);
   U166 : NOR2X1 port map( A => n24, B => n13, Y => n117);
   U167 : NOR2X1 port map( A => n46, B => n18, Y => n24);
   U168 : NOR2X1 port map( A => n40, B => n67, Y => n18);
   U169 : INVX1 port map( A => n39, Y => n67);
   U170 : NOR2X1 port map( A => state_1_port, B => state_2_port, Y => n39);
   U171 : INVX1 port map( A => n51, Y => n46);
   U172 : INVX1 port map( A => n141, Y => n122);
   U173 : NAND3X1 port map( A => n116, B => state_0_port, C => n142, Y => n141)
                           ;
   U174 : NOR2X1 port map( A => n14, B => N188, Y => n142);
   U175 : AOI22X1 port map( A => t_crc(8), B => n111, C => n112, D => 
                           PRGA_OUT(0), Y => n139);
   U176 : NOR2X1 port map( A => n26, B => n13, Y => n112);
   U177 : NAND2X1 port map( A => n65_port, B => n40, Y => n26);
   U178 : NOR2X1 port map( A => n83, B => n143, Y => n65_port);
   U179 : INVX1 port map( A => state_1_port, Y => n143);
   U180 : NOR2X1 port map( A => n27, B => n14, Y => n111);
   U181 : NAND2X1 port map( A => n116, B => n40, Y => n27);
   U182 : AOI22X1 port map( A => n118, B => current_send_data_0_port, C => 
                           send_data_0_port, D => n12, Y => n138);
   U183 : INVX1 port map( A => n144, Y => n118);
   U184 : NAND3X1 port map( A => state_0_port, B => n15, C => state_1_port, Y 
                           => n144);
   U185 : OAI21X1 port map( A => n51, B => n47, C => n145, Y => EOP);
   U186 : NAND3X1 port map( A => N188, B => n146, C => n49, Y => n145);
   U187 : NOR2X1 port map( A => n23, B => n147, Y => n49);
   U188 : OAI21X1 port map( A => n148, B => n149, C => state_0_port, Y => n147)
                           ;
   U189 : NAND3X1 port map( A => count_2_port, B => N188, C => count_3_port, Y 
                           => n149);
   U190 : NAND3X1 port map( A => n75, B => n73, C => n150, Y => n148);
   U191 : NOR2X1 port map( A => count_1_port, B => count_0_port, Y => n150);
   U192 : INVX1 port map( A => count_5_port, Y => n73);
   U193 : INVX1 port map( A => count_4_port, Y => n75);
   U194 : INVX1 port map( A => n116, Y => n23);
   U195 : NOR2X1 port map( A => n83, B => state_1_port, Y => n116);
   U196 : NAND3X1 port map( A => n19, B => n20, C => N188, Y => n47);
   U197 : INVX1 port map( A => count_0_port, Y => n20);
   U198 : NOR2X1 port map( A => n146, B => count_1_port, Y => n19);
   U199 : NAND3X1 port map( A => n79, B => n77, C => n151, Y => n146);
   U200 : NOR2X1 port map( A => count_5_port, B => count_4_port, Y => n151);
   U201 : INVX1 port map( A => count_3_port, Y => n77);
   U202 : INVX1 port map( A => count_2_port, Y => n79);
   U203 : NAND3X1 port map( A => n40, B => n83, C => state_1_port, Y => n51);
   U204 : INVX1 port map( A => state_2_port, Y => n83);
   U205 : INVX1 port map( A => state_0_port, Y => n40);

end SYN_behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_shiftreg_1 is

   port( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe : in std_logic;  
         send_data : in std_logic_vector (7 downto 0);  d_encode : out 
         std_logic);

end tx_shiftreg_1;

architecture SYN_dataflow of tx_shiftreg_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal d_encode_port, present_val_7_port, present_val_6_port, 
      present_val_5_port, present_val_4_port, present_val_3_port, 
      present_val_2_port, present_val_1_port, count_2_port, count_1_port, 
      count_0_port, n9, n10, n12, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n1, n2, n3, n4, n5, n6, n7, n8, n11, n13, n14, n15, n16, n17,
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n54 : std_logic;

begin
   d_encode <= d_encode_port;
   
   count_reg_0_inst : DFFSR port map( D => n53, CLK => clk, R => n12, S => n14,
                           Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => n51, CLK => clk, R => n10, S => n14,
                           Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n52, CLK => clk, R => n9, S => n14, 
                           Q => count_2_port);
   n9 <= '1';
   n10 <= '1';
   n12 <= '1';
   U30 : OAI21X1 port map( A => n13, B => n54, C => n29, Y => n43);
   U31 : AOI22X1 port map( A => send_data(0), B => n17, C => present_val_1_port
                           , D => n15, Y => n29);
   U32 : OAI21X1 port map( A => n13, B => n21, C => n30, Y => n44);
   U33 : NAND2X1 port map( A => send_data(7), B => n17, Y => n30);
   U34 : OAI21X1 port map( A => n13, B => n22, C => n31, Y => n45);
   U35 : AOI22X1 port map( A => send_data(6), B => n17, C => present_val_7_port
                           , D => n15, Y => n31);
   U36 : OAI21X1 port map( A => n13, B => n23, C => n32, Y => n46);
   U37 : AOI22X1 port map( A => send_data(5), B => n17, C => present_val_6_port
                           , D => n15, Y => n32);
   U38 : OAI21X1 port map( A => n13, B => n24, C => n33, Y => n47);
   U39 : AOI22X1 port map( A => send_data(4), B => n17, C => present_val_5_port
                           , D => n15, Y => n33);
   U40 : OAI21X1 port map( A => n13, B => n25, C => n34, Y => n48);
   U41 : AOI22X1 port map( A => send_data(3), B => n17, C => present_val_4_port
                           , D => n15, Y => n34);
   U42 : OAI21X1 port map( A => n13, B => n26, C => n35, Y => n49);
   U43 : AOI22X1 port map( A => send_data(2), B => n17, C => present_val_3_port
                           , D => n15, Y => n35);
   U44 : OAI21X1 port map( A => n27, B => n13, C => n36, Y => n50);
   U45 : AOI22X1 port map( A => send_data(1), B => n17, C => present_val_2_port
                           , D => n15, Y => n36);
   U46 : OAI21X1 port map( A => n37, B => n38, C => n39, Y => n51);
   U47 : OAI21X1 port map( A => n18, B => n11, C => count_1_port, Y => n39);
   U48 : NAND2X1 port map( A => count_0_port, B => n19, Y => n38);
   U49 : OAI21X1 port map( A => n17, B => n20, C => n40, Y => n52);
   U50 : NAND3X1 port map( A => count_1_port, B => count_0_port, C => n15, Y =>
                           n40);
   U51 : OAI22X1 port map( A => n18, B => n13, C => count_0_port, D => n37, Y 
                           => n53);
   U52 : NAND2X1 port map( A => n13, B => n41, Y => n37);
   U53 : OAI21X1 port map( A => t_bitstuff, B => n16, C => n41, Y => n28);
   U54 : NAND3X1 port map( A => SHIFT_ENABLE_R, B => count_0_port, C => n42, Y 
                           => n41);
   U55 : NOR2X1 port map( A => n19, B => n20, Y => n42);
   present_val_reg_7_inst : DFFSR port map( D => n44, CLK => clk, R => n14, S 
                           => n8, Q => present_val_7_port);
   present_val_reg_1_inst : DFFSR port map( D => n50, CLK => clk, R => n14, S 
                           => n7, Q => present_val_1_port);
   present_val_reg_6_inst : DFFSR port map( D => n45, CLK => clk, R => n14, S 
                           => n6, Q => present_val_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n46, CLK => clk, R => n14, S 
                           => n5, Q => present_val_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n47, CLK => clk, R => n14, S 
                           => n4, Q => present_val_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n48, CLK => clk, R => n14, S 
                           => n3, Q => present_val_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n49, CLK => clk, R => n14, S 
                           => n2, Q => present_val_2_port);
   present_val_reg_0_inst : DFFSR port map( D => n43, CLK => clk, R => n14, S 
                           => n1, Q => d_encode_port);
   U3 : INVX4 port map( A => n11, Y => n13);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   U15 : INVX2 port map( A => rst, Y => n14);
   U16 : INVX2 port map( A => n41, Y => n17);
   U17 : INVX2 port map( A => n28, Y => n11);
   U18 : INVX2 port map( A => n37, Y => n15);
   U19 : INVX2 port map( A => SHIFT_ENABLE_R, Y => n16);
   U20 : INVX2 port map( A => count_0_port, Y => n18);
   U21 : INVX2 port map( A => count_1_port, Y => n19);
   U22 : INVX2 port map( A => count_2_port, Y => n20);
   U23 : INVX2 port map( A => present_val_7_port, Y => n21);
   U24 : INVX2 port map( A => present_val_6_port, Y => n22);
   U25 : INVX2 port map( A => present_val_5_port, Y => n23);
   U26 : INVX2 port map( A => present_val_4_port, Y => n24);
   U27 : INVX2 port map( A => present_val_3_port, Y => n25);
   U28 : INVX2 port map( A => present_val_2_port, Y => n26);
   U29 : INVX2 port map( A => present_val_1_port, Y => n27);
   U56 : INVX2 port map( A => d_encode_port, Y => n54);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_encode_1 is

   port( clk, rst, SHIFT_ENABLE_E, d_encode, EOP : in std_logic;  t_bitstuff, 
         dp_tx_out, dm_tx_out : out std_logic);

end tx_encode_1;

architecture SYN_moore of tx_encode_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal DE_holdout, DE_holdout_BS, state_3_port, state_2_port, state_1_port, 
      state_0_port, nextstate_3_port, nextstate_2_port, nextstate_1_port, 
      nextstate_0_port, DE_holdout_last, DE_holdout_nxt, dm_tx_nxt, n1, n3, n5,
      n6, n9, n12, n13, n14, n15, n18, n19, n20, n22, n23, n24, n26, n27, n32, 
      n33, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n55, n61, n62, n64, n2, n4, n7, n8, n10, n11, n16, n17, n21, 
      n25, n28, n29, n30, n31, n34, n35, n42, n53, n54, n56, n57, n58, n59, n60
      , n63 : std_logic;

begin
   
   DE_holdout_reg : DFFSR port map( D => DE_holdout_nxt, CLK => clk, R => n62, 
                           S => n16, Q => DE_holdout);
   DE_holdout_last_reg : DFFPOSX1 port map( D => n61, CLK => clk, Q => 
                           DE_holdout_last);
   dp_tx_out_reg : DFFSR port map( D => DE_holdout_nxt, CLK => clk, R => n55, S
                           => n16, Q => dp_tx_out);
   U3 : AOI21X1 port map( A => state_3_port, B => n1, C => n30, Y => 
                           nextstate_3_port);
   U4 : OAI21X1 port map( A => n3, B => n60, C => n5, Y => nextstate_2_port);
   U5 : AOI21X1 port map( A => n6, B => n17, C => n34, Y => n5);
   U7 : NOR2X1 port map( A => state_2_port, B => n59, Y => n6);
   U8 : AOI21X1 port map( A => n35, B => n59, C => n12, Y => n3);
   U9 : OAI21X1 port map( A => state_1_port, B => n9, C => n13, Y => 
                           nextstate_1_port);
   U10 : AOI21X1 port map( A => state_1_port, B => n14, C => n34, Y => n13);
   U11 : OAI21X1 port map( A => state_0_port, B => n15, C => n21, Y => n14);
   U12 : NAND3X1 port map( A => SHIFT_ENABLE_E, B => n35, C => state_0_port, Y 
                           => n9);
   U14 : OAI21X1 port map( A => n58, B => n21, C => n18, Y => nextstate_0_port)
                           ;
   U15 : OAI21X1 port map( A => n19, B => n20, C => SHIFT_ENABLE_E, Y => n18);
   U16 : OAI21X1 port map( A => n31, B => n22, C => n23, Y => n20);
   U17 : NAND2X1 port map( A => n24, B => n42, Y => n22);
   U18 : NOR2X1 port map( A => state_0_port, B => n15, Y => n19);
   U19 : NAND3X1 port map( A => d_encode, B => n26, C => n27, Y => n15);
   U20 : XNOR2X1 port map( A => n54, B => n53, Y => n27);
   U22 : NOR2X1 port map( A => n31, B => SHIFT_ENABLE_E, Y => n12);
   U23 : OAI22X1 port map( A => n16, B => n54, C => rst, D => n53, Y => n61);
   U26 : OAI22X1 port map( A => n25, B => n63, C => n53, D => n32, Y => n64);
   U28 : NAND2X1 port map( A => n34, B => SHIFT_ENABLE_E, Y => n32);
   U30 : NAND3X1 port map( A => n24, B => n58, C => n26, Y => n23);
   U31 : NOR2X1 port map( A => state_3_port, B => n33, Y => t_bitstuff);
   U32 : OAI21X1 port map( A => n57, B => n56, C => n36, Y => dm_tx_nxt);
   U33 : AOI22X1 port map( A => n37, B => n24, C => n38, D => n39, Y => n36);
   U34 : NOR2X1 port map( A => n24, B => n31, Y => n38);
   U36 : NOR2X1 port map( A => EOP, B => state_3_port, Y => n26);
   U37 : NOR2X1 port map( A => EOP, B => n40, Y => n37);
   U38 : AOI22X1 port map( A => state_0_port, B => n41, C => n28, D => n58, Y 
                           => n40);
   U40 : XNOR2X1 port map( A => DE_holdout_BS, B => n44, Y => n41);
   U41 : OAI21X1 port map( A => n57, B => n56, C => n45, Y => DE_holdout_nxt);
   U42 : OAI21X1 port map( A => n46, B => n47, C => n30, Y => n45);
   U44 : OAI21X1 port map( A => n24, B => n39, C => n48, Y => n47);
   U45 : NAND3X1 port map( A => n43, B => n58, C => n24, Y => n48);
   U46 : XOR2X1 port map( A => DE_holdout, B => SHIFT_ENABLE_E, Y => n43);
   U47 : XNOR2X1 port map( A => n49, B => n53, Y => n39);
   U49 : NAND2X1 port map( A => SHIFT_ENABLE_E, B => n42, Y => n49);
   U51 : OAI21X1 port map( A => n33, B => n50, C => n51, Y => n46);
   U52 : AOI21X1 port map( A => n52, B => n29, C => state_3_port, Y => n51);
   U54 : NOR2X1 port map( A => n63, B => n33, Y => n52);
   U55 : NAND2X1 port map( A => n44, B => n63, Y => n50);
   U57 : NAND2X1 port map( A => SHIFT_ENABLE_E, B => d_encode, Y => n44);
   U58 : NAND2X1 port map( A => state_0_port, B => n24, Y => n33);
   U59 : NOR2X1 port map( A => n60, B => n59, Y => n24);
   U62 : NAND3X1 port map( A => n59, B => n60, C => n58, Y => n1);
   n55 <= '1';
   n62 <= '1';
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => clk, R => 
                           n16, S => n11, Q => state_3_port);
   dm_tx_out_reg : DFFSR port map( D => dm_tx_nxt, CLK => clk, R => n16, S => 
                           n10, Q => dm_tx_out);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n16, S => n8, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n16, S => n7, Q => state_1_port);
   DE_holdout_BS_reg : DFFSR port map( D => n64, CLK => clk, R => n16, S => n4,
                           Q => DE_holdout_BS);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n16, S => n2, Q => state_2_port);
   n2 <= '1';
   n4 <= '1';
   n7 <= '1';
   n8 <= '1';
   n10 <= '1';
   n11 <= '1';
   U29 : INVX2 port map( A => rst, Y => n16);
   U35 : INVX2 port map( A => n9, Y => n17);
   U39 : INVX2 port map( A => n12, Y => n21);
   U43 : INVX2 port map( A => n32, Y => n25);
   U48 : INVX2 port map( A => n43, Y => n28);
   U50 : INVX2 port map( A => n44, Y => n29);
   U53 : INVX2 port map( A => EOP, Y => n30);
   U56 : INVX2 port map( A => n26, Y => n31);
   U60 : INVX2 port map( A => n23, Y => n34);
   U61 : INVX2 port map( A => n15, Y => n35);
   U63 : INVX2 port map( A => d_encode, Y => n42);
   U64 : INVX2 port map( A => DE_holdout, Y => n53);
   U65 : INVX2 port map( A => DE_holdout_last, Y => n54);
   U66 : INVX2 port map( A => state_3_port, Y => n56);
   U68 : INVX2 port map( A => n1, Y => n57);
   U69 : INVX2 port map( A => state_0_port, Y => n58);
   U70 : INVX2 port map( A => state_1_port, Y => n59);
   U71 : INVX2 port map( A => state_2_port, Y => n60);
   U72 : INVX2 port map( A => DE_holdout_BS, Y => n63);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity tx_CRC_CALC_1 is

   port( CLK, RST, EOP, T_STROBE : in std_logic;  PRGA_OPCODE : in 
         std_logic_vector (1 downto 0);  PRGA_OUT : in std_logic_vector (7 
         downto 0);  TX_CRC : out std_logic_vector (15 downto 0));

end tx_CRC_CALC_1;

architecture SYN_txcrcm of tx_CRC_CALC_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal TX_CRC_15_port, TX_CRC_14_port, TX_CRC_13_port, TX_CRC_12_port, 
      TX_CRC_11_port, TX_CRC_10_port, TX_CRC_9_port, TX_CRC_8_port, 
      TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port, TX_CRC_4_port, TX_CRC_3_port
      , TX_CRC_2_port, TX_CRC_1_port, TX_CRC_0_port, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n79, 
      n80, n81 : std_logic;

begin
   TX_CRC <= ( TX_CRC_15_port, TX_CRC_14_port, TX_CRC_13_port, TX_CRC_12_port, 
      TX_CRC_11_port, TX_CRC_10_port, TX_CRC_9_port, TX_CRC_8_port, 
      TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port, TX_CRC_4_port, TX_CRC_3_port
      , TX_CRC_2_port, TX_CRC_1_port, TX_CRC_0_port );
   
   U39 : OAI22X1 port map( A => n25, B => n20, C => n38, D => n19, Y => n63);
   U40 : XNOR2X1 port map( A => n40, B => n80, Y => n38);
   U41 : OAI22X1 port map( A => n79, B => n20, C => n19, D => n37, Y => n64);
   U42 : OAI22X1 port map( A => n36, B => n20, C => n19, D => n35, Y => n65);
   U43 : OAI22X1 port map( A => n34, B => n20, C => n19, D => n33, Y => n66);
   U44 : OAI22X1 port map( A => n32, B => n20, C => n19, D => n31, Y => n67);
   U45 : OAI22X1 port map( A => n29, B => n20, C => n19, D => n28, Y => n68);
   U46 : OAI22X1 port map( A => n27, B => n20, C => n41, D => n19, Y => n69);
   U47 : XNOR2X1 port map( A => TX_CRC_1_port, B => n42, Y => n41);
   U48 : OAI22X1 port map( A => n24, B => n20, C => n43, D => n19, Y => n70);
   U49 : XOR2X1 port map( A => n44, B => n45, Y => n43);
   U50 : XNOR2X1 port map( A => TX_CRC_0_port, B => n42, Y => n44);
   U51 : OAI22X1 port map( A => n80, B => n20, C => n46, D => n19, Y => n71);
   U52 : OAI22X1 port map( A => n20, B => n37, C => n47, D => n19, Y => n72);
   U53 : XNOR2X1 port map( A => n48, B => n49, Y => n47);
   U54 : OAI22X1 port map( A => n20, B => n35, C => n50, D => n39, Y => n73);
   U55 : OAI22X1 port map( A => n20, B => n33, C => n51, D => n39, Y => n74);
   U56 : XNOR2X1 port map( A => n52, B => n53, Y => n51);
   U57 : OAI22X1 port map( A => n20, B => n31, C => n54, D => n39, Y => n75);
   U58 : OAI22X1 port map( A => n20, B => n28, C => n55, D => n39, Y => n76);
   U59 : XOR2X1 port map( A => n56, B => n57, Y => n55);
   U60 : OAI22X1 port map( A => n20, B => n26, C => n58, D => n39, Y => n77);
   U61 : XOR2X1 port map( A => n59, B => n60, Y => n58);
   U62 : XOR2X1 port map( A => n42, B => n46, Y => n59);
   U63 : OAI22X1 port map( A => n20, B => n23, C => n40, D => n39, Y => n78);
   U64 : XOR2X1 port map( A => n61, B => n62, Y => n40);
   U65 : XOR2X1 port map( A => n57, B => n42, Y => n62);
   U66 : XNOR2X1 port map( A => n25, B => PRGA_OUT(7), Y => n42);
   U67 : XNOR2X1 port map( A => n24, B => PRGA_OUT(0), Y => n57);
   U68 : XOR2X1 port map( A => n46, B => n60, Y => n61);
   U69 : XOR2X1 port map( A => n54, B => n50, Y => n60);
   U70 : XNOR2X1 port map( A => n53, B => n48, Y => n50);
   U71 : XOR2X1 port map( A => TX_CRC_12_port, B => PRGA_OUT(4), Y => n48);
   U72 : XOR2X1 port map( A => TX_CRC_11_port, B => PRGA_OUT(3), Y => n53);
   U73 : XNOR2X1 port map( A => n56, B => n30, Y => n54);
   U74 : XOR2X1 port map( A => TX_CRC_10_port, B => PRGA_OUT(2), Y => n52);
   U75 : XNOR2X1 port map( A => TX_CRC_9_port, B => PRGA_OUT(1), Y => n56);
   U76 : XNOR2X1 port map( A => n49, B => n45, Y => n46);
   U77 : XNOR2X1 port map( A => n79, B => PRGA_OUT(6), Y => n45);
   U78 : XOR2X1 port map( A => TX_CRC_13_port, B => PRGA_OUT(5), Y => n49);
   U80 : NAND3X1 port map( A => PRGA_OPCODE(0), B => n81, C => T_STROBE, Y => 
                           n39);
   current_crc_reg_6_inst : DFFSR port map( D => n72, CLK => CLK, R => n21, S 
                           => n17, Q => TX_CRC_6_port);
   current_crc_reg_5_inst : DFFSR port map( D => n73, CLK => CLK, R => n21, S 
                           => n16, Q => TX_CRC_5_port);
   current_crc_reg_4_inst : DFFSR port map( D => n74, CLK => CLK, R => n21, S 
                           => n15, Q => TX_CRC_4_port);
   current_crc_reg_3_inst : DFFSR port map( D => n75, CLK => CLK, R => n21, S 
                           => n14, Q => TX_CRC_3_port);
   current_crc_reg_2_inst : DFFSR port map( D => n76, CLK => CLK, R => n21, S 
                           => n13, Q => TX_CRC_2_port);
   current_crc_reg_1_inst : DFFSR port map( D => n77, CLK => CLK, R => n21, S 
                           => n12, Q => TX_CRC_1_port);
   current_crc_reg_0_inst : DFFSR port map( D => n78, CLK => CLK, R => n21, S 
                           => n11, Q => TX_CRC_0_port);
   current_crc_reg_15_inst : DFFSR port map( D => n63, CLK => CLK, R => n21, S 
                           => n10, Q => TX_CRC_15_port);
   current_crc_reg_14_inst : DFFSR port map( D => n64, CLK => CLK, R => n21, S 
                           => n9, Q => TX_CRC_14_port);
   current_crc_reg_13_inst : DFFSR port map( D => n65, CLK => CLK, R => n21, S 
                           => n8, Q => TX_CRC_13_port);
   current_crc_reg_12_inst : DFFSR port map( D => n66, CLK => CLK, R => n21, S 
                           => n7, Q => TX_CRC_12_port);
   current_crc_reg_11_inst : DFFSR port map( D => n67, CLK => CLK, R => n21, S 
                           => n6, Q => TX_CRC_11_port);
   current_crc_reg_10_inst : DFFSR port map( D => n68, CLK => CLK, R => n21, S 
                           => n5, Q => TX_CRC_10_port);
   current_crc_reg_9_inst : DFFSR port map( D => n69, CLK => CLK, R => n21, S 
                           => n4, Q => TX_CRC_9_port);
   current_crc_reg_8_inst : DFFSR port map( D => n70, CLK => CLK, R => n21, S 
                           => n3, Q => TX_CRC_8_port);
   current_crc_reg_7_inst : DFFSR port map( D => n71, CLK => CLK, R => n21, S 
                           => n2, Q => TX_CRC_7_port);
   U3 : AND2X2 port map( A => n19, B => n22, Y => n1);
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   U20 : INVX2 port map( A => n1, Y => n20);
   U21 : INVX2 port map( A => RST, Y => n21);
   U22 : INVX2 port map( A => n18, Y => n19);
   U23 : INVX2 port map( A => n39, Y => n18);
   U24 : INVX2 port map( A => EOP, Y => n22);
   U25 : INVX2 port map( A => TX_CRC_0_port, Y => n23);
   U26 : INVX2 port map( A => TX_CRC_8_port, Y => n24);
   U27 : INVX2 port map( A => TX_CRC_15_port, Y => n25);
   U28 : INVX2 port map( A => TX_CRC_1_port, Y => n26);
   U29 : INVX2 port map( A => TX_CRC_9_port, Y => n27);
   U30 : INVX2 port map( A => TX_CRC_2_port, Y => n28);
   U31 : INVX2 port map( A => TX_CRC_10_port, Y => n29);
   U32 : INVX2 port map( A => n52, Y => n30);
   U33 : INVX2 port map( A => TX_CRC_3_port, Y => n31);
   U34 : INVX2 port map( A => TX_CRC_11_port, Y => n32);
   U35 : INVX2 port map( A => TX_CRC_4_port, Y => n33);
   U36 : INVX2 port map( A => TX_CRC_12_port, Y => n34);
   U37 : INVX2 port map( A => TX_CRC_5_port, Y => n35);
   U38 : INVX2 port map( A => TX_CRC_13_port, Y => n36);
   U79 : INVX2 port map( A => TX_CRC_6_port, Y => n37);
   U81 : INVX2 port map( A => TX_CRC_14_port, Y => n79);
   U82 : INVX2 port map( A => TX_CRC_7_port, Y => n80);
   U83 : INVX2 port map( A => PRGA_OPCODE(1), Y => n81);

end SYN_txcrcm;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_timer_1 is

   port( CLK, RST, D_EDGE, RCVING : in std_logic;  SHIFT_ENABLE : out std_logic
         );

end rx_timer_1;

architecture SYN_moore of rx_timer_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   signal count_3_port, count_2_port, count_1_port, count_0_port, state, 
      nextcount_3_port, nextcount_2_port, nextcount_1_port, nextcount_0_port, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n1, n2, n3, n4, n5
      , n6, n7, n8, n9, n10, n11, n12, n24, n25 : std_logic;

begin
   
   U9 : AND2X2 port map( A => n25, B => state, Y => n19);
   U17 : NOR2X1 port map( A => n13, B => n14, Y => nextcount_3_port);
   U18 : AOI22X1 port map( A => n15, B => n16, C => n17, D => count_3_port, Y 
                           => n13);
   U19 : XOR2X1 port map( A => n18, B => n16, Y => n17);
   U20 : NOR2X1 port map( A => count_3_port, B => n11, Y => n15);
   U21 : AOI21X1 port map( A => n19, B => n20, C => n24, Y => nextcount_2_port)
                           ;
   U22 : XOR2X1 port map( A => n21, B => count_2_port, Y => n20);
   U23 : NOR2X1 port map( A => n22, B => n14, Y => nextcount_1_port);
   U24 : NAND2X1 port map( A => state, B => n23, Y => nextcount_0_port);
   U25 : OAI21X1 port map( A => D_EDGE, B => n10, C => RCVING, Y => n23);
   U28 : NAND3X1 port map( A => RCVING, B => n25, C => state, Y => n14);
   U29 : OAI21X1 port map( A => n22, B => n12, C => n21, Y => n18);
   U30 : NAND2X1 port map( A => count_0_port, B => count_1_port, Y => n21);
   U31 : XOR2X1 port map( A => n12, B => n22, Y => n16);
   U32 : XNOR2X1 port map( A => count_0_port, B => count_1_port, Y => n22);
   state_reg : DFFSR port map( D => RCVING, CLK => CLK, R => n8, S => n5, Q => 
                           state);
   count_reg_2_inst : DFFSR port map( D => nextcount_2_port, CLK => CLK, R => 
                           n8, S => n4, Q => count_2_port);
   count_reg_0_inst : DFFSR port map( D => nextcount_0_port, CLK => CLK, R => 
                           n8, S => n3, Q => count_0_port);
   count_reg_3_inst : DFFSR port map( D => nextcount_3_port, CLK => CLK, R => 
                           n8, S => n2, Q => count_3_port);
   count_reg_1_inst : DFFSR port map( D => nextcount_1_port, CLK => CLK, R => 
                           n8, S => n1, Q => count_1_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   U8 : INVX2 port map( A => RST, Y => n8);
   U10 : AND2X2 port map( A => n6, B => n7, Y => SHIFT_ENABLE);
   U11 : NOR2X1 port map( A => n16, B => n18, Y => n6);
   U12 : AND2X2 port map( A => n9, B => count_3_port, Y => n7);
   U13 : INVX2 port map( A => n14, Y => n9);
   U14 : INVX2 port map( A => count_0_port, Y => n10);
   U15 : INVX2 port map( A => n18, Y => n11);
   U16 : INVX2 port map( A => count_2_port, Y => n12);
   U26 : INVX2 port map( A => RCVING, Y => n24);
   U27 : INVX2 port map( A => D_EDGE, Y => n25);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_shift_reg_1 is

   port( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF : in std_logic;  RCV_DATA : 
         out std_logic_vector (7 downto 0));

end rx_shift_reg_1;

architecture SYN_dataflow of rx_shift_reg_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      present_val_7_port, present_val_6_port, present_val_5_port, 
      present_val_4_port, present_val_3_port, present_val_2_port, 
      present_val_1_port, present_val_0_port, n2, n4, n6, n8, n10, n12, n14, 
      n16, n18, n19, n21, n23, n24, n26, n27, n29, n30, n32, n33, n35, n36, n38
      , n39, n41, n42, n44, n1, n3, n5, n7, n9, n11, n13, n15, n17, n20, n22, 
      n25, n28, n31, n34, n37, n40, n43, n45 : std_logic;

begin
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   
   RCV_DATA_reg_7_inst : DFFPOSX1 port map( D => n42, CLK => CLK, Q => 
                           RCV_DATA_7_port);
   RCV_DATA_reg_6_inst : DFFPOSX1 port map( D => n39, CLK => CLK, Q => 
                           RCV_DATA_6_port);
   RCV_DATA_reg_5_inst : DFFPOSX1 port map( D => n36, CLK => CLK, Q => 
                           RCV_DATA_5_port);
   RCV_DATA_reg_4_inst : DFFPOSX1 port map( D => n33, CLK => CLK, Q => 
                           RCV_DATA_4_port);
   RCV_DATA_reg_3_inst : DFFPOSX1 port map( D => n30, CLK => CLK, Q => 
                           RCV_DATA_3_port);
   RCV_DATA_reg_2_inst : DFFPOSX1 port map( D => n27, CLK => CLK, Q => 
                           RCV_DATA_2_port);
   RCV_DATA_reg_1_inst : DFFPOSX1 port map( D => n24, CLK => CLK, Q => 
                           RCV_DATA_1_port);
   RCV_DATA_reg_0_inst : DFFPOSX1 port map( D => n21, CLK => CLK, Q => 
                           RCV_DATA_0_port);
   U2 : OAI21X1 port map( A => RST, B => n43, C => n2, Y => n21);
   U3 : NAND2X1 port map( A => RCV_DATA_0_port, B => RST, Y => n2);
   U4 : OAI22X1 port map( A => n20, B => n43, C => n4, D => n40, Y => n23);
   U6 : OAI21X1 port map( A => RST, B => n40, C => n6, Y => n24);
   U7 : NAND2X1 port map( A => RCV_DATA_1_port, B => RST, Y => n6);
   U8 : OAI22X1 port map( A => n20, B => n40, C => n4, D => n37, Y => n26);
   U10 : OAI21X1 port map( A => RST, B => n37, C => n8, Y => n27);
   U11 : NAND2X1 port map( A => RCV_DATA_2_port, B => RST, Y => n8);
   U12 : OAI22X1 port map( A => n20, B => n37, C => n4, D => n34, Y => n29);
   U14 : OAI21X1 port map( A => RST, B => n34, C => n10, Y => n30);
   U15 : NAND2X1 port map( A => RCV_DATA_3_port, B => RST, Y => n10);
   U16 : OAI22X1 port map( A => n20, B => n34, C => n4, D => n31, Y => n32);
   U18 : OAI21X1 port map( A => RST, B => n31, C => n12, Y => n33);
   U19 : NAND2X1 port map( A => RCV_DATA_4_port, B => RST, Y => n12);
   U20 : OAI22X1 port map( A => n20, B => n31, C => n4, D => n28, Y => n35);
   U22 : OAI21X1 port map( A => RST, B => n28, C => n14, Y => n36);
   U23 : NAND2X1 port map( A => RCV_DATA_5_port, B => RST, Y => n14);
   U24 : OAI22X1 port map( A => n20, B => n28, C => n4, D => n25, Y => n38);
   U26 : OAI21X1 port map( A => RST, B => n25, C => n16, Y => n39);
   U27 : NAND2X1 port map( A => RCV_DATA_6_port, B => RST, Y => n16);
   U28 : OAI22X1 port map( A => n20, B => n25, C => n4, D => n22, Y => n41);
   U30 : OAI21X1 port map( A => RST, B => n22, C => n18, Y => n42);
   U31 : NAND2X1 port map( A => RCV_DATA_7_port, B => RST, Y => n18);
   U32 : OAI21X1 port map( A => n20, B => n22, C => n19, Y => n44);
   U33 : NAND2X1 port map( A => D_ORIG, B => n20, Y => n19);
   U36 : NAND2X1 port map( A => SHIFT_ENABLE, B => n45, Y => n4);
   present_val_reg_7_inst : DFFSR port map( D => n44, CLK => CLK, R => n17, S 
                           => n15, Q => present_val_7_port);
   present_val_reg_6_inst : DFFSR port map( D => n41, CLK => CLK, R => n17, S 
                           => n13, Q => present_val_6_port);
   present_val_reg_5_inst : DFFSR port map( D => n38, CLK => CLK, R => n17, S 
                           => n11, Q => present_val_5_port);
   present_val_reg_4_inst : DFFSR port map( D => n35, CLK => CLK, R => n17, S 
                           => n9, Q => present_val_4_port);
   present_val_reg_3_inst : DFFSR port map( D => n32, CLK => CLK, R => n17, S 
                           => n7, Q => present_val_3_port);
   present_val_reg_2_inst : DFFSR port map( D => n29, CLK => CLK, R => n17, S 
                           => n5, Q => present_val_2_port);
   present_val_reg_1_inst : DFFSR port map( D => n26, CLK => CLK, R => n17, S 
                           => n3, Q => present_val_1_port);
   present_val_reg_0_inst : DFFSR port map( D => n23, CLK => CLK, R => n17, S 
                           => n1, Q => present_val_0_port);
   U5 : INVX2 port map( A => n4, Y => n20);
   n1 <= '1';
   n3 <= '1';
   n5 <= '1';
   n7 <= '1';
   n9 <= '1';
   n11 <= '1';
   n13 <= '1';
   n15 <= '1';
   U37 : INVX2 port map( A => RST, Y => n17);
   U38 : INVX2 port map( A => present_val_7_port, Y => n22);
   U39 : INVX2 port map( A => present_val_6_port, Y => n25);
   U40 : INVX2 port map( A => present_val_5_port, Y => n28);
   U41 : INVX2 port map( A => present_val_4_port, Y => n31);
   U42 : INVX2 port map( A => present_val_3_port, Y => n34);
   U43 : INVX2 port map( A => present_val_2_port, Y => n37);
   U44 : INVX2 port map( A => present_val_1_port, Y => n40);
   U45 : INVX2 port map( A => present_val_0_port, Y => n43);
   U46 : INVX2 port map( A => BITSTUFF, Y => n45);

end SYN_dataflow;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_rcu_1 is

   port( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR : in std_logic
         ;  RX_CRC, RX_CHECK_CRC : in std_logic_vector (15 downto 0);  RCV_DATA
         : in std_logic_vector (7 downto 0);  RCVING, W_ENABLE, R_ERROR, 
         CRC_ERROR : out std_logic;  OPCODE : out std_logic_vector (1 downto 0)
         );

end rx_rcu_1;

architecture SYN_moore of rx_rcu_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal CRC_ERROR_port, n192, state_3_port, state_2_port, state_1_port, 
      state_0_port, count_3_port, count_2_port, count_1_port, count_0_port, 
      nextstate_3_port, nextstate_2_port, nextstate_1_port, nextstate_0_port, 
      nxtR_ERROR, curR_ERROR, curCRC_ERROR, n9, n11, n12, n14, n15, n16, n20, 
      n21, n22, n27, n29, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41, n42
      , n45, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n59, n60, 
      n61, n62, n63, n65, n66, n67, n70, n71, n72, n74, n75, n77, n78, n79, n80
      , n81, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95, n96, 
      n97, n98, n99, n100, n102, n103, n105, n106, n107, n109, n111, n113, n116
      , n117, n119, n120, n121, n122, n123, n125, n126, n127, n129, n133, n134,
      n136, n137, n138, n139, n140, n142, n144, n145, n146, n147, n150, n151, 
      n161, n162, n163, n1, n2, n3, n4, n5, n6, n7, n8, n10, n13, n17, n18, n19
      , n23, n24, n25, n28, n30, n35, n43, n44, n49, n58, n64, n68, n69, n73, 
      n76, n82, n93, n101, n104, n108, n110, n112, n114, n115, n118, n124, n128
      , n130, n131, n132, n135, n141, n143, n148, n149, n152, n153, n154, n155,
      n156, n157, n158, n159, n160, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191 : std_logic;

begin
   CRC_ERROR <= CRC_ERROR_port;
   
   curCRC_ERROR_reg : DFFPOSX1 port map( D => n151, CLK => CLK, Q => 
                           curCRC_ERROR);
   curR_ERROR_reg : DFFPOSX1 port map( D => n150, CLK => CLK, Q => curR_ERROR);
   CRC_ERROR_reg : DFFPOSX1 port map( D => n169, CLK => CLK, Q => 
                           CRC_ERROR_port);
   U5 : OAI21X1 port map( A => EOP, B => n43, C => n14, Y => n12);
   U6 : AOI22X1 port map( A => BS_ERROR, B => n15, C => n16, D => n30, Y => n14
                           );
   U7 : OAI21X1 port map( A => n191, B => n25, C => n20, Y => n16);
   U8 : AOI22X1 port map( A => n21, B => D_EDGE, C => n1, D => n22, Y => n20);
   U9 : OAI21X1 port map( A => n181, B => n189, C => n182, Y => n22);
   U11 : NOR2X1 port map( A => n181, B => n175, Y => n21);
   U12 : OAI21X1 port map( A => n27, B => n183, C => n29, Y => n15);
   U13 : OAI21X1 port map( A => n3, B => n31, C => n32, Y => n11);
   U15 : NAND2X1 port map( A => n176, B => n36, Y => n31);
   U16 : NAND2X1 port map( A => n37, B => n38, Y => nextstate_2_port);
   U17 : NOR2X1 port map( A => n39, B => n40, Y => n38);
   U18 : OAI21X1 port map( A => n25, B => n41, C => n34, Y => n40);
   U19 : OAI21X1 port map( A => n3, B => n42, C => n35, Y => n41);
   U20 : NAND2X1 port map( A => n177, B => n186, Y => n42);
   U21 : NAND2X1 port map( A => n45, B => n46, Y => n39);
   U22 : NOR2X1 port map( A => n47, B => n48, Y => n37);
   U23 : OAI22X1 port map( A => n23, B => n30, C => n50, D => n189, Y => n48);
   U24 : OAI21X1 port map( A => n35, B => n51, C => n52, Y => n47);
   U25 : OAI21X1 port map( A => n53, B => n54, C => n55, Y => n52);
   U26 : AOI22X1 port map( A => n56, B => n57, C => n36, D => n191, Y => n51);
   U27 : NOR2X1 port map( A => D_EDGE, B => n181, Y => n56);
   U28 : OAI21X1 port map( A => n168, B => n191, C => n59, Y => 
                           nextstate_1_port);
   U30 : OAI21X1 port map( A => n62, B => n63, C => n189, Y => n60);
   U31 : OAI21X1 port map( A => n29, B => n178, C => n65, Y => n63);
   U33 : OAI21X1 port map( A => n43, B => n67, C => n172, Y => n62);
   U34 : NAND2X1 port map( A => n179, B => n191, Y => n67);
   U35 : OAI22X1 port map( A => n70, B => n71, C => n30, D => n72, Y => 
                           nextstate_0_port);
   U36 : OAI21X1 port map( A => n181, B => n24, C => n74, Y => n72);
   U37 : NAND3X1 port map( A => n189, B => n181, C => n75, Y => n74);
   U38 : OAI21X1 port map( A => n19, B => n191, C => n77, Y => n75);
   U39 : AOI22X1 port map( A => n66, B => n78, C => n79, D => n80, Y => n77);
   U42 : OAI22X1 port map( A => state_0_port, B => n182, C => n81, D => n181, Y
                           => n71);
   U43 : AOI22X1 port map( A => EOP, B => n78, C => D_EDGE, D => n171, Y => n81
                           );
   U45 : OAI21X1 port map( A => state_2_port, B => n84, C => n85, Y => n70);
   U46 : NOR2X1 port map( A => n35, B => n36, Y => n85);
   U47 : AOI22X1 port map( A => n86, B => n66, C => D_EDGE, D => n78, Y => n84)
                           ;
   U48 : NOR2X1 port map( A => n179, B => EOP, Y => n66);
   U50 : NOR2X1 port map( A => BS_ERROR, B => n19, Y => n86);
   U52 : AOI21X1 port map( A => CRC_ERROR_port, B => RST, C => n88, Y => n87);
   U53 : OAI21X1 port map( A => n89, B => n90, C => n91, Y => n88);
   U54 : NAND2X1 port map( A => curCRC_ERROR, B => n92, Y => n90);
   U55 : NAND2X1 port map( A => n44, B => n30, Y => n89);
   U56 : OAI21X1 port map( A => n44, B => n188, C => n94, Y => n150);
   U57 : AOI21X1 port map( A => n9, B => n44, C => n170, Y => n94);
   U59 : NAND3X1 port map( A => n96, B => n30, C => curR_ERROR, Y => n95);
   U60 : OAI21X1 port map( A => n1, B => n181, C => n97, Y => n96);
   U61 : OAI21X1 port map( A => n176, B => n25, C => n98, Y => n9);
   U64 : OAI21X1 port map( A => n1, B => n80, C => n175, Y => n100);
   U65 : OAI21X1 port map( A => n54, B => n173, C => EOP, Y => n99);
   U69 : OAI21X1 port map( A => n103, B => n187, C => n91, Y => n151);
   U70 : NAND3X1 port map( A => n3, B => n44, C => n105, Y => n91);
   U71 : NOR2X1 port map( A => n25, B => n102, Y => n105);
   U72 : NAND3X1 port map( A => n35, B => n186, C => n177, Y => n102);
   U76 : AOI21X1 port map( A => n92, B => n30, C => RST, Y => n103);
   U77 : OAI21X1 port map( A => n181, B => n19, C => n97, Y => n92);
   U78 : NAND2X1 port map( A => n27, B => n83, Y => n97);
   U79 : NOR2X1 port map( A => D_EDGE, B => state_2_port, Y => n83);
   U81 : OAI21X1 port map( A => n107, B => n184, C => n109, Y => n161);
   U82 : NAND3X1 port map( A => n160, B => n184, C => count_0_port, Y => n109);
   U83 : AOI21X1 port map( A => n111, B => n180, C => n113, Y => n107);
   U84 : OAI21X1 port map( A => n157, B => n185, C => n116, Y => n162);
   U85 : NAND3X1 port map( A => n117, B => n185, C => n158, Y => n116);
   U87 : OAI21X1 port map( A => n120, B => n186, C => n121, Y => n163);
   U88 : NAND3X1 port map( A => n117, B => n186, C => n122, Y => n121);
   U89 : NOR2X1 port map( A => n123, B => n185, Y => n122);
   U90 : AOI21X1 port map( A => n111, B => n185, C => n119, Y => n120);
   U91 : OAI21X1 port map( A => n158, B => n166, C => n46, Y => n119);
   U93 : NAND3X1 port map( A => count_1_port, B => count_0_port, C => n125, Y 
                           => n123);
   U95 : AOI22X1 port map( A => n113, B => count_0_port, C => n180, D => n160, 
                           Y => n126);
   U97 : NAND3X1 port map( A => n117, B => n190, C => SHIFT_ENABLE, Y => n127);
   U100 : OAI21X1 port map( A => n125, B => n166, C => n46, Y => n113);
   U101 : NAND2X1 port map( A => EOP, B => n129, Y => n46);
   U103 : NOR2X1 port map( A => n55, B => n167, Y => n111);
   U104 : NOR2X1 port map( A => n186, B => n106, Y => n55);
   U105 : NAND3X1 port map( A => n184, B => n185, C => n180, Y => n106);
   U110 : NOR2X1 port map( A => BITSTUFF, B => n159, Y => n125);
   U115 : NAND3X1 port map( A => n134, B => n164, C => n79, Y => n33);
   U117 : NAND3X1 port map( A => n136, B => n137, C => n138, Y => n80);
   U119 : NOR2X1 port map( A => RCV_DATA(6), B => RCV_DATA(5), Y => n140);
   U120 : NOR2X1 port map( A => RCV_DATA(4), B => RCV_DATA(3), Y => n139);
   U121 : NOR2X1 port map( A => RCV_DATA(2), B => RCV_DATA(1), Y => n137);
   U122 : NOR2X1 port map( A => RCV_DATA(0), B => n165, Y => n136);
   U124 : NAND3X1 port map( A => n168, B => n61, C => n50, Y => RCVING);
   U125 : NOR2X1 port map( A => n129, B => n142, Y => n50);
   U126 : OAI21X1 port map( A => n183, B => n174, C => n133, Y => n142);
   U127 : NAND3X1 port map( A => state_2_port, B => n30, C => n27, Y => n133);
   U129 : OAI21X1 port map( A => n35, B => n25, C => n34, Y => n144);
   U130 : NAND3X1 port map( A => state_2_port, B => n30, C => n78, Y => n34);
   U133 : NAND3X1 port map( A => n43, B => n29, C => n172, Y => n129);
   U135 : NOR2X1 port map( A => n19, B => n183, Y => n53);
   U137 : NAND3X1 port map( A => n30, B => n181, C => n57, Y => n29);
   U141 : NOR2X1 port map( A => n30, B => state_2_port, Y => n134);
   U143 : NOR2X1 port map( A => n175, B => n171, Y => n78);
   U144 : OAI21X1 port map( A => n181, B => n23, C => n30, Y => n146);
   U148 : OAI21X1 port map( A => n147, B => n1, C => n35, Y => n145);
   U149 : NOR2X1 port map( A => state_0_port, B => n181, Y => n147);
   U150 : OAI21X1 port map( A => n30, B => n25, C => n61, Y => n192);
   U151 : NAND3X1 port map( A => n35, B => state_2_port, C => n57, Y => n61);
   U155 : NOR2X1 port map( A => n174, B => n181, Y => n36);
   U158 : NOR2X1 port map( A => state_0_port, B => n1, Y => n79);
   U3 : OR2X2 port map( A => n9, B => n170, Y => nxtR_ERROR);
   U4 : OR2X2 port map( A => n11, B => n12, Y => nextstate_3_port);
   U14 : AND2X2 port map( A => n33, B => n34, Y => n32);
   U29 : AND2X2 port map( A => n60, B => n61, Y => n59);
   U62 : AND2X2 port map( A => n99, B => n45, Y => n98);
   U63 : OR2X2 port map( A => n183, B => n100, Y => n45);
   U99 : AND2X2 port map( A => n111, B => n46, Y => n117);
   U114 : AND2X2 port map( A => n33, B => n133, Y => n65);
   U118 : AND2X2 port map( A => n139, B => n140, Y => n138);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => CLK, R => 
                           n44, S => n18, Q => state_1_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => CLK, R => 
                           n44, S => n17, Q => state_0_port);
   R_ERROR_reg : DFFSR port map( D => nxtR_ERROR, CLK => CLK, R => n44, S => 
                           n13, Q => R_ERROR);
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => CLK, R => 
                           n44, S => n10, Q => state_3_port);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => CLK, R => 
                           n44, S => n8, Q => state_2_port);
   count_reg_0_inst : DFFSR port map( D => n156, CLK => CLK, R => n44, S => n7,
                           Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => n161, CLK => CLK, R => n44, S => n6,
                           Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n162, CLK => CLK, R => n44, S => n5,
                           Q => count_2_port);
   count_reg_3_inst : DFFSR port map( D => n163, CLK => CLK, R => n44, S => n4,
                           Q => count_3_port);
   U10 : BUFX2 port map( A => state_3_port, Y => n1);
   U32 : INVX2 port map( A => state_0_port, Y => n175);
   U40 : AND2X2 port map( A => n146, B => n145, Y => n2);
   U41 : NAND2X1 port map( A => n152, B => n149, Y => n3);
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n10 <= '1';
   n13 <= '1';
   n17 <= '1';
   n18 <= '1';
   U75 : INVX2 port map( A => n1, Y => n171);
   U80 : OR2X2 port map( A => n175, B => n1, Y => n19);
   U86 : INVX2 port map( A => n19, Y => n57);
   U92 : OR2X2 port map( A => n171, B => state_0_port, Y => n23);
   U94 : INVX2 port map( A => n23, Y => n27);
   U96 : NAND2X1 port map( A => n167, B => n2, Y => OPCODE(1));
   U98 : OR2X2 port map( A => n175, B => n171, Y => n24);
   U102 : INVX2 port map( A => state_2_port, Y => n181);
   U106 : OR2X2 port map( A => n174, B => n181, Y => n25);
   U107 : OAI21X1 port map( A => n30, B => n25, C => n61, Y => OPCODE(0));
   U108 : INVX2 port map( A => n65, Y => n28);
   U109 : OR2X2 port map( A => n28, B => n192, Y => W_ENABLE);
   U111 : INVX2 port map( A => RST, Y => n44);
   U112 : INVX2 port map( A => n134, Y => n183);
   U113 : INVX2 port map( A => state_1_port, Y => n30);
   U116 : INVX1 port map( A => n30, Y => n35);
   U123 : OR2X2 port map( A => n24, B => n183, Y => n43);
   U128 : INVX1 port map( A => n43, Y => n54);
   U131 : XNOR2X1 port map( A => RX_CHECK_CRC(10), B => RX_CRC(10), Y => n69);
   U132 : XNOR2X1 port map( A => RX_CHECK_CRC(9), B => RX_CRC(9), Y => n68);
   U134 : XOR2X1 port map( A => RX_CHECK_CRC(7), B => RX_CRC(7), Y => n58);
   U136 : XOR2X1 port map( A => RX_CHECK_CRC(8), B => RX_CRC(8), Y => n49);
   U138 : NOR2X1 port map( A => n58, B => n49, Y => n64);
   U139 : NAND3X1 port map( A => n69, B => n68, C => n64, Y => n108);
   U140 : XNOR2X1 port map( A => RX_CHECK_CRC(14), B => RX_CRC(14), Y => n101);
   U142 : XNOR2X1 port map( A => RX_CHECK_CRC(13), B => RX_CRC(13), Y => n93);
   U145 : XOR2X1 port map( A => RX_CHECK_CRC(11), B => RX_CRC(11), Y => n76);
   U146 : XOR2X1 port map( A => RX_CHECK_CRC(12), B => RX_CRC(12), Y => n73);
   U147 : NOR2X1 port map( A => n76, B => n73, Y => n82);
   U152 : NAND3X1 port map( A => n101, B => n93, C => n82, Y => n104);
   U153 : NOR2X1 port map( A => n108, B => n104, Y => n152);
   U154 : NOR2X1 port map( A => n153, B => RX_CHECK_CRC(0), Y => n110);
   U156 : OAI22X1 port map( A => RX_CRC(1), B => n110, C => n110, D => n155, Y 
                           => n128);
   U157 : AND2X1 port map( A => RX_CHECK_CRC(0), B => n153, Y => n112);
   U159 : OAI22X1 port map( A => n112, B => n154, C => RX_CHECK_CRC(1), D => 
                           n112, Y => n124);
   U160 : XOR2X1 port map( A => RX_CHECK_CRC(15), B => RX_CRC(15), Y => n115);
   U161 : XOR2X1 port map( A => RX_CHECK_CRC(2), B => RX_CRC(2), Y => n114);
   U162 : NOR2X1 port map( A => n115, B => n114, Y => n118);
   U163 : NAND3X1 port map( A => n128, B => n124, C => n118, Y => n148);
   U164 : XNOR2X1 port map( A => RX_CHECK_CRC(6), B => RX_CRC(6), Y => n141);
   U165 : XNOR2X1 port map( A => RX_CHECK_CRC(5), B => RX_CRC(5), Y => n135);
   U166 : XOR2X1 port map( A => RX_CHECK_CRC(3), B => RX_CRC(3), Y => n131);
   U167 : XOR2X1 port map( A => RX_CHECK_CRC(4), B => RX_CRC(4), Y => n130);
   U168 : NOR2X1 port map( A => n131, B => n130, Y => n132);
   U169 : NAND3X1 port map( A => n141, B => n135, C => n132, Y => n143);
   U170 : NOR2X1 port map( A => n148, B => n143, Y => n149);
   U171 : INVX2 port map( A => RX_CRC(0), Y => n153);
   U172 : INVX2 port map( A => RX_CRC(1), Y => n154);
   U173 : INVX2 port map( A => RX_CHECK_CRC(1), Y => n155);
   U174 : INVX2 port map( A => n126, Y => n156);
   U175 : INVX2 port map( A => n119, Y => n157);
   U176 : INVX2 port map( A => n123, Y => n158);
   U177 : INVX2 port map( A => SHIFT_ENABLE, Y => n159);
   U178 : INVX2 port map( A => n127, Y => n160);
   U179 : INVX2 port map( A => n80, Y => n164);
   U180 : INVX2 port map( A => RCV_DATA(7), Y => n165);
   U181 : INVX2 port map( A => n111, Y => n166);
   U182 : INVX2 port map( A => n129, Y => n167);
   U183 : INVX2 port map( A => n144, Y => n168);
   U184 : INVX2 port map( A => n87, Y => n169);
   U185 : INVX2 port map( A => n95, Y => n170);
   U186 : INVX2 port map( A => n53, Y => n172);
   U187 : INVX2 port map( A => n29, Y => n173);
   U188 : INVX2 port map( A => n79, Y => n174);
   U189 : INVX2 port map( A => n102, Y => n176);
   U190 : INVX2 port map( A => n106, Y => n177);
   U191 : INVX2 port map( A => n66, Y => n178);
   U192 : INVX2 port map( A => n55, Y => n179);
   U193 : INVX2 port map( A => count_0_port, Y => n180);
   U194 : INVX2 port map( A => n83, Y => n182);
   U195 : INVX2 port map( A => count_1_port, Y => n184);
   U196 : INVX2 port map( A => count_2_port, Y => n185);
   U197 : INVX2 port map( A => count_3_port, Y => n186);
   U198 : INVX2 port map( A => curCRC_ERROR, Y => n187);
   U199 : INVX2 port map( A => curR_ERROR, Y => n188);
   U200 : INVX2 port map( A => BS_ERROR, Y => n189);
   U201 : INVX2 port map( A => BITSTUFF, Y => n190);
   U202 : INVX2 port map( A => EOP, Y => n191);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_eopdetect_1 is

   port( DP1_RX, DM1_RX : in std_logic;  EOP : out std_logic);

end rx_eopdetect_1;

architecture SYN_Behavioral of rx_eopdetect_1 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;

begin
   
   U1 : NOR2X1 port map( A => DP1_RX, B => DM1_RX, Y => EOP);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_edgedetect_1 is

   port( CLK, RST, DP1_RX : in std_logic;  D_EDGE : out std_logic);

end rx_edgedetect_1;

architecture SYN_Behavioral of rx_edgedetect_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal DP_hold1, DP_hold2, n1, n3, n4, n2 : std_logic;

begin
   
   DP_hold1_reg : DFFSR port map( D => DP1_RX, CLK => CLK, R => n3, S => n2, Q 
                           => DP_hold1);
   DP_hold2_reg : DFFSR port map( D => DP_hold1, CLK => CLK, R => n1, S => n2, 
                           Q => DP_hold2);
   n1 <= '1';
   n3 <= '1';
   U6 : NOR2X1 port map( A => RST, B => n4, Y => D_EDGE);
   U7 : XNOR2X1 port map( A => DP_hold2, B => DP_hold1, Y => n4);
   U4 : INVX2 port map( A => RST, Y => n2);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_decode_1 is

   port( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP : in std_logic;  D_ORIG, BITSTUFF,
         BS_ERROR : out std_logic);

end rx_decode_1;

architecture SYN_moore of rx_decode_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal DP_hold1, DP_hold2, state_3_port, state_2_port, state_1_port, 
      state_0_port, N29, N30, N31, N32, n1, n7, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29_port, n30_port, n31_port, n32_port, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, BITSTUFF_port, 
      n2, n3, n4, n5, n6, n8, n9, n10, BS_ERROR_port, n12, n13, n14, n15, n16 :
      std_logic;

begin
   BITSTUFF <= BITSTUFF_port;
   BS_ERROR <= BS_ERROR_port;
   
   DP_hold2_reg : DFFSR port map( D => n44, CLK => CLK, R => n7, S => n6, Q => 
                           DP_hold2);
   DP_hold1_reg : DFFSR port map( D => n43, CLK => CLK, R => n1, S => n6, Q => 
                           DP_hold1);
   n1 <= '1';
   n7 <= '1';
   U10 : OR2X2 port map( A => n8, B => state_1_port, Y => n36);
   U20 : NAND2X1 port map( A => n17, B => n18, Y => n43);
   U21 : AOI22X1 port map( A => DP_hold1, B => n12, C => DP1_RX, D => n19, Y =>
                           n17);
   U22 : NAND2X1 port map( A => n20, B => n18, Y => n44);
   U23 : AOI22X1 port map( A => n10, B => DP_hold1, C => DP_hold2, D => n21, Y 
                           => n20);
   U24 : NAND2X1 port map( A => SHIFT_ENABLE, B => n19, Y => n21);
   U25 : XNOR2X1 port map( A => DP_hold1, B => DP_hold2, Y => D_ORIG);
   U26 : NOR2X1 port map( A => n22, B => EOP, Y => N32);
   U27 : AOI21X1 port map( A => n23, B => BITSTUFF_port, C => BS_ERROR_port, Y 
                           => n22);
   U28 : NAND3X1 port map( A => state_3_port, B => n16, C => n25, Y => n24);
   U29 : NOR2X1 port map( A => state_2_port, B => state_1_port, Y => n25);
   U30 : NOR2X1 port map( A => n19, B => state_3_port, Y => BITSTUFF_port);
   U31 : NOR2X1 port map( A => n26, B => n14, Y => N31);
   U32 : AOI21X1 port map( A => state_2_port, B => n27, C => n28, Y => n26);
   U33 : OAI21X1 port map( A => n29_port, B => n30_port, C => n31_port, Y => 
                           n28);
   U34 : NAND2X1 port map( A => state_0_port, B => n23, Y => n30_port);
   U35 : NAND2X1 port map( A => state_1_port, B => n15, Y => n29_port);
   U36 : OAI21X1 port map( A => state_1_port, B => n32_port, C => SHIFT_ENABLE,
                           Y => n27);
   U37 : NOR2X1 port map( A => n33, B => n14, Y => N30);
   U38 : AOI21X1 port map( A => state_1_port, B => n34, C => n35, Y => n33);
   U39 : OAI21X1 port map( A => n16, B => n36, C => n31_port, Y => n35);
   U40 : NAND2X1 port map( A => n12, B => n32_port, Y => n31_port);
   U41 : NAND2X1 port map( A => n13, B => n16, Y => n19);
   U42 : OAI21X1 port map( A => n32_port, B => n37, C => SHIFT_ENABLE, Y => n34
                           );
   U43 : NAND2X1 port map( A => n16, B => n15, Y => n37);
   U44 : NOR2X1 port map( A => n38, B => n14, Y => N29);
   U45 : NOR2X1 port map( A => EOP, B => state_3_port, Y => n18);
   U46 : AOI21X1 port map( A => state_0_port, B => n9, C => n39, Y => n38);
   U47 : OAI21X1 port map( A => n8, B => n40, C => n41, Y => n39);
   U48 : NAND3X1 port map( A => n13, B => n32_port, C => SHIFT_ENABLE, Y => n41
                           );
   U49 : NAND2X1 port map( A => n42, B => n16, Y => n40);
   U50 : NAND2X1 port map( A => state_2_port, B => state_1_port, Y => n42);
   U51 : NOR2X1 port map( A => n32_port, B => n9, Y => n23);
   U52 : XOR2X1 port map( A => DP1_RX, B => DP_hold2, Y => n32_port);
   state_reg_3_inst : DFFSR port map( D => N32, CLK => CLK, R => n6, S => n5, Q
                           => state_3_port);
   state_reg_0_inst : DFFSR port map( D => N29, CLK => CLK, R => n6, S => n4, Q
                           => state_0_port);
   state_reg_2_inst : DFFSR port map( D => N31, CLK => CLK, R => n6, S => n3, Q
                           => state_2_port);
   state_reg_1_inst : DFFSR port map( D => N30, CLK => CLK, R => n6, S => n2, Q
                           => state_1_port);
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   n5 <= '1';
   U8 : INVX2 port map( A => RST, Y => n6);
   U11 : INVX2 port map( A => n23, Y => n8);
   U12 : INVX2 port map( A => SHIFT_ENABLE, Y => n9);
   U13 : INVX2 port map( A => n21, Y => n10);
   U14 : INVX2 port map( A => n24, Y => BS_ERROR_port);
   U15 : INVX2 port map( A => n19, Y => n12);
   U16 : INVX2 port map( A => n42, Y => n13);
   U17 : INVX2 port map( A => n18, Y => n14);
   U18 : INVX2 port map( A => state_2_port, Y => n15);
   U19 : INVX2 port map( A => state_0_port, Y => n16);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_accumulator_1 is

   port( CLK, RST : in std_logic;  RCV_DATA : in std_logic_vector (7 downto 0);
         W_ENABLE : in std_logic;  rx_CHECK_CRC : out std_logic_vector (15 
         downto 0));

end rx_accumulator_1;

architecture SYN_Behavioral of rx_accumulator_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, rx_CHECK_CRC_13_port, 
      rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, rx_CHECK_CRC_10_port, 
      rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, rx_CHECK_CRC_7_port, 
      rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, rx_CHECK_CRC_4_port, 
      rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, rx_CHECK_CRC_1_port, 
      rx_CHECK_CRC_0_port, n3, n4, n6, n7, n9, n10, n12, n13, n15, n16, n18, 
      n19, n21, n22, n24, n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n45
      , n47, n49, n51, n53, n55, n58, n1, n2, n5, n8, n11, n14, n17, n20, n23, 
      n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54
      , n56, n57, n59 : std_logic;

begin
   rx_CHECK_CRC <= ( rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, 
      rx_CHECK_CRC_13_port, rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, 
      rx_CHECK_CRC_10_port, rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, 
      rx_CHECK_CRC_7_port, rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, 
      rx_CHECK_CRC_4_port, rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, 
      rx_CHECK_CRC_1_port, rx_CHECK_CRC_0_port );
   
   U2 : OAI21X1 port map( A => n40, B => n59, C => n3, Y => n27);
   U3 : NAND2X1 port map( A => rx_CHECK_CRC_8_port, B => n40, Y => n3);
   U4 : OAI21X1 port map( A => n42, B => n59, C => n4, Y => n29);
   U5 : NAND2X1 port map( A => RCV_DATA(0), B => n42, Y => n4);
   U7 : OAI21X1 port map( A => n40, B => n57, C => n6, Y => n31);
   U8 : NAND2X1 port map( A => rx_CHECK_CRC_9_port, B => n40, Y => n6);
   U9 : OAI21X1 port map( A => n42, B => n57, C => n7, Y => n33);
   U10 : NAND2X1 port map( A => RCV_DATA(1), B => n42, Y => n7);
   U12 : OAI21X1 port map( A => n40, B => n56, C => n9, Y => n35);
   U13 : NAND2X1 port map( A => rx_CHECK_CRC_10_port, B => n40, Y => n9);
   U14 : OAI21X1 port map( A => n42, B => n56, C => n10, Y => n37);
   U15 : NAND2X1 port map( A => RCV_DATA(2), B => n42, Y => n10);
   U17 : OAI21X1 port map( A => n40, B => n54, C => n12, Y => n39);
   U18 : NAND2X1 port map( A => rx_CHECK_CRC_11_port, B => n40, Y => n12);
   U19 : OAI21X1 port map( A => n42, B => n54, C => n13, Y => n41);
   U20 : NAND2X1 port map( A => RCV_DATA(3), B => n42, Y => n13);
   U22 : OAI21X1 port map( A => n40, B => n52, C => n15, Y => n43);
   U23 : NAND2X1 port map( A => rx_CHECK_CRC_12_port, B => n40, Y => n15);
   U24 : OAI21X1 port map( A => n42, B => n52, C => n16, Y => n45);
   U25 : NAND2X1 port map( A => RCV_DATA(4), B => n42, Y => n16);
   U27 : OAI21X1 port map( A => n40, B => n50, C => n18, Y => n47);
   U28 : NAND2X1 port map( A => rx_CHECK_CRC_13_port, B => n40, Y => n18);
   U29 : OAI21X1 port map( A => n42, B => n50, C => n19, Y => n49);
   U30 : NAND2X1 port map( A => RCV_DATA(5), B => n42, Y => n19);
   U32 : OAI21X1 port map( A => n40, B => n48, C => n21, Y => n51);
   U33 : NAND2X1 port map( A => rx_CHECK_CRC_14_port, B => n40, Y => n21);
   U34 : OAI21X1 port map( A => n42, B => n48, C => n22, Y => n53);
   U35 : NAND2X1 port map( A => RCV_DATA(6), B => n42, Y => n22);
   U37 : OAI21X1 port map( A => n40, B => n46, C => n24, Y => n55);
   U38 : NAND2X1 port map( A => rx_CHECK_CRC_15_port, B => n40, Y => n24);
   U41 : OAI21X1 port map( A => n42, B => n46, C => n25, Y => n58);
   U42 : NAND2X1 port map( A => RCV_DATA(7), B => n42, Y => n25);
   present_CHECK_CRC_reg_7_inst : DFFSR port map( D => n58, CLK => CLK, R => 
                           n44, S => n38, Q => rx_CHECK_CRC_7_port);
   present_CHECK_CRC_reg_6_inst : DFFSR port map( D => n53, CLK => CLK, R => 
                           n44, S => n36, Q => rx_CHECK_CRC_6_port);
   present_CHECK_CRC_reg_5_inst : DFFSR port map( D => n49, CLK => CLK, R => 
                           n44, S => n34, Q => rx_CHECK_CRC_5_port);
   present_CHECK_CRC_reg_4_inst : DFFSR port map( D => n45, CLK => CLK, R => 
                           n44, S => n32, Q => rx_CHECK_CRC_4_port);
   present_CHECK_CRC_reg_3_inst : DFFSR port map( D => n41, CLK => CLK, R => 
                           n44, S => n30, Q => rx_CHECK_CRC_3_port);
   present_CHECK_CRC_reg_2_inst : DFFSR port map( D => n37, CLK => CLK, R => 
                           n44, S => n28, Q => rx_CHECK_CRC_2_port);
   present_CHECK_CRC_reg_1_inst : DFFSR port map( D => n33, CLK => CLK, R => 
                           n44, S => n26, Q => rx_CHECK_CRC_1_port);
   present_CHECK_CRC_reg_0_inst : DFFSR port map( D => n29, CLK => CLK, R => 
                           n44, S => n23, Q => rx_CHECK_CRC_0_port);
   present_CHECK_CRC_reg_15_inst : DFFSR port map( D => n55, CLK => CLK, R => 
                           n44, S => n20, Q => rx_CHECK_CRC_15_port);
   present_CHECK_CRC_reg_14_inst : DFFSR port map( D => n51, CLK => CLK, R => 
                           n44, S => n17, Q => rx_CHECK_CRC_14_port);
   present_CHECK_CRC_reg_13_inst : DFFSR port map( D => n47, CLK => CLK, R => 
                           n44, S => n14, Q => rx_CHECK_CRC_13_port);
   present_CHECK_CRC_reg_12_inst : DFFSR port map( D => n43, CLK => CLK, R => 
                           n44, S => n11, Q => rx_CHECK_CRC_12_port);
   present_CHECK_CRC_reg_11_inst : DFFSR port map( D => n39, CLK => CLK, R => 
                           n44, S => n8, Q => rx_CHECK_CRC_11_port);
   present_CHECK_CRC_reg_10_inst : DFFSR port map( D => n35, CLK => CLK, R => 
                           n44, S => n5, Q => rx_CHECK_CRC_10_port);
   present_CHECK_CRC_reg_9_inst : DFFSR port map( D => n31, CLK => CLK, R => 
                           n44, S => n2, Q => rx_CHECK_CRC_9_port);
   present_CHECK_CRC_reg_8_inst : DFFSR port map( D => n27, CLK => CLK, R => 
                           n44, S => n1, Q => rx_CHECK_CRC_8_port);
   U6 : INVX2 port map( A => W_ENABLE, Y => n40);
   n1 <= '1';
   n2 <= '1';
   n5 <= '1';
   n8 <= '1';
   n11 <= '1';
   n14 <= '1';
   n17 <= '1';
   n20 <= '1';
   n23 <= '1';
   n26 <= '1';
   n28 <= '1';
   n30 <= '1';
   n32 <= '1';
   n34 <= '1';
   n36 <= '1';
   n38 <= '1';
   U51 : INVX2 port map( A => n40, Y => n42);
   U52 : INVX2 port map( A => RST, Y => n44);
   U53 : INVX2 port map( A => rx_CHECK_CRC_7_port, Y => n46);
   U54 : INVX2 port map( A => rx_CHECK_CRC_6_port, Y => n48);
   U55 : INVX2 port map( A => rx_CHECK_CRC_5_port, Y => n50);
   U56 : INVX2 port map( A => rx_CHECK_CRC_4_port, Y => n52);
   U57 : INVX2 port map( A => rx_CHECK_CRC_3_port, Y => n54);
   U58 : INVX2 port map( A => rx_CHECK_CRC_2_port, Y => n56);
   U59 : INVX2 port map( A => rx_CHECK_CRC_1_port, Y => n57);
   U60 : INVX2 port map( A => rx_CHECK_CRC_0_port, Y => n59);

end SYN_Behavioral;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rx_CRC_CALC_1 is

   port( CLK, RST, W_ENABLE : in std_logic;  OPCODE : in std_logic_vector (1 
         downto 0);  RCV_DATA : in std_logic_vector (7 downto 0);  RX_CRC : out
         std_logic_vector (15 downto 0));

end rx_CRC_CALC_1;

architecture SYN_moore of rx_CRC_CALC_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port, current_crc_15_port, 
      current_crc_14_port, current_crc_13_port, current_crc_12_port, 
      current_crc_11_port, current_crc_10_port, current_crc_9_port, 
      current_crc_8_port, current_crc_7_port, current_crc_6_port, 
      current_crc_5_port, current_crc_4_port, current_crc_3_port, 
      current_crc_2_port, current_crc_1_port, current_crc_0_port, 
      cache_1_15_port, cache_1_14_port, cache_1_13_port, cache_1_12_port, 
      cache_1_11_port, cache_1_10_port, cache_1_9_port, cache_1_8_port, 
      cache_1_7_port, cache_1_6_port, cache_1_5_port, cache_1_4_port, 
      cache_1_3_port, cache_1_2_port, cache_1_1_port, cache_1_0_port, n3, n5, 
      n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, n33, n51, 
      n52, n53, n54, n55, n57, n58, n59, n61, n62, n63, n64, n65, n66, n67, n68
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n101, 
      n103, n105, n107, n109, n111, n113, n115, n117, n119, n121, n123, n125, 
      n127, n129, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n1, n2, n4, n6, n8, n10, n12, n14, 
      n16, n18, n20, n22, n24, n26, n28, n30, n32, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n56, n60, n79, 
      n80, n81, n82, n100, n102, n104, n106, n108, n110, n112, n114, n116, n118
      , n120, n122, n124, n126, n128, n130, n131, n148, n149, n150, n151, n152,
      n153, n154, n155, n156 : std_logic;

begin
   RX_CRC <= ( RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, RX_CRC_12_port, 
      RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, RX_CRC_8_port, 
      RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port, RX_CRC_3_port
      , RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port );
   
   cache_1_reg_0_inst : DFFPOSX1 port map( D => n129, CLK => CLK, Q => 
                           cache_1_0_port);
   cache_1_reg_8_inst : DFFPOSX1 port map( D => n127, CLK => CLK, Q => 
                           cache_1_8_port);
   cache_1_reg_15_inst : DFFPOSX1 port map( D => n125, CLK => CLK, Q => 
                           cache_1_15_port);
   cache_1_reg_1_inst : DFFPOSX1 port map( D => n123, CLK => CLK, Q => 
                           cache_1_1_port);
   cache_1_reg_9_inst : DFFPOSX1 port map( D => n121, CLK => CLK, Q => 
                           cache_1_9_port);
   cache_1_reg_2_inst : DFFPOSX1 port map( D => n119, CLK => CLK, Q => 
                           cache_1_2_port);
   cache_1_reg_10_inst : DFFPOSX1 port map( D => n117, CLK => CLK, Q => 
                           cache_1_10_port);
   cache_1_reg_3_inst : DFFPOSX1 port map( D => n115, CLK => CLK, Q => 
                           cache_1_3_port);
   cache_1_reg_11_inst : DFFPOSX1 port map( D => n113, CLK => CLK, Q => 
                           cache_1_11_port);
   cache_1_reg_4_inst : DFFPOSX1 port map( D => n111, CLK => CLK, Q => 
                           cache_1_4_port);
   cache_1_reg_12_inst : DFFPOSX1 port map( D => n109, CLK => CLK, Q => 
                           cache_1_12_port);
   cache_1_reg_5_inst : DFFPOSX1 port map( D => n107, CLK => CLK, Q => 
                           cache_1_5_port);
   cache_1_reg_13_inst : DFFPOSX1 port map( D => n105, CLK => CLK, Q => 
                           cache_1_13_port);
   cache_1_reg_6_inst : DFFPOSX1 port map( D => n103, CLK => CLK, Q => 
                           cache_1_6_port);
   cache_1_reg_14_inst : DFFPOSX1 port map( D => n101, CLK => CLK, Q => 
                           cache_1_14_port);
   cache_1_reg_7_inst : DFFPOSX1 port map( D => n99, CLK => CLK, Q => 
                           cache_1_7_port);
   cache_2_reg_15_inst : DFFPOSX1 port map( D => n98, CLK => CLK, Q => 
                           RX_CRC_15_port);
   cache_2_reg_14_inst : DFFPOSX1 port map( D => n97, CLK => CLK, Q => 
                           RX_CRC_14_port);
   cache_2_reg_13_inst : DFFPOSX1 port map( D => n96, CLK => CLK, Q => 
                           RX_CRC_13_port);
   cache_2_reg_12_inst : DFFPOSX1 port map( D => n95, CLK => CLK, Q => 
                           RX_CRC_12_port);
   cache_2_reg_11_inst : DFFPOSX1 port map( D => n94, CLK => CLK, Q => 
                           RX_CRC_11_port);
   cache_2_reg_10_inst : DFFPOSX1 port map( D => n93, CLK => CLK, Q => 
                           RX_CRC_10_port);
   cache_2_reg_9_inst : DFFPOSX1 port map( D => n92, CLK => CLK, Q => 
                           RX_CRC_9_port);
   cache_2_reg_8_inst : DFFPOSX1 port map( D => n91, CLK => CLK, Q => 
                           RX_CRC_8_port);
   cache_2_reg_7_inst : DFFPOSX1 port map( D => n90, CLK => CLK, Q => 
                           RX_CRC_7_port);
   cache_2_reg_6_inst : DFFPOSX1 port map( D => n89, CLK => CLK, Q => 
                           RX_CRC_6_port);
   cache_2_reg_5_inst : DFFPOSX1 port map( D => n88, CLK => CLK, Q => 
                           RX_CRC_5_port);
   cache_2_reg_4_inst : DFFPOSX1 port map( D => n87, CLK => CLK, Q => 
                           RX_CRC_4_port);
   cache_2_reg_3_inst : DFFPOSX1 port map( D => n86, CLK => CLK, Q => 
                           RX_CRC_3_port);
   cache_2_reg_2_inst : DFFPOSX1 port map( D => n85, CLK => CLK, Q => 
                           RX_CRC_2_port);
   cache_2_reg_1_inst : DFFPOSX1 port map( D => n84, CLK => CLK, Q => 
                           RX_CRC_1_port);
   cache_2_reg_0_inst : DFFPOSX1 port map( D => n83, CLK => CLK, Q => 
                           RX_CRC_0_port);
   U3 : OAI21X1 port map( A => n42, B => n60, C => n3, Y => n83);
   U4 : NAND2X1 port map( A => RX_CRC_0_port, B => n43, Y => n3);
   U5 : OAI21X1 port map( A => n41, B => n102, C => n5, Y => n84);
   U6 : NAND2X1 port map( A => RX_CRC_1_port, B => n43, Y => n5);
   U7 : OAI21X1 port map( A => n41, B => n110, C => n7, Y => n85);
   U8 : NAND2X1 port map( A => RX_CRC_2_port, B => n43, Y => n7);
   U9 : OAI21X1 port map( A => n41, B => n118, C => n9, Y => n86);
   U10 : NAND2X1 port map( A => RX_CRC_3_port, B => n43, Y => n9);
   U11 : OAI21X1 port map( A => n41, B => n126, C => n11, Y => n87);
   U12 : NAND2X1 port map( A => RX_CRC_4_port, B => n43, Y => n11);
   U13 : OAI21X1 port map( A => n41, B => n148, C => n13, Y => n88);
   U14 : NAND2X1 port map( A => RX_CRC_5_port, B => n42, Y => n13);
   U15 : OAI21X1 port map( A => n41, B => n152, C => n15, Y => n89);
   U16 : NAND2X1 port map( A => RX_CRC_6_port, B => n42, Y => n15);
   U17 : OAI21X1 port map( A => n41, B => n156, C => n17, Y => n90);
   U18 : NAND2X1 port map( A => RX_CRC_7_port, B => n42, Y => n17);
   U19 : OAI21X1 port map( A => n41, B => n80, C => n19, Y => n91);
   U20 : NAND2X1 port map( A => RX_CRC_8_port, B => n42, Y => n19);
   U21 : OAI21X1 port map( A => n41, B => n106, C => n21, Y => n92);
   U22 : NAND2X1 port map( A => RX_CRC_9_port, B => n42, Y => n21);
   U23 : OAI21X1 port map( A => n42, B => n114, C => n23, Y => n93);
   U24 : NAND2X1 port map( A => RX_CRC_10_port, B => n42, Y => n23);
   U25 : OAI21X1 port map( A => n42, B => n122, C => n25, Y => n94);
   U26 : NAND2X1 port map( A => RX_CRC_11_port, B => n42, Y => n25);
   U27 : OAI21X1 port map( A => n42, B => n130, C => n27, Y => n95);
   U28 : NAND2X1 port map( A => RX_CRC_12_port, B => n42, Y => n27);
   U29 : OAI21X1 port map( A => n42, B => n150, C => n29, Y => n96);
   U30 : NAND2X1 port map( A => RX_CRC_13_port, B => n43, Y => n29);
   U31 : OAI21X1 port map( A => n42, B => n154, C => n31, Y => n97);
   U32 : NAND2X1 port map( A => RX_CRC_14_port, B => n43, Y => n31);
   U33 : OAI21X1 port map( A => n42, B => n82, C => n33, Y => n98);
   U34 : NAND2X1 port map( A => RX_CRC_15_port, B => n43, Y => n33);
   U35 : OAI22X1 port map( A => n41, B => n155, C => n39, D => n156, Y => n99);
   U37 : OAI22X1 port map( A => n41, B => n153, C => n39, D => n154, Y => n101)
                           ;
   U39 : OAI22X1 port map( A => n41, B => n151, C => n39, D => n152, Y => n103)
                           ;
   U41 : OAI22X1 port map( A => n41, B => n149, C => n39, D => n150, Y => n105)
                           ;
   U43 : OAI22X1 port map( A => n40, B => n131, C => n39, D => n148, Y => n107)
                           ;
   U45 : OAI22X1 port map( A => n40, B => n128, C => n39, D => n130, Y => n109)
                           ;
   U47 : OAI22X1 port map( A => n40, B => n124, C => n39, D => n126, Y => n111)
                           ;
   U49 : OAI22X1 port map( A => n40, B => n120, C => n39, D => n122, Y => n113)
                           ;
   U51 : OAI22X1 port map( A => n40, B => n116, C => n39, D => n118, Y => n115)
                           ;
   U53 : OAI22X1 port map( A => n40, B => n112, C => n38, D => n114, Y => n117)
                           ;
   U55 : OAI22X1 port map( A => n40, B => n108, C => n38, D => n110, Y => n119)
                           ;
   U57 : OAI22X1 port map( A => n40, B => n104, C => n38, D => n106, Y => n121)
                           ;
   U59 : OAI22X1 port map( A => n40, B => n100, C => n38, D => n102, Y => n123)
                           ;
   U61 : OAI22X1 port map( A => n40, B => n81, C => n38, D => n82, Y => n125);
   U63 : OAI22X1 port map( A => n40, B => n79, C => n38, D => n80, Y => n127);
   U65 : OAI22X1 port map( A => n40, B => n56, C => n38, D => n60, Y => n129);
   U70 : OAI22X1 port map( A => n81, B => n37, C => n53, D => n35, Y => n132);
   U71 : XOR2X1 port map( A => n54, B => current_crc_7_port, Y => n53);
   U72 : OAI22X1 port map( A => n35, B => n151, C => n153, D => n37, Y => n133)
                           ;
   U73 : OAI22X1 port map( A => n35, B => n131, C => n149, D => n52, Y => n134)
                           ;
   U74 : OAI22X1 port map( A => n51, B => n124, C => n128, D => n37, Y => n135)
                           ;
   U75 : OAI22X1 port map( A => n35, B => n116, C => n120, D => n52, Y => n136)
                           ;
   U77 : OAI22X1 port map( A => n51, B => n108, C => n112, D => n37, Y => n137)
                           ;
   U78 : OAI22X1 port map( A => n104, B => n37, C => n55, D => n51, Y => n138);
   U79 : XOR2X1 port map( A => n100, B => n45, Y => n55);
   U80 : OAI22X1 port map( A => n79, B => n52, C => n57, D => n35, Y => n139);
   U81 : XOR2X1 port map( A => n58, B => n59, Y => n57);
   U82 : XOR2X1 port map( A => n56, B => n45, Y => n58);
   U84 : OAI22X1 port map( A => n155, B => n37, C => n46, D => n51, Y => n140);
   U86 : OAI22X1 port map( A => n151, B => n52, C => n61, D => n35, Y => n141);
   U87 : XOR2X1 port map( A => n62, B => n63, Y => n61);
   U89 : OAI22X1 port map( A => n131, B => n37, C => n64, D => n51, Y => n142);
   U91 : OAI22X1 port map( A => n124, B => n52, C => n65, D => n35, Y => n143);
   U92 : XOR2X1 port map( A => n66, B => n67, Y => n65);
   U94 : OAI22X1 port map( A => n116, B => n37, C => n68, D => n51, Y => n144);
   U96 : OAI22X1 port map( A => n108, B => n52, C => n69, D => n35, Y => n145);
   U97 : XOR2X1 port map( A => n70, B => n71, Y => n69);
   U99 : OAI22X1 port map( A => n100, B => n37, C => n72, D => n51, Y => n146);
   U100 : XOR2X1 port map( A => n73, B => n74, Y => n72);
   U101 : XOR2X1 port map( A => n75, B => n76, Y => n73);
   U103 : OAI22X1 port map( A => n56, B => n52, C => n54, D => n35, Y => n147);
   U104 : XOR2X1 port map( A => n77, B => n78, Y => n54);
   U105 : XOR2X1 port map( A => n45, B => n71, Y => n78);
   U106 : XOR2X1 port map( A => current_crc_8_port, B => RCV_DATA(0), Y => n71)
                           ;
   U108 : XOR2X1 port map( A => n81, B => RCV_DATA(7), Y => n75);
   U110 : XOR2X1 port map( A => n46, B => n76, Y => n77);
   U111 : XOR2X1 port map( A => n68, B => n64, Y => n76);
   U112 : XNOR2X1 port map( A => n63, B => n67, Y => n64);
   U113 : XOR2X1 port map( A => current_crc_11_port, B => RCV_DATA(3), Y => n67
                           );
   U114 : XNOR2X1 port map( A => n128, B => RCV_DATA(4), Y => n63);
   U116 : XOR2X1 port map( A => n70, B => n48, Y => n68);
   U118 : XOR2X1 port map( A => n112, B => RCV_DATA(2), Y => n66);
   U120 : XOR2X1 port map( A => n104, B => RCV_DATA(1), Y => n70);
   U123 : XOR2X1 port map( A => n59, B => n47, Y => n74);
   U125 : XOR2X1 port map( A => n149, B => RCV_DATA(5), Y => n62);
   U127 : XNOR2X1 port map( A => n153, B => RCV_DATA(6), Y => n59);
   U129 : OAI21X1 port map( A => n50, B => n49, C => n51, Y => n52);
   U130 : NAND3X1 port map( A => OPCODE(0), B => n49, C => W_ENABLE, Y => n51);
   current_crc_reg_14_inst : DFFSR port map( D => n133, CLK => CLK, R => n44, S
                           => n30, Q => current_crc_14_port);
   current_crc_reg_12_inst : DFFSR port map( D => n135, CLK => CLK, R => n44, S
                           => n28, Q => current_crc_12_port);
   current_crc_reg_10_inst : DFFSR port map( D => n137, CLK => CLK, R => n44, S
                           => n26, Q => current_crc_10_port);
   current_crc_reg_13_inst : DFFSR port map( D => n134, CLK => CLK, R => n44, S
                           => n24, Q => current_crc_13_port);
   current_crc_reg_11_inst : DFFSR port map( D => n136, CLK => CLK, R => n44, S
                           => n22, Q => current_crc_11_port);
   current_crc_reg_15_inst : DFFSR port map( D => n132, CLK => CLK, R => n44, S
                           => n20, Q => current_crc_15_port);
   current_crc_reg_8_inst : DFFSR port map( D => n139, CLK => CLK, R => n44, S 
                           => n18, Q => current_crc_8_port);
   current_crc_reg_6_inst : DFFSR port map( D => n141, CLK => CLK, R => n44, S 
                           => n16, Q => current_crc_6_port);
   current_crc_reg_4_inst : DFFSR port map( D => n143, CLK => CLK, R => n44, S 
                           => n14, Q => current_crc_4_port);
   current_crc_reg_2_inst : DFFSR port map( D => n145, CLK => CLK, R => n44, S 
                           => n12, Q => current_crc_2_port);
   current_crc_reg_0_inst : DFFSR port map( D => n147, CLK => CLK, R => n44, S 
                           => n10, Q => current_crc_0_port);
   current_crc_reg_9_inst : DFFSR port map( D => n138, CLK => CLK, R => n44, S 
                           => n8, Q => current_crc_9_port);
   current_crc_reg_7_inst : DFFSR port map( D => n140, CLK => CLK, R => n44, S 
                           => n6, Q => current_crc_7_port);
   current_crc_reg_5_inst : DFFSR port map( D => n142, CLK => CLK, R => n44, S 
                           => n4, Q => current_crc_5_port);
   current_crc_reg_3_inst : DFFSR port map( D => n144, CLK => CLK, R => n44, S 
                           => n2, Q => current_crc_3_port);
   current_crc_reg_1_inst : DFFSR port map( D => n146, CLK => CLK, R => n44, S 
                           => n1, Q => current_crc_1_port);
   U36 : INVX2 port map( A => OPCODE(1), Y => n49);
   U38 : INVX2 port map( A => n32, Y => n38);
   n1 <= '1';
   n2 <= '1';
   n4 <= '1';
   n6 <= '1';
   n8 <= '1';
   n10 <= '1';
   n12 <= '1';
   n14 <= '1';
   n16 <= '1';
   n18 <= '1';
   n20 <= '1';
   n22 <= '1';
   n24 <= '1';
   n26 <= '1';
   n28 <= '1';
   n30 <= '1';
   U69 : INVX2 port map( A => n51, Y => n34);
   U76 : BUFX2 port map( A => n32, Y => n40);
   U83 : BUFX2 port map( A => n32, Y => n43);
   U85 : INVX2 port map( A => n32, Y => n39);
   U88 : OR2X2 port map( A => n35, B => RST, Y => n32);
   U90 : INVX2 port map( A => n34, Y => n35);
   U93 : INVX2 port map( A => n36, Y => n37);
   U95 : INVX2 port map( A => n52, Y => n36);
   U98 : INVX2 port map( A => RST, Y => n44);
   U102 : INVX1 port map( A => OPCODE(0), Y => n50);
   U107 : BUFX4 port map( A => n32, Y => n41);
   U109 : BUFX4 port map( A => n32, Y => n42);
   U115 : INVX2 port map( A => n75, Y => n45);
   U117 : INVX2 port map( A => n74, Y => n46);
   U119 : INVX2 port map( A => n62, Y => n47);
   U121 : INVX2 port map( A => n66, Y => n48);
   U122 : INVX2 port map( A => current_crc_0_port, Y => n56);
   U124 : INVX2 port map( A => cache_1_0_port, Y => n60);
   U126 : INVX2 port map( A => current_crc_8_port, Y => n79);
   U128 : INVX2 port map( A => cache_1_8_port, Y => n80);
   U131 : INVX2 port map( A => current_crc_15_port, Y => n81);
   U132 : INVX2 port map( A => cache_1_15_port, Y => n82);
   U133 : INVX2 port map( A => current_crc_1_port, Y => n100);
   U134 : INVX2 port map( A => cache_1_1_port, Y => n102);
   U135 : INVX2 port map( A => current_crc_9_port, Y => n104);
   U136 : INVX2 port map( A => cache_1_9_port, Y => n106);
   U137 : INVX2 port map( A => current_crc_2_port, Y => n108);
   U138 : INVX2 port map( A => cache_1_2_port, Y => n110);
   U139 : INVX2 port map( A => current_crc_10_port, Y => n112);
   U140 : INVX2 port map( A => cache_1_10_port, Y => n114);
   U141 : INVX2 port map( A => current_crc_3_port, Y => n116);
   U142 : INVX2 port map( A => cache_1_3_port, Y => n118);
   U143 : INVX2 port map( A => current_crc_11_port, Y => n120);
   U144 : INVX2 port map( A => cache_1_11_port, Y => n122);
   U145 : INVX2 port map( A => current_crc_4_port, Y => n124);
   U146 : INVX2 port map( A => cache_1_4_port, Y => n126);
   U147 : INVX2 port map( A => current_crc_12_port, Y => n128);
   U148 : INVX2 port map( A => cache_1_12_port, Y => n130);
   U149 : INVX2 port map( A => current_crc_5_port, Y => n131);
   U150 : INVX2 port map( A => cache_1_5_port, Y => n148);
   U151 : INVX2 port map( A => current_crc_13_port, Y => n149);
   U152 : INVX2 port map( A => cache_1_13_port, Y => n150);
   U153 : INVX2 port map( A => current_crc_6_port, Y => n151);
   U154 : INVX2 port map( A => cache_1_6_port, Y => n152);
   U155 : INVX2 port map( A => current_crc_14_port, Y => n153);
   U156 : INVX2 port map( A => cache_1_14_port, Y => n154);
   U157 : INVX2 port map( A => current_crc_7_port, Y => n155);
   U158 : INVX2 port map( A => cache_1_7_port, Y => n156);

end SYN_moore;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RFIFO_1 is

   port( CLK, RST, W_ENABLE, R_ENABLE : in std_logic;  RCV_DATA : in 
         std_logic_vector (7 downto 0);  RCV_OPCODE : in std_logic_vector (1 
         downto 0);  DATA : out std_logic_vector (7 downto 0);  OUT_OPCODE : 
         out std_logic_vector (1 downto 0);  BYTE_COUNT : out std_logic_vector 
         (4 downto 0);  EMPTY, FULL : out std_logic);

end RFIFO_1;

architecture SYN_BRFIFO of RFIFO_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, 
      DATA_3_port, DATA_2_port, DATA_1_port, DATA_0_port, OUT_OPCODE_1_port, 
      OUT_OPCODE_0_port, EMPTY_port, FULL_port, readptr_4_port, readptr_3_port,
      readptr_2_port, readptr_1_port, readptr_0_port, writeptr_4_port, 
      writeptr_3_port, writeptr_2_port, writeptr_1_port, writeptr_0_port, state
      , N32, N33, N34, N43, N44, N45, N46, opcode_0_1_port, opcode_0_0_port, 
      opcode_1_1_port, opcode_1_0_port, opcode_2_1_port, opcode_2_0_port, 
      opcode_3_1_port, opcode_3_0_port, opcode_4_1_port, opcode_4_0_port, 
      opcode_5_1_port, opcode_5_0_port, opcode_6_1_port, opcode_6_0_port, 
      opcode_7_1_port, opcode_7_0_port, opcode_8_1_port, opcode_8_0_port, 
      opcode_9_1_port, opcode_9_0_port, opcode_10_1_port, opcode_10_0_port, 
      opcode_11_1_port, opcode_11_0_port, opcode_12_1_port, opcode_12_0_port, 
      opcode_13_1_port, opcode_13_0_port, opcode_14_1_port, opcode_14_0_port, 
      opcode_15_1_port, opcode_15_0_port, opcode_16_1_port, opcode_16_0_port, 
      opcode_17_1_port, opcode_17_0_port, opcode_18_1_port, opcode_18_0_port, 
      opcode_19_1_port, opcode_19_0_port, opcode_20_1_port, opcode_20_0_port, 
      opcode_21_1_port, opcode_21_0_port, opcode_22_1_port, opcode_22_0_port, 
      opcode_23_1_port, opcode_23_0_port, opcode_24_1_port, opcode_24_0_port, 
      opcode_25_1_port, opcode_25_0_port, opcode_26_1_port, opcode_26_0_port, 
      opcode_27_1_port, opcode_27_0_port, opcode_28_1_port, opcode_28_0_port, 
      opcode_29_1_port, opcode_29_0_port, opcode_30_1_port, opcode_30_0_port, 
      opcode_31_1_port, opcode_31_0_port, memory_0_7_port, memory_0_6_port, 
      memory_0_5_port, memory_0_4_port, memory_0_3_port, memory_0_2_port, 
      memory_0_1_port, memory_0_0_port, memory_1_7_port, memory_1_6_port, 
      memory_1_5_port, memory_1_4_port, memory_1_3_port, memory_1_2_port, 
      memory_1_1_port, memory_1_0_port, memory_2_7_port, memory_2_6_port, 
      memory_2_5_port, memory_2_4_port, memory_2_3_port, memory_2_2_port, 
      memory_2_1_port, memory_2_0_port, memory_3_7_port, memory_3_6_port, 
      memory_3_5_port, memory_3_4_port, memory_3_3_port, memory_3_2_port, 
      memory_3_1_port, memory_3_0_port, memory_4_7_port, memory_4_6_port, 
      memory_4_5_port, memory_4_4_port, memory_4_3_port, memory_4_2_port, 
      memory_4_1_port, memory_4_0_port, memory_5_7_port, memory_5_6_port, 
      memory_5_5_port, memory_5_4_port, memory_5_3_port, memory_5_2_port, 
      memory_5_1_port, memory_5_0_port, memory_6_7_port, memory_6_6_port, 
      memory_6_5_port, memory_6_4_port, memory_6_3_port, memory_6_2_port, 
      memory_6_1_port, memory_6_0_port, memory_7_7_port, memory_7_6_port, 
      memory_7_5_port, memory_7_4_port, memory_7_3_port, memory_7_2_port, 
      memory_7_1_port, memory_7_0_port, memory_8_7_port, memory_8_6_port, 
      memory_8_5_port, memory_8_4_port, memory_8_3_port, memory_8_2_port, 
      memory_8_1_port, memory_8_0_port, memory_9_7_port, memory_9_6_port, 
      memory_9_5_port, memory_9_4_port, memory_9_3_port, memory_9_2_port, 
      memory_9_1_port, memory_9_0_port, memory_10_7_port, memory_10_6_port, 
      memory_10_5_port, memory_10_4_port, memory_10_3_port, memory_10_2_port, 
      memory_10_1_port, memory_10_0_port, memory_11_7_port, memory_11_6_port, 
      memory_11_5_port, memory_11_4_port, memory_11_3_port, memory_11_2_port, 
      memory_11_1_port, memory_11_0_port, memory_12_7_port, memory_12_6_port, 
      memory_12_5_port, memory_12_4_port, memory_12_3_port, memory_12_2_port, 
      memory_12_1_port, memory_12_0_port, memory_13_7_port, memory_13_6_port, 
      memory_13_5_port, memory_13_4_port, memory_13_3_port, memory_13_2_port, 
      memory_13_1_port, memory_13_0_port, memory_14_7_port, memory_14_6_port, 
      memory_14_5_port, memory_14_4_port, memory_14_3_port, memory_14_2_port, 
      memory_14_1_port, memory_14_0_port, memory_15_7_port, memory_15_6_port, 
      memory_15_5_port, memory_15_4_port, memory_15_3_port, memory_15_2_port, 
      memory_15_1_port, memory_15_0_port, memory_16_7_port, memory_16_6_port, 
      memory_16_5_port, memory_16_4_port, memory_16_3_port, memory_16_2_port, 
      memory_16_1_port, memory_16_0_port, memory_17_7_port, memory_17_6_port, 
      memory_17_5_port, memory_17_4_port, memory_17_3_port, memory_17_2_port, 
      memory_17_1_port, memory_17_0_port, memory_18_7_port, memory_18_6_port, 
      memory_18_5_port, memory_18_4_port, memory_18_3_port, memory_18_2_port, 
      memory_18_1_port, memory_18_0_port, memory_19_7_port, memory_19_6_port, 
      memory_19_5_port, memory_19_4_port, memory_19_3_port, memory_19_2_port, 
      memory_19_1_port, memory_19_0_port, memory_20_7_port, memory_20_6_port, 
      memory_20_5_port, memory_20_4_port, memory_20_3_port, memory_20_2_port, 
      memory_20_1_port, memory_20_0_port, memory_21_7_port, memory_21_6_port, 
      memory_21_5_port, memory_21_4_port, memory_21_3_port, memory_21_2_port, 
      memory_21_1_port, memory_21_0_port, memory_22_7_port, memory_22_6_port, 
      memory_22_5_port, memory_22_4_port, memory_22_3_port, memory_22_2_port, 
      memory_22_1_port, memory_22_0_port, memory_23_7_port, memory_23_6_port, 
      memory_23_5_port, memory_23_4_port, memory_23_3_port, memory_23_2_port, 
      memory_23_1_port, memory_23_0_port, memory_24_7_port, memory_24_6_port, 
      memory_24_5_port, memory_24_4_port, memory_24_3_port, memory_24_2_port, 
      memory_24_1_port, memory_24_0_port, memory_25_7_port, memory_25_6_port, 
      memory_25_5_port, memory_25_4_port, memory_25_3_port, memory_25_2_port, 
      memory_25_1_port, memory_25_0_port, memory_26_7_port, memory_26_6_port, 
      memory_26_5_port, memory_26_4_port, memory_26_3_port, memory_26_2_port, 
      memory_26_1_port, memory_26_0_port, memory_27_7_port, memory_27_6_port, 
      memory_27_5_port, memory_27_4_port, memory_27_3_port, memory_27_2_port, 
      memory_27_1_port, memory_27_0_port, memory_28_7_port, memory_28_6_port, 
      memory_28_5_port, memory_28_4_port, memory_28_3_port, memory_28_2_port, 
      memory_28_1_port, memory_28_0_port, memory_29_7_port, memory_29_6_port, 
      memory_29_5_port, memory_29_4_port, memory_29_3_port, memory_29_2_port, 
      memory_29_1_port, memory_29_0_port, memory_30_7_port, memory_30_6_port, 
      memory_30_5_port, memory_30_4_port, memory_30_3_port, memory_30_2_port, 
      memory_30_1_port, memory_30_0_port, memory_31_7_port, memory_31_6_port, 
      memory_31_5_port, memory_31_4_port, memory_31_3_port, memory_31_2_port, 
      memory_31_1_port, memory_31_0_port, N48, N49, N50, N51, N189, N190, N191,
      N192, N193, N195, N333, N334, N335, N336, N337, N338, N339, N340, N341, 
      N342, N343, N344, N345, N346, N347, n854, n856, n858, n860, n862, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1072, n1073, n1074, 
      n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
      n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
      n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, 
      n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
      n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
      n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
      n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
      n1165, n1166, n1167, add_76_aco_carry_1_port, add_76_aco_carry_2_port, 
      add_76_aco_carry_3_port, add_76_aco_carry_4_port, sub_72_carry_1_port, 
      sub_72_carry_2_port, sub_72_carry_3_port, sub_72_carry_4_port, 
      add_67_carry_2_port, add_67_carry_3_port, add_67_carry_4_port, 
      r83_carry_2_port, r83_carry_3_port, r83_carry_4_port, n1, n2, n3, n4, n5,
      n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32_port, n33_port
      , n34_port, n35, n36, n37, n38, n39, n40, n41, n42, n43_port, n44_port, 
      n45_port, n46_port, n47, n48_port, n49_port, n50_port, n51_port, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n187, n188, n189_port, n190_port, n191_port
      , n192_port, n193_port, n194, n195_port, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333_port, n334_port, n335_port, n336_port, n337_port, n338_port, 
      n339_port, n340_port, n341_port, n342_port, n343_port, n344_port, 
      n345_port, n346_port, n347_port, n348, n349, n350, n351, n352, n353, n354
      , n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n855, n857, n859, n861, n863, 
      n864, n865, n866, n867, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1064, 
      n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198 : std_logic;

begin
   DATA <= ( DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, 
      DATA_2_port, DATA_1_port, DATA_0_port );
   OUT_OPCODE <= ( OUT_OPCODE_1_port, OUT_OPCODE_0_port );
   EMPTY <= EMPTY_port;
   FULL <= FULL_port;
   
   X_Logic1_port <= '1';
   state_reg : DFFSR port map( D => X_Logic1_port, CLK => CLK, R => n85, S => 
                           n868, Q => state);
   FULL_reg : DFFPOSX1 port map( D => n1197, CLK => CLK, Q => FULL_port);
   memory_reg_0_7_inst : DFFPOSX1 port map( D => n1172, CLK => CLK, Q => 
                           memory_0_7_port);
   memory_reg_0_6_inst : DFFPOSX1 port map( D => n1171, CLK => CLK, Q => 
                           memory_0_6_port);
   memory_reg_0_5_inst : DFFPOSX1 port map( D => n1170, CLK => CLK, Q => 
                           memory_0_5_port);
   memory_reg_0_4_inst : DFFPOSX1 port map( D => n1169, CLK => CLK, Q => 
                           memory_0_4_port);
   memory_reg_0_3_inst : DFFPOSX1 port map( D => n1168, CLK => CLK, Q => 
                           memory_0_3_port);
   memory_reg_0_2_inst : DFFPOSX1 port map( D => n1071, CLK => CLK, Q => 
                           memory_0_2_port);
   memory_reg_0_1_inst : DFFPOSX1 port map( D => n1070, CLK => CLK, Q => 
                           memory_0_1_port);
   memory_reg_0_0_inst : DFFPOSX1 port map( D => n1069, CLK => CLK, Q => 
                           memory_0_0_port);
   memory_reg_1_7_inst : DFFPOSX1 port map( D => n1180, CLK => CLK, Q => 
                           memory_1_7_port);
   memory_reg_1_6_inst : DFFPOSX1 port map( D => n1179, CLK => CLK, Q => 
                           memory_1_6_port);
   memory_reg_1_5_inst : DFFPOSX1 port map( D => n1178, CLK => CLK, Q => 
                           memory_1_5_port);
   memory_reg_1_4_inst : DFFPOSX1 port map( D => n1177, CLK => CLK, Q => 
                           memory_1_4_port);
   memory_reg_1_3_inst : DFFPOSX1 port map( D => n1176, CLK => CLK, Q => 
                           memory_1_3_port);
   memory_reg_1_2_inst : DFFPOSX1 port map( D => n1175, CLK => CLK, Q => 
                           memory_1_2_port);
   memory_reg_1_1_inst : DFFPOSX1 port map( D => n1174, CLK => CLK, Q => 
                           memory_1_1_port);
   memory_reg_1_0_inst : DFFPOSX1 port map( D => n1173, CLK => CLK, Q => 
                           memory_1_0_port);
   memory_reg_2_7_inst : DFFPOSX1 port map( D => n1188, CLK => CLK, Q => 
                           memory_2_7_port);
   memory_reg_2_6_inst : DFFPOSX1 port map( D => n1187, CLK => CLK, Q => 
                           memory_2_6_port);
   memory_reg_2_5_inst : DFFPOSX1 port map( D => n1186, CLK => CLK, Q => 
                           memory_2_5_port);
   memory_reg_2_4_inst : DFFPOSX1 port map( D => n1185, CLK => CLK, Q => 
                           memory_2_4_port);
   memory_reg_2_3_inst : DFFPOSX1 port map( D => n1184, CLK => CLK, Q => 
                           memory_2_3_port);
   memory_reg_2_2_inst : DFFPOSX1 port map( D => n1183, CLK => CLK, Q => 
                           memory_2_2_port);
   memory_reg_2_1_inst : DFFPOSX1 port map( D => n1182, CLK => CLK, Q => 
                           memory_2_1_port);
   memory_reg_2_0_inst : DFFPOSX1 port map( D => n1181, CLK => CLK, Q => 
                           memory_2_0_port);
   memory_reg_3_7_inst : DFFPOSX1 port map( D => n1196, CLK => CLK, Q => 
                           memory_3_7_port);
   memory_reg_3_6_inst : DFFPOSX1 port map( D => n1195, CLK => CLK, Q => 
                           memory_3_6_port);
   memory_reg_3_5_inst : DFFPOSX1 port map( D => n1194, CLK => CLK, Q => 
                           memory_3_5_port);
   memory_reg_3_4_inst : DFFPOSX1 port map( D => n1193, CLK => CLK, Q => 
                           memory_3_4_port);
   memory_reg_3_3_inst : DFFPOSX1 port map( D => n1192, CLK => CLK, Q => 
                           memory_3_3_port);
   memory_reg_3_2_inst : DFFPOSX1 port map( D => n1191, CLK => CLK, Q => 
                           memory_3_2_port);
   memory_reg_3_1_inst : DFFPOSX1 port map( D => n1190, CLK => CLK, Q => 
                           memory_3_1_port);
   memory_reg_3_0_inst : DFFPOSX1 port map( D => n1189, CLK => CLK, Q => 
                           memory_3_0_port);
   memory_reg_4_7_inst : DFFPOSX1 port map( D => n869, CLK => CLK, Q => 
                           memory_4_7_port);
   memory_reg_4_6_inst : DFFPOSX1 port map( D => n870, CLK => CLK, Q => 
                           memory_4_6_port);
   memory_reg_4_5_inst : DFFPOSX1 port map( D => n871, CLK => CLK, Q => 
                           memory_4_5_port);
   memory_reg_4_4_inst : DFFPOSX1 port map( D => n872, CLK => CLK, Q => 
                           memory_4_4_port);
   memory_reg_4_3_inst : DFFPOSX1 port map( D => n873, CLK => CLK, Q => 
                           memory_4_3_port);
   memory_reg_4_2_inst : DFFPOSX1 port map( D => n874, CLK => CLK, Q => 
                           memory_4_2_port);
   memory_reg_4_1_inst : DFFPOSX1 port map( D => n875, CLK => CLK, Q => 
                           memory_4_1_port);
   memory_reg_4_0_inst : DFFPOSX1 port map( D => n876, CLK => CLK, Q => 
                           memory_4_0_port);
   memory_reg_5_7_inst : DFFPOSX1 port map( D => n879, CLK => CLK, Q => 
                           memory_5_7_port);
   memory_reg_5_6_inst : DFFPOSX1 port map( D => n880, CLK => CLK, Q => 
                           memory_5_6_port);
   memory_reg_5_5_inst : DFFPOSX1 port map( D => n881, CLK => CLK, Q => 
                           memory_5_5_port);
   memory_reg_5_4_inst : DFFPOSX1 port map( D => n882, CLK => CLK, Q => 
                           memory_5_4_port);
   memory_reg_5_3_inst : DFFPOSX1 port map( D => n883, CLK => CLK, Q => 
                           memory_5_3_port);
   memory_reg_5_2_inst : DFFPOSX1 port map( D => n884, CLK => CLK, Q => 
                           memory_5_2_port);
   memory_reg_5_1_inst : DFFPOSX1 port map( D => n885, CLK => CLK, Q => 
                           memory_5_1_port);
   memory_reg_5_0_inst : DFFPOSX1 port map( D => n886, CLK => CLK, Q => 
                           memory_5_0_port);
   memory_reg_6_7_inst : DFFPOSX1 port map( D => n889, CLK => CLK, Q => 
                           memory_6_7_port);
   memory_reg_6_6_inst : DFFPOSX1 port map( D => n890, CLK => CLK, Q => 
                           memory_6_6_port);
   memory_reg_6_5_inst : DFFPOSX1 port map( D => n891, CLK => CLK, Q => 
                           memory_6_5_port);
   memory_reg_6_4_inst : DFFPOSX1 port map( D => n892, CLK => CLK, Q => 
                           memory_6_4_port);
   memory_reg_6_3_inst : DFFPOSX1 port map( D => n893, CLK => CLK, Q => 
                           memory_6_3_port);
   memory_reg_6_2_inst : DFFPOSX1 port map( D => n894, CLK => CLK, Q => 
                           memory_6_2_port);
   memory_reg_6_1_inst : DFFPOSX1 port map( D => n895, CLK => CLK, Q => 
                           memory_6_1_port);
   memory_reg_6_0_inst : DFFPOSX1 port map( D => n896, CLK => CLK, Q => 
                           memory_6_0_port);
   memory_reg_7_7_inst : DFFPOSX1 port map( D => n899, CLK => CLK, Q => 
                           memory_7_7_port);
   memory_reg_7_6_inst : DFFPOSX1 port map( D => n900, CLK => CLK, Q => 
                           memory_7_6_port);
   memory_reg_7_5_inst : DFFPOSX1 port map( D => n901, CLK => CLK, Q => 
                           memory_7_5_port);
   memory_reg_7_4_inst : DFFPOSX1 port map( D => n902, CLK => CLK, Q => 
                           memory_7_4_port);
   memory_reg_7_3_inst : DFFPOSX1 port map( D => n903, CLK => CLK, Q => 
                           memory_7_3_port);
   memory_reg_7_2_inst : DFFPOSX1 port map( D => n904, CLK => CLK, Q => 
                           memory_7_2_port);
   memory_reg_7_1_inst : DFFPOSX1 port map( D => n905, CLK => CLK, Q => 
                           memory_7_1_port);
   memory_reg_7_0_inst : DFFPOSX1 port map( D => n906, CLK => CLK, Q => 
                           memory_7_0_port);
   memory_reg_8_7_inst : DFFPOSX1 port map( D => n1167, CLK => CLK, Q => 
                           memory_8_7_port);
   memory_reg_8_6_inst : DFFPOSX1 port map( D => n1166, CLK => CLK, Q => 
                           memory_8_6_port);
   memory_reg_8_5_inst : DFFPOSX1 port map( D => n1165, CLK => CLK, Q => 
                           memory_8_5_port);
   memory_reg_8_4_inst : DFFPOSX1 port map( D => n1164, CLK => CLK, Q => 
                           memory_8_4_port);
   memory_reg_8_3_inst : DFFPOSX1 port map( D => n1163, CLK => CLK, Q => 
                           memory_8_3_port);
   memory_reg_8_2_inst : DFFPOSX1 port map( D => n1162, CLK => CLK, Q => 
                           memory_8_2_port);
   memory_reg_8_1_inst : DFFPOSX1 port map( D => n1161, CLK => CLK, Q => 
                           memory_8_1_port);
   memory_reg_8_0_inst : DFFPOSX1 port map( D => n1160, CLK => CLK, Q => 
                           memory_8_0_port);
   memory_reg_9_7_inst : DFFPOSX1 port map( D => n1159, CLK => CLK, Q => 
                           memory_9_7_port);
   memory_reg_9_6_inst : DFFPOSX1 port map( D => n1158, CLK => CLK, Q => 
                           memory_9_6_port);
   memory_reg_9_5_inst : DFFPOSX1 port map( D => n1157, CLK => CLK, Q => 
                           memory_9_5_port);
   memory_reg_9_4_inst : DFFPOSX1 port map( D => n1156, CLK => CLK, Q => 
                           memory_9_4_port);
   memory_reg_9_3_inst : DFFPOSX1 port map( D => n1155, CLK => CLK, Q => 
                           memory_9_3_port);
   memory_reg_9_2_inst : DFFPOSX1 port map( D => n1154, CLK => CLK, Q => 
                           memory_9_2_port);
   memory_reg_9_1_inst : DFFPOSX1 port map( D => n1153, CLK => CLK, Q => 
                           memory_9_1_port);
   memory_reg_9_0_inst : DFFPOSX1 port map( D => n1152, CLK => CLK, Q => 
                           memory_9_0_port);
   memory_reg_10_7_inst : DFFPOSX1 port map( D => n1151, CLK => CLK, Q => 
                           memory_10_7_port);
   memory_reg_10_6_inst : DFFPOSX1 port map( D => n1150, CLK => CLK, Q => 
                           memory_10_6_port);
   memory_reg_10_5_inst : DFFPOSX1 port map( D => n1149, CLK => CLK, Q => 
                           memory_10_5_port);
   memory_reg_10_4_inst : DFFPOSX1 port map( D => n1148, CLK => CLK, Q => 
                           memory_10_4_port);
   memory_reg_10_3_inst : DFFPOSX1 port map( D => n1147, CLK => CLK, Q => 
                           memory_10_3_port);
   memory_reg_10_2_inst : DFFPOSX1 port map( D => n1146, CLK => CLK, Q => 
                           memory_10_2_port);
   memory_reg_10_1_inst : DFFPOSX1 port map( D => n1145, CLK => CLK, Q => 
                           memory_10_1_port);
   memory_reg_10_0_inst : DFFPOSX1 port map( D => n1144, CLK => CLK, Q => 
                           memory_10_0_port);
   memory_reg_11_7_inst : DFFPOSX1 port map( D => n1143, CLK => CLK, Q => 
                           memory_11_7_port);
   memory_reg_11_6_inst : DFFPOSX1 port map( D => n1142, CLK => CLK, Q => 
                           memory_11_6_port);
   memory_reg_11_5_inst : DFFPOSX1 port map( D => n1141, CLK => CLK, Q => 
                           memory_11_5_port);
   memory_reg_11_4_inst : DFFPOSX1 port map( D => n1140, CLK => CLK, Q => 
                           memory_11_4_port);
   memory_reg_11_3_inst : DFFPOSX1 port map( D => n1139, CLK => CLK, Q => 
                           memory_11_3_port);
   memory_reg_11_2_inst : DFFPOSX1 port map( D => n1138, CLK => CLK, Q => 
                           memory_11_2_port);
   memory_reg_11_1_inst : DFFPOSX1 port map( D => n1137, CLK => CLK, Q => 
                           memory_11_1_port);
   memory_reg_11_0_inst : DFFPOSX1 port map( D => n1136, CLK => CLK, Q => 
                           memory_11_0_port);
   memory_reg_12_7_inst : DFFPOSX1 port map( D => n1027, CLK => CLK, Q => 
                           memory_12_7_port);
   memory_reg_12_6_inst : DFFPOSX1 port map( D => n1028, CLK => CLK, Q => 
                           memory_12_6_port);
   memory_reg_12_5_inst : DFFPOSX1 port map( D => n1029, CLK => CLK, Q => 
                           memory_12_5_port);
   memory_reg_12_4_inst : DFFPOSX1 port map( D => n1064, CLK => CLK, Q => 
                           memory_12_4_port);
   memory_reg_12_3_inst : DFFPOSX1 port map( D => n1065, CLK => CLK, Q => 
                           memory_12_3_port);
   memory_reg_12_2_inst : DFFPOSX1 port map( D => n1066, CLK => CLK, Q => 
                           memory_12_2_port);
   memory_reg_12_1_inst : DFFPOSX1 port map( D => n1067, CLK => CLK, Q => 
                           memory_12_1_port);
   memory_reg_12_0_inst : DFFPOSX1 port map( D => n1068, CLK => CLK, Q => 
                           memory_12_0_port);
   memory_reg_13_7_inst : DFFPOSX1 port map( D => n1019, CLK => CLK, Q => 
                           memory_13_7_port);
   memory_reg_13_6_inst : DFFPOSX1 port map( D => n1020, CLK => CLK, Q => 
                           memory_13_6_port);
   memory_reg_13_5_inst : DFFPOSX1 port map( D => n1021, CLK => CLK, Q => 
                           memory_13_5_port);
   memory_reg_13_4_inst : DFFPOSX1 port map( D => n1022, CLK => CLK, Q => 
                           memory_13_4_port);
   memory_reg_13_3_inst : DFFPOSX1 port map( D => n1023, CLK => CLK, Q => 
                           memory_13_3_port);
   memory_reg_13_2_inst : DFFPOSX1 port map( D => n1024, CLK => CLK, Q => 
                           memory_13_2_port);
   memory_reg_13_1_inst : DFFPOSX1 port map( D => n1025, CLK => CLK, Q => 
                           memory_13_1_port);
   memory_reg_13_0_inst : DFFPOSX1 port map( D => n1026, CLK => CLK, Q => 
                           memory_13_0_port);
   memory_reg_14_7_inst : DFFPOSX1 port map( D => n1011, CLK => CLK, Q => 
                           memory_14_7_port);
   memory_reg_14_6_inst : DFFPOSX1 port map( D => n1012, CLK => CLK, Q => 
                           memory_14_6_port);
   memory_reg_14_5_inst : DFFPOSX1 port map( D => n1013, CLK => CLK, Q => 
                           memory_14_5_port);
   memory_reg_14_4_inst : DFFPOSX1 port map( D => n1014, CLK => CLK, Q => 
                           memory_14_4_port);
   memory_reg_14_3_inst : DFFPOSX1 port map( D => n1015, CLK => CLK, Q => 
                           memory_14_3_port);
   memory_reg_14_2_inst : DFFPOSX1 port map( D => n1016, CLK => CLK, Q => 
                           memory_14_2_port);
   memory_reg_14_1_inst : DFFPOSX1 port map( D => n1017, CLK => CLK, Q => 
                           memory_14_1_port);
   memory_reg_14_0_inst : DFFPOSX1 port map( D => n1018, CLK => CLK, Q => 
                           memory_14_0_port);
   memory_reg_15_7_inst : DFFPOSX1 port map( D => n1003, CLK => CLK, Q => 
                           memory_15_7_port);
   memory_reg_15_6_inst : DFFPOSX1 port map( D => n1004, CLK => CLK, Q => 
                           memory_15_6_port);
   memory_reg_15_5_inst : DFFPOSX1 port map( D => n1005, CLK => CLK, Q => 
                           memory_15_5_port);
   memory_reg_15_4_inst : DFFPOSX1 port map( D => n1006, CLK => CLK, Q => 
                           memory_15_4_port);
   memory_reg_15_3_inst : DFFPOSX1 port map( D => n1007, CLK => CLK, Q => 
                           memory_15_3_port);
   memory_reg_15_2_inst : DFFPOSX1 port map( D => n1008, CLK => CLK, Q => 
                           memory_15_2_port);
   memory_reg_15_1_inst : DFFPOSX1 port map( D => n1009, CLK => CLK, Q => 
                           memory_15_1_port);
   memory_reg_15_0_inst : DFFPOSX1 port map( D => n1010, CLK => CLK, Q => 
                           memory_15_0_port);
   memory_reg_16_7_inst : DFFPOSX1 port map( D => n1135, CLK => CLK, Q => 
                           memory_16_7_port);
   memory_reg_16_6_inst : DFFPOSX1 port map( D => n1134, CLK => CLK, Q => 
                           memory_16_6_port);
   memory_reg_16_5_inst : DFFPOSX1 port map( D => n1133, CLK => CLK, Q => 
                           memory_16_5_port);
   memory_reg_16_4_inst : DFFPOSX1 port map( D => n1132, CLK => CLK, Q => 
                           memory_16_4_port);
   memory_reg_16_3_inst : DFFPOSX1 port map( D => n1131, CLK => CLK, Q => 
                           memory_16_3_port);
   memory_reg_16_2_inst : DFFPOSX1 port map( D => n1130, CLK => CLK, Q => 
                           memory_16_2_port);
   memory_reg_16_1_inst : DFFPOSX1 port map( D => n1129, CLK => CLK, Q => 
                           memory_16_1_port);
   memory_reg_16_0_inst : DFFPOSX1 port map( D => n1128, CLK => CLK, Q => 
                           memory_16_0_port);
   memory_reg_17_7_inst : DFFPOSX1 port map( D => n1127, CLK => CLK, Q => 
                           memory_17_7_port);
   memory_reg_17_6_inst : DFFPOSX1 port map( D => n1126, CLK => CLK, Q => 
                           memory_17_6_port);
   memory_reg_17_5_inst : DFFPOSX1 port map( D => n1125, CLK => CLK, Q => 
                           memory_17_5_port);
   memory_reg_17_4_inst : DFFPOSX1 port map( D => n1124, CLK => CLK, Q => 
                           memory_17_4_port);
   memory_reg_17_3_inst : DFFPOSX1 port map( D => n1123, CLK => CLK, Q => 
                           memory_17_3_port);
   memory_reg_17_2_inst : DFFPOSX1 port map( D => n1122, CLK => CLK, Q => 
                           memory_17_2_port);
   memory_reg_17_1_inst : DFFPOSX1 port map( D => n1121, CLK => CLK, Q => 
                           memory_17_1_port);
   memory_reg_17_0_inst : DFFPOSX1 port map( D => n1120, CLK => CLK, Q => 
                           memory_17_0_port);
   memory_reg_18_7_inst : DFFPOSX1 port map( D => n1119, CLK => CLK, Q => 
                           memory_18_7_port);
   memory_reg_18_6_inst : DFFPOSX1 port map( D => n1118, CLK => CLK, Q => 
                           memory_18_6_port);
   memory_reg_18_5_inst : DFFPOSX1 port map( D => n1117, CLK => CLK, Q => 
                           memory_18_5_port);
   memory_reg_18_4_inst : DFFPOSX1 port map( D => n1116, CLK => CLK, Q => 
                           memory_18_4_port);
   memory_reg_18_3_inst : DFFPOSX1 port map( D => n1115, CLK => CLK, Q => 
                           memory_18_3_port);
   memory_reg_18_2_inst : DFFPOSX1 port map( D => n1114, CLK => CLK, Q => 
                           memory_18_2_port);
   memory_reg_18_1_inst : DFFPOSX1 port map( D => n1113, CLK => CLK, Q => 
                           memory_18_1_port);
   memory_reg_18_0_inst : DFFPOSX1 port map( D => n1112, CLK => CLK, Q => 
                           memory_18_0_port);
   memory_reg_19_7_inst : DFFPOSX1 port map( D => n1111, CLK => CLK, Q => 
                           memory_19_7_port);
   memory_reg_19_6_inst : DFFPOSX1 port map( D => n1110, CLK => CLK, Q => 
                           memory_19_6_port);
   memory_reg_19_5_inst : DFFPOSX1 port map( D => n1109, CLK => CLK, Q => 
                           memory_19_5_port);
   memory_reg_19_4_inst : DFFPOSX1 port map( D => n1108, CLK => CLK, Q => 
                           memory_19_4_port);
   memory_reg_19_3_inst : DFFPOSX1 port map( D => n1107, CLK => CLK, Q => 
                           memory_19_3_port);
   memory_reg_19_2_inst : DFFPOSX1 port map( D => n1106, CLK => CLK, Q => 
                           memory_19_2_port);
   memory_reg_19_1_inst : DFFPOSX1 port map( D => n1105, CLK => CLK, Q => 
                           memory_19_1_port);
   memory_reg_19_0_inst : DFFPOSX1 port map( D => n1104, CLK => CLK, Q => 
                           memory_19_0_port);
   memory_reg_20_7_inst : DFFPOSX1 port map( D => n995, CLK => CLK, Q => 
                           memory_20_7_port);
   memory_reg_20_6_inst : DFFPOSX1 port map( D => n996, CLK => CLK, Q => 
                           memory_20_6_port);
   memory_reg_20_5_inst : DFFPOSX1 port map( D => n997, CLK => CLK, Q => 
                           memory_20_5_port);
   memory_reg_20_4_inst : DFFPOSX1 port map( D => n998, CLK => CLK, Q => 
                           memory_20_4_port);
   memory_reg_20_3_inst : DFFPOSX1 port map( D => n999, CLK => CLK, Q => 
                           memory_20_3_port);
   memory_reg_20_2_inst : DFFPOSX1 port map( D => n1000, CLK => CLK, Q => 
                           memory_20_2_port);
   memory_reg_20_1_inst : DFFPOSX1 port map( D => n1001, CLK => CLK, Q => 
                           memory_20_1_port);
   memory_reg_20_0_inst : DFFPOSX1 port map( D => n1002, CLK => CLK, Q => 
                           memory_20_0_port);
   memory_reg_21_7_inst : DFFPOSX1 port map( D => n987, CLK => CLK, Q => 
                           memory_21_7_port);
   memory_reg_21_6_inst : DFFPOSX1 port map( D => n988, CLK => CLK, Q => 
                           memory_21_6_port);
   memory_reg_21_5_inst : DFFPOSX1 port map( D => n989, CLK => CLK, Q => 
                           memory_21_5_port);
   memory_reg_21_4_inst : DFFPOSX1 port map( D => n990, CLK => CLK, Q => 
                           memory_21_4_port);
   memory_reg_21_3_inst : DFFPOSX1 port map( D => n991, CLK => CLK, Q => 
                           memory_21_3_port);
   memory_reg_21_2_inst : DFFPOSX1 port map( D => n992, CLK => CLK, Q => 
                           memory_21_2_port);
   memory_reg_21_1_inst : DFFPOSX1 port map( D => n993, CLK => CLK, Q => 
                           memory_21_1_port);
   memory_reg_21_0_inst : DFFPOSX1 port map( D => n994, CLK => CLK, Q => 
                           memory_21_0_port);
   memory_reg_22_7_inst : DFFPOSX1 port map( D => n979, CLK => CLK, Q => 
                           memory_22_7_port);
   memory_reg_22_6_inst : DFFPOSX1 port map( D => n980, CLK => CLK, Q => 
                           memory_22_6_port);
   memory_reg_22_5_inst : DFFPOSX1 port map( D => n981, CLK => CLK, Q => 
                           memory_22_5_port);
   memory_reg_22_4_inst : DFFPOSX1 port map( D => n982, CLK => CLK, Q => 
                           memory_22_4_port);
   memory_reg_22_3_inst : DFFPOSX1 port map( D => n983, CLK => CLK, Q => 
                           memory_22_3_port);
   memory_reg_22_2_inst : DFFPOSX1 port map( D => n984, CLK => CLK, Q => 
                           memory_22_2_port);
   memory_reg_22_1_inst : DFFPOSX1 port map( D => n985, CLK => CLK, Q => 
                           memory_22_1_port);
   memory_reg_22_0_inst : DFFPOSX1 port map( D => n986, CLK => CLK, Q => 
                           memory_22_0_port);
   memory_reg_23_7_inst : DFFPOSX1 port map( D => n971, CLK => CLK, Q => 
                           memory_23_7_port);
   memory_reg_23_6_inst : DFFPOSX1 port map( D => n972, CLK => CLK, Q => 
                           memory_23_6_port);
   memory_reg_23_5_inst : DFFPOSX1 port map( D => n973, CLK => CLK, Q => 
                           memory_23_5_port);
   memory_reg_23_4_inst : DFFPOSX1 port map( D => n974, CLK => CLK, Q => 
                           memory_23_4_port);
   memory_reg_23_3_inst : DFFPOSX1 port map( D => n975, CLK => CLK, Q => 
                           memory_23_3_port);
   memory_reg_23_2_inst : DFFPOSX1 port map( D => n976, CLK => CLK, Q => 
                           memory_23_2_port);
   memory_reg_23_1_inst : DFFPOSX1 port map( D => n977, CLK => CLK, Q => 
                           memory_23_1_port);
   memory_reg_23_0_inst : DFFPOSX1 port map( D => n978, CLK => CLK, Q => 
                           memory_23_0_port);
   memory_reg_24_7_inst : DFFPOSX1 port map( D => n963, CLK => CLK, Q => 
                           memory_24_7_port);
   memory_reg_24_6_inst : DFFPOSX1 port map( D => n964, CLK => CLK, Q => 
                           memory_24_6_port);
   memory_reg_24_5_inst : DFFPOSX1 port map( D => n965, CLK => CLK, Q => 
                           memory_24_5_port);
   memory_reg_24_4_inst : DFFPOSX1 port map( D => n966, CLK => CLK, Q => 
                           memory_24_4_port);
   memory_reg_24_3_inst : DFFPOSX1 port map( D => n967, CLK => CLK, Q => 
                           memory_24_3_port);
   memory_reg_24_2_inst : DFFPOSX1 port map( D => n968, CLK => CLK, Q => 
                           memory_24_2_port);
   memory_reg_24_1_inst : DFFPOSX1 port map( D => n969, CLK => CLK, Q => 
                           memory_24_1_port);
   memory_reg_24_0_inst : DFFPOSX1 port map( D => n970, CLK => CLK, Q => 
                           memory_24_0_port);
   memory_reg_25_7_inst : DFFPOSX1 port map( D => n955, CLK => CLK, Q => 
                           memory_25_7_port);
   memory_reg_25_6_inst : DFFPOSX1 port map( D => n956, CLK => CLK, Q => 
                           memory_25_6_port);
   memory_reg_25_5_inst : DFFPOSX1 port map( D => n957, CLK => CLK, Q => 
                           memory_25_5_port);
   memory_reg_25_4_inst : DFFPOSX1 port map( D => n958, CLK => CLK, Q => 
                           memory_25_4_port);
   memory_reg_25_3_inst : DFFPOSX1 port map( D => n959, CLK => CLK, Q => 
                           memory_25_3_port);
   memory_reg_25_2_inst : DFFPOSX1 port map( D => n960, CLK => CLK, Q => 
                           memory_25_2_port);
   memory_reg_25_1_inst : DFFPOSX1 port map( D => n961, CLK => CLK, Q => 
                           memory_25_1_port);
   memory_reg_25_0_inst : DFFPOSX1 port map( D => n962, CLK => CLK, Q => 
                           memory_25_0_port);
   memory_reg_26_7_inst : DFFPOSX1 port map( D => n947, CLK => CLK, Q => 
                           memory_26_7_port);
   memory_reg_26_6_inst : DFFPOSX1 port map( D => n948, CLK => CLK, Q => 
                           memory_26_6_port);
   memory_reg_26_5_inst : DFFPOSX1 port map( D => n949, CLK => CLK, Q => 
                           memory_26_5_port);
   memory_reg_26_4_inst : DFFPOSX1 port map( D => n950, CLK => CLK, Q => 
                           memory_26_4_port);
   memory_reg_26_3_inst : DFFPOSX1 port map( D => n951, CLK => CLK, Q => 
                           memory_26_3_port);
   memory_reg_26_2_inst : DFFPOSX1 port map( D => n952, CLK => CLK, Q => 
                           memory_26_2_port);
   memory_reg_26_1_inst : DFFPOSX1 port map( D => n953, CLK => CLK, Q => 
                           memory_26_1_port);
   memory_reg_26_0_inst : DFFPOSX1 port map( D => n954, CLK => CLK, Q => 
                           memory_26_0_port);
   memory_reg_27_7_inst : DFFPOSX1 port map( D => n939, CLK => CLK, Q => 
                           memory_27_7_port);
   memory_reg_27_6_inst : DFFPOSX1 port map( D => n940, CLK => CLK, Q => 
                           memory_27_6_port);
   memory_reg_27_5_inst : DFFPOSX1 port map( D => n941, CLK => CLK, Q => 
                           memory_27_5_port);
   memory_reg_27_4_inst : DFFPOSX1 port map( D => n942, CLK => CLK, Q => 
                           memory_27_4_port);
   memory_reg_27_3_inst : DFFPOSX1 port map( D => n943, CLK => CLK, Q => 
                           memory_27_3_port);
   memory_reg_27_2_inst : DFFPOSX1 port map( D => n944, CLK => CLK, Q => 
                           memory_27_2_port);
   memory_reg_27_1_inst : DFFPOSX1 port map( D => n945, CLK => CLK, Q => 
                           memory_27_1_port);
   memory_reg_27_0_inst : DFFPOSX1 port map( D => n946, CLK => CLK, Q => 
                           memory_27_0_port);
   memory_reg_28_7_inst : DFFPOSX1 port map( D => n1103, CLK => CLK, Q => 
                           memory_28_7_port);
   memory_reg_28_6_inst : DFFPOSX1 port map( D => n1102, CLK => CLK, Q => 
                           memory_28_6_port);
   memory_reg_28_5_inst : DFFPOSX1 port map( D => n1101, CLK => CLK, Q => 
                           memory_28_5_port);
   memory_reg_28_4_inst : DFFPOSX1 port map( D => n1100, CLK => CLK, Q => 
                           memory_28_4_port);
   memory_reg_28_3_inst : DFFPOSX1 port map( D => n1099, CLK => CLK, Q => 
                           memory_28_3_port);
   memory_reg_28_2_inst : DFFPOSX1 port map( D => n1098, CLK => CLK, Q => 
                           memory_28_2_port);
   memory_reg_28_1_inst : DFFPOSX1 port map( D => n1097, CLK => CLK, Q => 
                           memory_28_1_port);
   memory_reg_28_0_inst : DFFPOSX1 port map( D => n1096, CLK => CLK, Q => 
                           memory_28_0_port);
   memory_reg_29_7_inst : DFFPOSX1 port map( D => n1095, CLK => CLK, Q => 
                           memory_29_7_port);
   memory_reg_29_6_inst : DFFPOSX1 port map( D => n1094, CLK => CLK, Q => 
                           memory_29_6_port);
   memory_reg_29_5_inst : DFFPOSX1 port map( D => n1093, CLK => CLK, Q => 
                           memory_29_5_port);
   memory_reg_29_4_inst : DFFPOSX1 port map( D => n1092, CLK => CLK, Q => 
                           memory_29_4_port);
   memory_reg_29_3_inst : DFFPOSX1 port map( D => n1091, CLK => CLK, Q => 
                           memory_29_3_port);
   memory_reg_29_2_inst : DFFPOSX1 port map( D => n1090, CLK => CLK, Q => 
                           memory_29_2_port);
   memory_reg_29_1_inst : DFFPOSX1 port map( D => n1089, CLK => CLK, Q => 
                           memory_29_1_port);
   memory_reg_29_0_inst : DFFPOSX1 port map( D => n1088, CLK => CLK, Q => 
                           memory_29_0_port);
   memory_reg_30_7_inst : DFFPOSX1 port map( D => n1087, CLK => CLK, Q => 
                           memory_30_7_port);
   memory_reg_30_6_inst : DFFPOSX1 port map( D => n1086, CLK => CLK, Q => 
                           memory_30_6_port);
   memory_reg_30_5_inst : DFFPOSX1 port map( D => n1085, CLK => CLK, Q => 
                           memory_30_5_port);
   memory_reg_30_4_inst : DFFPOSX1 port map( D => n1084, CLK => CLK, Q => 
                           memory_30_4_port);
   memory_reg_30_3_inst : DFFPOSX1 port map( D => n1083, CLK => CLK, Q => 
                           memory_30_3_port);
   memory_reg_30_2_inst : DFFPOSX1 port map( D => n1082, CLK => CLK, Q => 
                           memory_30_2_port);
   memory_reg_30_1_inst : DFFPOSX1 port map( D => n1081, CLK => CLK, Q => 
                           memory_30_1_port);
   memory_reg_30_0_inst : DFFPOSX1 port map( D => n1080, CLK => CLK, Q => 
                           memory_30_0_port);
   memory_reg_31_7_inst : DFFPOSX1 port map( D => n1079, CLK => CLK, Q => 
                           memory_31_7_port);
   memory_reg_31_6_inst : DFFPOSX1 port map( D => n1078, CLK => CLK, Q => 
                           memory_31_6_port);
   memory_reg_31_5_inst : DFFPOSX1 port map( D => n1077, CLK => CLK, Q => 
                           memory_31_5_port);
   memory_reg_31_4_inst : DFFPOSX1 port map( D => n1076, CLK => CLK, Q => 
                           memory_31_4_port);
   memory_reg_31_3_inst : DFFPOSX1 port map( D => n1075, CLK => CLK, Q => 
                           memory_31_3_port);
   memory_reg_31_2_inst : DFFPOSX1 port map( D => n1074, CLK => CLK, Q => 
                           memory_31_2_port);
   memory_reg_31_1_inst : DFFPOSX1 port map( D => n1073, CLK => CLK, Q => 
                           memory_31_1_port);
   memory_reg_31_0_inst : DFFPOSX1 port map( D => n1072, CLK => CLK, Q => 
                           memory_31_0_port);
   opcode_reg_0_1_inst : DFFPOSX1 port map( D => n932, CLK => CLK, Q => 
                           opcode_0_1_port);
   opcode_reg_0_0_inst : DFFPOSX1 port map( D => n931, CLK => CLK, Q => 
                           opcode_0_0_port);
   opcode_reg_1_1_inst : DFFPOSX1 port map( D => n934, CLK => CLK, Q => 
                           opcode_1_1_port);
   opcode_reg_1_0_inst : DFFPOSX1 port map( D => n933, CLK => CLK, Q => 
                           opcode_1_0_port);
   opcode_reg_2_1_inst : DFFPOSX1 port map( D => n936, CLK => CLK, Q => 
                           opcode_2_1_port);
   opcode_reg_2_0_inst : DFFPOSX1 port map( D => n935, CLK => CLK, Q => 
                           opcode_2_0_port);
   opcode_reg_3_1_inst : DFFPOSX1 port map( D => n938, CLK => CLK, Q => 
                           opcode_3_1_port);
   opcode_reg_3_0_inst : DFFPOSX1 port map( D => n937, CLK => CLK, Q => 
                           opcode_3_0_port);
   opcode_reg_4_1_inst : DFFPOSX1 port map( D => n877, CLK => CLK, Q => 
                           opcode_4_1_port);
   opcode_reg_4_0_inst : DFFPOSX1 port map( D => n878, CLK => CLK, Q => 
                           opcode_4_0_port);
   opcode_reg_5_1_inst : DFFPOSX1 port map( D => n887, CLK => CLK, Q => 
                           opcode_5_1_port);
   opcode_reg_5_0_inst : DFFPOSX1 port map( D => n888, CLK => CLK, Q => 
                           opcode_5_0_port);
   opcode_reg_6_1_inst : DFFPOSX1 port map( D => n897, CLK => CLK, Q => 
                           opcode_6_1_port);
   opcode_reg_6_0_inst : DFFPOSX1 port map( D => n898, CLK => CLK, Q => 
                           opcode_6_0_port);
   opcode_reg_7_1_inst : DFFPOSX1 port map( D => n907, CLK => CLK, Q => 
                           opcode_7_1_port);
   opcode_reg_7_0_inst : DFFPOSX1 port map( D => n908, CLK => CLK, Q => 
                           opcode_7_0_port);
   opcode_reg_8_1_inst : DFFPOSX1 port map( D => n1063, CLK => CLK, Q => 
                           opcode_8_1_port);
   opcode_reg_8_0_inst : DFFPOSX1 port map( D => n1062, CLK => CLK, Q => 
                           opcode_8_0_port);
   opcode_reg_9_1_inst : DFFPOSX1 port map( D => n1061, CLK => CLK, Q => 
                           opcode_9_1_port);
   opcode_reg_9_0_inst : DFFPOSX1 port map( D => n1060, CLK => CLK, Q => 
                           opcode_9_0_port);
   opcode_reg_10_1_inst : DFFPOSX1 port map( D => n1059, CLK => CLK, Q => 
                           opcode_10_1_port);
   opcode_reg_10_0_inst : DFFPOSX1 port map( D => n1058, CLK => CLK, Q => 
                           opcode_10_0_port);
   opcode_reg_11_1_inst : DFFPOSX1 port map( D => n1057, CLK => CLK, Q => 
                           opcode_11_1_port);
   opcode_reg_11_0_inst : DFFPOSX1 port map( D => n1056, CLK => CLK, Q => 
                           opcode_11_0_port);
   opcode_reg_12_1_inst : DFFPOSX1 port map( D => n929, CLK => CLK, Q => 
                           opcode_12_1_port);
   opcode_reg_12_0_inst : DFFPOSX1 port map( D => n930, CLK => CLK, Q => 
                           opcode_12_0_port);
   opcode_reg_13_1_inst : DFFPOSX1 port map( D => n927, CLK => CLK, Q => 
                           opcode_13_1_port);
   opcode_reg_13_0_inst : DFFPOSX1 port map( D => n928, CLK => CLK, Q => 
                           opcode_13_0_port);
   opcode_reg_14_1_inst : DFFPOSX1 port map( D => n925, CLK => CLK, Q => 
                           opcode_14_1_port);
   opcode_reg_14_0_inst : DFFPOSX1 port map( D => n926, CLK => CLK, Q => 
                           opcode_14_0_port);
   opcode_reg_15_1_inst : DFFPOSX1 port map( D => n923, CLK => CLK, Q => 
                           opcode_15_1_port);
   opcode_reg_15_0_inst : DFFPOSX1 port map( D => n924, CLK => CLK, Q => 
                           opcode_15_0_port);
   opcode_reg_16_1_inst : DFFPOSX1 port map( D => n1055, CLK => CLK, Q => 
                           opcode_16_1_port);
   opcode_reg_16_0_inst : DFFPOSX1 port map( D => n1054, CLK => CLK, Q => 
                           opcode_16_0_port);
   opcode_reg_17_1_inst : DFFPOSX1 port map( D => n1053, CLK => CLK, Q => 
                           opcode_17_1_port);
   opcode_reg_17_0_inst : DFFPOSX1 port map( D => n1052, CLK => CLK, Q => 
                           opcode_17_0_port);
   opcode_reg_18_1_inst : DFFPOSX1 port map( D => n1051, CLK => CLK, Q => 
                           opcode_18_1_port);
   opcode_reg_18_0_inst : DFFPOSX1 port map( D => n1050, CLK => CLK, Q => 
                           opcode_18_0_port);
   opcode_reg_19_1_inst : DFFPOSX1 port map( D => n1049, CLK => CLK, Q => 
                           opcode_19_1_port);
   opcode_reg_19_0_inst : DFFPOSX1 port map( D => n1048, CLK => CLK, Q => 
                           opcode_19_0_port);
   opcode_reg_20_1_inst : DFFPOSX1 port map( D => n921, CLK => CLK, Q => 
                           opcode_20_1_port);
   opcode_reg_20_0_inst : DFFPOSX1 port map( D => n922, CLK => CLK, Q => 
                           opcode_20_0_port);
   opcode_reg_21_1_inst : DFFPOSX1 port map( D => n919, CLK => CLK, Q => 
                           opcode_21_1_port);
   opcode_reg_21_0_inst : DFFPOSX1 port map( D => n920, CLK => CLK, Q => 
                           opcode_21_0_port);
   opcode_reg_22_1_inst : DFFPOSX1 port map( D => n917, CLK => CLK, Q => 
                           opcode_22_1_port);
   opcode_reg_22_0_inst : DFFPOSX1 port map( D => n918, CLK => CLK, Q => 
                           opcode_22_0_port);
   opcode_reg_23_1_inst : DFFPOSX1 port map( D => n915, CLK => CLK, Q => 
                           opcode_23_1_port);
   opcode_reg_23_0_inst : DFFPOSX1 port map( D => n916, CLK => CLK, Q => 
                           opcode_23_0_port);
   opcode_reg_24_1_inst : DFFPOSX1 port map( D => n913, CLK => CLK, Q => 
                           opcode_24_1_port);
   opcode_reg_24_0_inst : DFFPOSX1 port map( D => n914, CLK => CLK, Q => 
                           opcode_24_0_port);
   opcode_reg_25_1_inst : DFFPOSX1 port map( D => n911, CLK => CLK, Q => 
                           opcode_25_1_port);
   opcode_reg_25_0_inst : DFFPOSX1 port map( D => n912, CLK => CLK, Q => 
                           opcode_25_0_port);
   opcode_reg_26_1_inst : DFFPOSX1 port map( D => n909, CLK => CLK, Q => 
                           opcode_26_1_port);
   opcode_reg_26_0_inst : DFFPOSX1 port map( D => n910, CLK => CLK, Q => 
                           opcode_26_0_port);
   opcode_reg_27_1_inst : DFFPOSX1 port map( D => n866, CLK => CLK, Q => 
                           opcode_27_1_port);
   opcode_reg_27_0_inst : DFFPOSX1 port map( D => n867, CLK => CLK, Q => 
                           opcode_27_0_port);
   opcode_reg_28_1_inst : DFFPOSX1 port map( D => n1047, CLK => CLK, Q => 
                           opcode_28_1_port);
   opcode_reg_28_0_inst : DFFPOSX1 port map( D => n1046, CLK => CLK, Q => 
                           opcode_28_0_port);
   opcode_reg_29_1_inst : DFFPOSX1 port map( D => n1045, CLK => CLK, Q => 
                           opcode_29_1_port);
   opcode_reg_29_0_inst : DFFPOSX1 port map( D => n1044, CLK => CLK, Q => 
                           opcode_29_0_port);
   opcode_reg_30_1_inst : DFFPOSX1 port map( D => n1043, CLK => CLK, Q => 
                           opcode_30_1_port);
   opcode_reg_30_0_inst : DFFPOSX1 port map( D => n1042, CLK => CLK, Q => 
                           opcode_30_0_port);
   opcode_reg_31_1_inst : DFFPOSX1 port map( D => n1041, CLK => CLK, Q => 
                           opcode_31_1_port);
   opcode_reg_31_0_inst : DFFPOSX1 port map( D => n1040, CLK => CLK, Q => 
                           opcode_31_0_port);
   DATA_reg_7_inst : DFFPOSX1 port map( D => n1039, CLK => CLK, Q => 
                           DATA_7_port);
   DATA_reg_6_inst : DFFPOSX1 port map( D => n1038, CLK => CLK, Q => 
                           DATA_6_port);
   DATA_reg_5_inst : DFFPOSX1 port map( D => n1037, CLK => CLK, Q => 
                           DATA_5_port);
   DATA_reg_4_inst : DFFPOSX1 port map( D => n1036, CLK => CLK, Q => 
                           DATA_4_port);
   DATA_reg_3_inst : DFFPOSX1 port map( D => n1035, CLK => CLK, Q => 
                           DATA_3_port);
   DATA_reg_2_inst : DFFPOSX1 port map( D => n1034, CLK => CLK, Q => 
                           DATA_2_port);
   DATA_reg_1_inst : DFFPOSX1 port map( D => n1033, CLK => CLK, Q => 
                           DATA_1_port);
   DATA_reg_0_inst : DFFPOSX1 port map( D => n1032, CLK => CLK, Q => 
                           DATA_0_port);
   OUT_OPCODE_reg_1_inst : DFFPOSX1 port map( D => n1031, CLK => CLK, Q => 
                           OUT_OPCODE_1_port);
   OUT_OPCODE_reg_0_inst : DFFPOSX1 port map( D => n1030, CLK => CLK, Q => 
                           OUT_OPCODE_0_port);
   EMPTY_reg : DFFPOSX1 port map( D => n1198, CLK => CLK, Q => EMPTY_port);
   n868 <= '1';
   sub_72_U2_1 : FAX1 port map( A => n67, B => n514, C => sub_72_carry_1_port, 
                           YC => sub_72_carry_2_port, YS => N190);
   sub_72_U2_2 : FAX1 port map( A => n65, B => n851, C => sub_72_carry_2_port, 
                           YC => sub_72_carry_3_port, YS => N191);
   sub_72_U2_3 : FAX1 port map( A => n71, B => n821, C => sub_72_carry_3_port, 
                           YC => sub_72_carry_4_port, YS => N192);
   sub_72_U2_4 : FAX1 port map( A => writeptr_4_port, B => n842, C => 
                           sub_72_carry_4_port, YC => n90, YS => N193);
   add_67_U1_1_1 : HAX1 port map( A => n67, B => n69, YC => add_67_carry_2_port
                           , YS => N48);
   add_67_U1_1_2 : HAX1 port map( A => n65, B => add_67_carry_2_port, YC => 
                           add_67_carry_3_port, YS => N49);
   add_67_U1_1_3 : HAX1 port map( A => n71, B => add_67_carry_3_port, YC => 
                           add_67_carry_4_port, YS => N50);
   r83_U1_1_1 : HAX1 port map( A => writeptr_1_port, B => writeptr_0_port, YC 
                           => r83_carry_2_port, YS => N32);
   r83_U1_1_2 : HAX1 port map( A => writeptr_2_port, B => r83_carry_2_port, YC 
                           => r83_carry_3_port, YS => N33);
   r83_U1_1_3 : HAX1 port map( A => writeptr_3_port, B => r83_carry_3_port, YC 
                           => r83_carry_4_port, YS => N34);
   BYTE_COUNT_reg_0_inst : DFFSR port map( D => N338, CLK => CLK, R => n85, S 
                           => n18, Q => BYTE_COUNT(0));
   BYTE_COUNT_reg_1_inst : DFFSR port map( D => N339, CLK => CLK, R => n85, S 
                           => n17, Q => BYTE_COUNT(1));
   BYTE_COUNT_reg_2_inst : DFFSR port map( D => N340, CLK => CLK, R => n85, S 
                           => n16, Q => BYTE_COUNT(2));
   readptr_reg_0_inst : DFFSR port map( D => N343, CLK => CLK, R => n85, S => 
                           n15, Q => readptr_0_port);
   BYTE_COUNT_reg_3_inst : DFFSR port map( D => N341, CLK => CLK, R => n85, S 
                           => n14, Q => BYTE_COUNT(3));
   readptr_reg_1_inst : DFFSR port map( D => N344, CLK => CLK, R => n85, S => 
                           n13, Q => readptr_1_port);
   BYTE_COUNT_reg_4_inst : DFFSR port map( D => N342, CLK => CLK, R => n85, S 
                           => n12, Q => BYTE_COUNT(4));
   readptr_reg_2_inst : DFFSR port map( D => N345, CLK => CLK, R => n85, S => 
                           n11, Q => readptr_2_port);
   readptr_reg_3_inst : DFFSR port map( D => N346, CLK => CLK, R => n85, S => 
                           n10, Q => readptr_3_port);
   writeptr_reg_4_inst : DFFSR port map( D => n862, CLK => CLK, R => n85, S => 
                           n9, Q => writeptr_4_port);
   writeptr_reg_3_inst : DFFSR port map( D => n860, CLK => CLK, R => n85, S => 
                           n8, Q => writeptr_3_port);
   writeptr_reg_2_inst : DFFSR port map( D => n854, CLK => CLK, R => n85, S => 
                           n7, Q => writeptr_2_port);
   writeptr_reg_1_inst : DFFSR port map( D => n856, CLK => CLK, R => n85, S => 
                           n6, Q => writeptr_1_port);
   writeptr_reg_0_inst : DFFSR port map( D => n858, CLK => CLK, R => n85, S => 
                           n5, Q => writeptr_0_port);
   readptr_reg_4_inst : DFFSR port map( D => N347, CLK => CLK, R => n85, S => 
                           n4, Q => readptr_4_port);
   U3 : BUFX2 port map( A => n351, Y => n63);
   U4 : BUFX2 port map( A => n277, Y => n20);
   U5 : BUFX2 port map( A => n449, Y => n62);
   U6 : INVX2 port map( A => n34_port, Y => n61);
   U7 : INVX2 port map( A => n33_port, Y => n45_port);
   U8 : BUFX2 port map( A => n116, Y => n46_port);
   U9 : INVX4 port map( A => n26, Y => n121);
   U10 : INVX2 port map( A => n27, Y => n47);
   U11 : INVX2 port map( A => n28, Y => n48_port);
   U12 : INVX2 port map( A => n29, Y => n60);
   U13 : INVX2 port map( A => n30, Y => n59);
   U14 : INVX2 port map( A => n31, Y => n58);
   U15 : INVX2 port map( A => n32_port, Y => n57);
   U16 : INVX2 port map( A => n35, Y => n53);
   U17 : INVX2 port map( A => n36, Y => n54);
   U18 : INVX2 port map( A => n40, Y => n55);
   U19 : INVX2 port map( A => n41, Y => n56);
   U20 : INVX2 port map( A => n39, Y => n52);
   U21 : INVX2 port map( A => n37, Y => n51_port);
   U22 : INVX2 port map( A => n2, Y => n50_port);
   U23 : INVX2 port map( A => n38, Y => n49_port);
   U24 : AND2X2 port map( A => n493, B => n70, Y => n1);
   U25 : OR2X2 port map( A => n19, B => n134, Y => n2);
   U26 : AND2X2 port map( A => n493, B => n71, Y => n3);
   n4 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n15 <= '1';
   n16 <= '1';
   n17 <= '1';
   n18 <= '1';
   U42 : INVX2 port map( A => n146, Y => n309);
   U43 : NAND2X1 port map( A => n63, B => n3, Y => n174);
   U44 : NAND2X1 port map( A => n63, B => n1, Y => n209);
   U45 : BUFX2 port map( A => n277, Y => n19);
   U46 : INVX2 port map( A => n135, Y => n126);
   U47 : INVX2 port map( A => writeptr_0_port, Y => n68);
   U48 : INVX2 port map( A => writeptr_1_port, Y => n66);
   U49 : OR2X2 port map( A => n145, B => n174, Y => n21);
   U50 : INVX4 port map( A => n21, Y => n458);
   U51 : OR2X2 port map( A => n134, B => n174, Y => n22);
   U52 : INVX4 port map( A => n22, Y => n106);
   U53 : OR2X2 port map( A => n184, B => n174, Y => n23);
   U54 : INVX4 port map( A => n23, Y => n101);
   U55 : OR2X2 port map( A => n140, B => n174, Y => n24);
   U56 : INVX4 port map( A => n24, Y => n111);
   U57 : OR2X2 port map( A => n235, B => n174, Y => n25);
   U58 : INVX4 port map( A => n25, Y => n432);
   U59 : OR2X2 port map( A => n151, B => n209, Y => n26);
   U60 : OR2X2 port map( A => n209, B => n226, Y => n27);
   U61 : OR2X2 port map( A => n209, B => n235, Y => n28);
   U62 : OR2X2 port map( A => n209, B => n175, Y => n29);
   U63 : OR2X2 port map( A => n209, B => n184, Y => n30);
   U64 : OR2X2 port map( A => n209, B => n134, Y => n31);
   U65 : OR2X2 port map( A => n209, B => n140, Y => n32_port);
   U66 : OR2X2 port map( A => n174, B => n175, Y => n33_port);
   U67 : OR2X2 port map( A => n174, B => n226, Y => n34_port);
   U68 : INVX2 port map( A => RCV_OPCODE(0), Y => n76);
   U69 : OR2X2 port map( A => n20, B => n145, Y => n35);
   U70 : OR2X2 port map( A => n20, B => n151, Y => n36);
   U71 : INVX2 port map( A => n500, Y => n96);
   U72 : XNOR2X1 port map( A => readptr_0_port, B => n69, Y => n516);
   U73 : OR2X2 port map( A => n19, B => n184, Y => n37);
   U74 : OR2X2 port map( A => n19, B => n140, Y => n38);
   U75 : OR2X2 port map( A => n20, B => n175, Y => n39);
   U76 : OR2X2 port map( A => n20, B => n226, Y => n40);
   U77 : OR2X2 port map( A => n20, B => n235, Y => n41);
   U78 : INVX2 port map( A => RST, Y => n85);
   U79 : INVX2 port map( A => n508, Y => n156);
   U80 : INVX2 port map( A => n68, Y => n69);
   U81 : INVX2 port map( A => n66, Y => n67);
   U82 : INVX2 port map( A => n70, Y => n71);
   U83 : INVX2 port map( A => n64, Y => n65);
   U84 : INVX2 port map( A => RCV_DATA(7), Y => n77);
   U85 : INVX2 port map( A => RCV_DATA(1), Y => n83);
   U86 : INVX2 port map( A => RCV_DATA(3), Y => n81);
   U87 : INVX2 port map( A => RCV_DATA(5), Y => n79);
   U88 : INVX2 port map( A => RCV_DATA(0), Y => n84);
   U89 : INVX2 port map( A => RCV_DATA(2), Y => n82);
   U90 : INVX2 port map( A => RCV_DATA(4), Y => n80);
   U91 : INVX2 port map( A => RCV_DATA(6), Y => n78);
   U92 : XNOR2X1 port map( A => readptr_4_port, B => n42, Y => n513);
   U93 : XNOR2X1 port map( A => r83_carry_4_port, B => writeptr_4_port, Y => 
                           n42);
   U94 : INVX2 port map( A => writeptr_2_port, Y => n64);
   U95 : INVX2 port map( A => writeptr_3_port, Y => n70);
   U96 : BUFX2 port map( A => state, Y => n72);
   U97 : INVX2 port map( A => RCV_OPCODE(0), Y => n93);
   U98 : INVX2 port map( A => n507, Y => n353);
   U99 : INVX1 port map( A => n63, Y => n43_port);
   U100 : INVX2 port map( A => n43_port, Y => n44_port);
   U101 : AND2X2 port map( A => n475, B => n63, Y => n244);
   U102 : INVX1 port map( A => RCV_OPCODE(1), Y => n73);
   U103 : INVX1 port map( A => RCV_OPCODE(1), Y => n74);
   U104 : AND2X2 port map( A => RCV_OPCODE(1), B => RCV_OPCODE(0), Y => n480);
   U105 : INVX1 port map( A => RCV_OPCODE(1), Y => n75);
   U106 : AND2X2 port map( A => n480, B => n353, Y => n356);
   U107 : AND2X2 port map( A => n815, B => n817, Y => n534);
   U108 : AND2X2 port map( A => n813, B => n817, Y => n533);
   U109 : AND2X2 port map( A => n815, B => n818, Y => n536);
   U110 : AND2X2 port map( A => n813, B => n818, Y => n535);
   U111 : AND2X2 port map( A => n829, B => n817, Y => n547);
   U112 : AND2X2 port map( A => n817, B => n828, Y => n546);
   U113 : AND2X2 port map( A => n818, B => n829, Y => n549);
   U114 : AND2X2 port map( A => n818, B => n828, Y => n548);
   U115 : AND2X2 port map( A => n840, B => n818, Y => n562);
   U116 : AND2X2 port map( A => n839, B => n818, Y => n561);
   U117 : AND2X2 port map( A => n840, B => n817, Y => n564);
   U118 : AND2X2 port map( A => n839, B => n817, Y => n563);
   U119 : AND2X2 port map( A => n850, B => n817, Y => n575);
   U120 : AND2X2 port map( A => n849, B => n817, Y => n574);
   U121 : AND2X2 port map( A => n850, B => n818, Y => n577);
   U122 : AND2X2 port map( A => n849, B => n818, Y => n576);
   U123 : OR2X1 port map( A => n820, B => n69, Y => sub_72_carry_1_port);
   U124 : XNOR2X1 port map( A => n69, B => n820, Y => N189);
   U125 : XOR2X1 port map( A => readptr_4_port, B => add_76_aco_carry_4_port, Y
                           => N337);
   U126 : AND2X1 port map( A => readptr_3_port, B => add_76_aco_carry_3_port, Y
                           => add_76_aco_carry_4_port);
   U127 : XOR2X1 port map( A => add_76_aco_carry_3_port, B => readptr_3_port, Y
                           => N336);
   U128 : AND2X1 port map( A => readptr_2_port, B => add_76_aco_carry_2_port, Y
                           => add_76_aco_carry_3_port);
   U129 : XOR2X1 port map( A => add_76_aco_carry_2_port, B => readptr_2_port, Y
                           => N335);
   U130 : AND2X1 port map( A => readptr_1_port, B => add_76_aco_carry_1_port, Y
                           => add_76_aco_carry_2_port);
   U131 : XOR2X1 port map( A => add_76_aco_carry_1_port, B => readptr_1_port, Y
                           => N334);
   U132 : AND2X1 port map( A => readptr_0_port, B => N195, Y => 
                           add_76_aco_carry_1_port);
   U133 : XOR2X1 port map( A => N195, B => readptr_0_port, Y => N333);
   U134 : NOR2X1 port map( A => n67, B => n69, Y => n87);
   U135 : AOI21X1 port map( A => n69, B => n67, C => n87, Y => n86);
   U136 : NAND2X1 port map( A => n87, B => n64, Y => n88);
   U137 : OAI21X1 port map( A => n87, B => n64, C => n88, Y => N44);
   U138 : XNOR2X1 port map( A => n71, B => n88, Y => N45);
   U139 : NOR2X1 port map( A => n71, B => n88, Y => n89);
   U140 : XOR2X1 port map( A => writeptr_4_port, B => n89, Y => N46);
   U141 : INVX2 port map( A => n86, Y => N43);
   U142 : XOR2X1 port map( A => add_67_carry_4_port, B => writeptr_4_port, Y =>
                           N51);
   U143 : MUX2X1 port map( B => n74, A => n91, S => n92, Y => n866);
   U144 : MUX2X1 port map( B => n76, A => n94, S => n92, Y => n867);
   U145 : AOI21X1 port map( A => n95, B => n96, C => n45_port, Y => n92);
   U146 : MUX2X1 port map( B => n73, A => n97, S => n98, Y => n909);
   U147 : MUX2X1 port map( B => n76, A => n99, S => n98, Y => n910);
   U148 : AOI21X1 port map( A => n96, B => n100, C => n101, Y => n98);
   U149 : MUX2X1 port map( B => n73, A => n102, S => n103, Y => n911);
   U150 : MUX2X1 port map( B => n76, A => n104, S => n103, Y => n912);
   U151 : AOI21X1 port map( A => n96, B => n105, C => n106, Y => n103);
   U152 : MUX2X1 port map( B => n73, A => n107, S => n108, Y => n913);
   U153 : MUX2X1 port map( B => n76, A => n109, S => n108, Y => n914);
   U154 : AOI21X1 port map( A => n96, B => n110, C => n111, Y => n108);
   U155 : MUX2X1 port map( B => n73, A => n112, S => n113, Y => n915);
   U156 : INVX1 port map( A => opcode_23_1_port, Y => n112);
   U157 : MUX2X1 port map( B => n76, A => n114, S => n113, Y => n916);
   U158 : AOI21X1 port map( A => n96, B => n115, C => n46_port, Y => n113);
   U159 : INVX1 port map( A => opcode_23_0_port, Y => n114);
   U160 : MUX2X1 port map( B => n73, A => n117, S => n118, Y => n917);
   U161 : INVX1 port map( A => opcode_22_1_port, Y => n117);
   U162 : MUX2X1 port map( B => n76, A => n119, S => n118, Y => n918);
   U163 : AOI21X1 port map( A => n96, B => n120, C => n121, Y => n118);
   U164 : INVX1 port map( A => opcode_22_0_port, Y => n119);
   U165 : MUX2X1 port map( B => n73, A => n122, S => n123, Y => n919);
   U166 : INVX1 port map( A => opcode_21_1_port, Y => n122);
   U167 : MUX2X1 port map( B => n76, A => n124, S => n123, Y => n920);
   U168 : AOI21X1 port map( A => n125, B => n126, C => n47, Y => n123);
   U169 : INVX1 port map( A => opcode_21_0_port, Y => n124);
   U170 : MUX2X1 port map( B => n73, A => n127, S => n128, Y => n921);
   U171 : INVX1 port map( A => opcode_20_1_port, Y => n127);
   U172 : MUX2X1 port map( B => n76, A => n129, S => n128, Y => n922);
   U173 : AOI21X1 port map( A => n130, B => n126, C => n48_port, Y => n128);
   U174 : INVX1 port map( A => opcode_20_0_port, Y => n129);
   U175 : INVX1 port map( A => n131, Y => n923);
   U176 : MUX2X1 port map( B => opcode_15_1_port, A => RCV_OPCODE(1), S => n132
                           , Y => n131);
   U177 : INVX1 port map( A => n133, Y => n924);
   U178 : MUX2X1 port map( B => opcode_15_0_port, A => RCV_OPCODE(0), S => n132
                           , Y => n133);
   U179 : OAI21X1 port map( A => n134, B => n135, C => n136, Y => n132);
   U180 : INVX1 port map( A => n137, Y => n925);
   U181 : MUX2X1 port map( B => opcode_14_1_port, A => RCV_OPCODE(1), S => n138
                           , Y => n137);
   U182 : INVX1 port map( A => n139, Y => n926);
   U183 : MUX2X1 port map( B => opcode_14_0_port, A => RCV_OPCODE(0), S => n138
                           , Y => n139);
   U184 : OAI21X1 port map( A => n140, B => n135, C => n141, Y => n138);
   U185 : MUX2X1 port map( B => n142, A => n75, S => n143, Y => n927);
   U186 : INVX1 port map( A => opcode_13_1_port, Y => n142);
   U187 : MUX2X1 port map( B => n144, A => n76, S => n143, Y => n928);
   U188 : OAI21X1 port map( A => n145, B => n146, C => n147, Y => n143);
   U189 : INVX1 port map( A => opcode_13_0_port, Y => n144);
   U190 : MUX2X1 port map( B => n148, A => n75, S => n149, Y => n929);
   U191 : INVX1 port map( A => opcode_12_1_port, Y => n148);
   U192 : MUX2X1 port map( B => n150, A => n76, S => n149, Y => n930);
   U193 : OAI21X1 port map( A => n151, B => n146, C => n152, Y => n149);
   U194 : INVX1 port map( A => opcode_12_0_port, Y => n150);
   U195 : MUX2X1 port map( B => n76, A => n153, S => n154, Y => n931);
   U196 : MUX2X1 port map( B => n73, A => n155, S => n154, Y => n932);
   U197 : AOI21X1 port map( A => n110, B => n156, C => n49_port, Y => n154);
   U198 : MUX2X1 port map( B => n76, A => n157, S => n158, Y => n933);
   U199 : MUX2X1 port map( B => n73, A => n159, S => n158, Y => n934);
   U200 : AOI21X1 port map( A => n105, B => n156, C => n50_port, Y => n158);
   U201 : MUX2X1 port map( B => n76, A => n160, S => n161, Y => n935);
   U202 : MUX2X1 port map( B => n73, A => n162, S => n161, Y => n936);
   U203 : AOI21X1 port map( A => n100, B => n156, C => n51_port, Y => n161);
   U204 : MUX2X1 port map( B => n76, A => n163, S => n164, Y => n937);
   U205 : MUX2X1 port map( B => n73, A => n165, S => n164, Y => n938);
   U206 : AOI21X1 port map( A => n95, B => n156, C => n52, Y => n164);
   U207 : MUX2X1 port map( B => n166, A => n77, S => n45_port, Y => n939);
   U208 : MUX2X1 port map( B => n167, A => n78, S => n45_port, Y => n940);
   U209 : MUX2X1 port map( B => n168, A => n79, S => n45_port, Y => n941);
   U210 : MUX2X1 port map( B => n169, A => n80, S => n45_port, Y => n942);
   U211 : MUX2X1 port map( B => n170, A => n81, S => n45_port, Y => n943);
   U212 : MUX2X1 port map( B => n171, A => n82, S => n45_port, Y => n944);
   U213 : MUX2X1 port map( B => n172, A => n83, S => n45_port, Y => n945);
   U214 : MUX2X1 port map( B => n173, A => n84, S => n45_port, Y => n946);
   U215 : MUX2X1 port map( B => n176, A => n77, S => n101, Y => n947);
   U216 : MUX2X1 port map( B => n177, A => n78, S => n101, Y => n948);
   U217 : MUX2X1 port map( B => n178, A => n79, S => n101, Y => n949);
   U218 : MUX2X1 port map( B => n179, A => n80, S => n101, Y => n950);
   U219 : MUX2X1 port map( B => n180, A => n81, S => n101, Y => n951);
   U220 : MUX2X1 port map( B => n181, A => n82, S => n101, Y => n952);
   U221 : MUX2X1 port map( B => n182, A => n83, S => n101, Y => n953);
   U222 : MUX2X1 port map( B => n183, A => n84, S => n101, Y => n954);
   U223 : MUX2X1 port map( B => n185, A => n77, S => n106, Y => n955);
   U224 : MUX2X1 port map( B => n186, A => n78, S => n106, Y => n956);
   U225 : MUX2X1 port map( B => n187, A => n79, S => n106, Y => n957);
   U226 : MUX2X1 port map( B => n188, A => n80, S => n106, Y => n958);
   U227 : MUX2X1 port map( B => n189_port, A => n81, S => n106, Y => n959);
   U228 : MUX2X1 port map( B => n190_port, A => n82, S => n106, Y => n960);
   U229 : MUX2X1 port map( B => n191_port, A => n83, S => n106, Y => n961);
   U230 : MUX2X1 port map( B => n192_port, A => n84, S => n106, Y => n962);
   U231 : MUX2X1 port map( B => n193_port, A => n77, S => n111, Y => n963);
   U232 : MUX2X1 port map( B => n194, A => n78, S => n111, Y => n964);
   U233 : MUX2X1 port map( B => n195_port, A => n79, S => n111, Y => n965);
   U234 : MUX2X1 port map( B => n196, A => n80, S => n111, Y => n966);
   U235 : MUX2X1 port map( B => n197, A => n81, S => n111, Y => n967);
   U236 : MUX2X1 port map( B => n198, A => n82, S => n111, Y => n968);
   U237 : MUX2X1 port map( B => n199, A => n83, S => n111, Y => n969);
   U238 : MUX2X1 port map( B => n200, A => n84, S => n111, Y => n970);
   U239 : MUX2X1 port map( B => n201, A => n77, S => n46_port, Y => n971);
   U240 : INVX1 port map( A => memory_23_7_port, Y => n201);
   U241 : MUX2X1 port map( B => n202, A => n78, S => n46_port, Y => n972);
   U242 : INVX1 port map( A => memory_23_6_port, Y => n202);
   U243 : MUX2X1 port map( B => n203, A => n79, S => n46_port, Y => n973);
   U244 : INVX1 port map( A => memory_23_5_port, Y => n203);
   U245 : MUX2X1 port map( B => n204, A => n80, S => n46_port, Y => n974);
   U246 : INVX1 port map( A => memory_23_4_port, Y => n204);
   U247 : MUX2X1 port map( B => n205, A => n81, S => n46_port, Y => n975);
   U248 : INVX1 port map( A => memory_23_3_port, Y => n205);
   U249 : MUX2X1 port map( B => n206, A => n82, S => n46_port, Y => n976);
   U250 : INVX1 port map( A => memory_23_2_port, Y => n206);
   U251 : MUX2X1 port map( B => n207, A => n83, S => n46_port, Y => n977);
   U252 : INVX1 port map( A => memory_23_1_port, Y => n207);
   U253 : MUX2X1 port map( B => n208, A => n84, S => n46_port, Y => n978);
   U254 : NOR2X1 port map( A => n145, B => n209, Y => n116);
   U255 : INVX1 port map( A => memory_23_0_port, Y => n208);
   U256 : MUX2X1 port map( B => n210, A => n77, S => n121, Y => n979);
   U257 : INVX1 port map( A => memory_22_7_port, Y => n210);
   U258 : MUX2X1 port map( B => n211, A => n78, S => n121, Y => n980);
   U259 : INVX1 port map( A => memory_22_6_port, Y => n211);
   U260 : MUX2X1 port map( B => n212, A => n79, S => n121, Y => n981);
   U261 : INVX1 port map( A => memory_22_5_port, Y => n212);
   U262 : MUX2X1 port map( B => n213, A => n80, S => n121, Y => n982);
   U263 : INVX1 port map( A => memory_22_4_port, Y => n213);
   U264 : MUX2X1 port map( B => n214, A => n81, S => n121, Y => n983);
   U265 : INVX1 port map( A => memory_22_3_port, Y => n214);
   U266 : MUX2X1 port map( B => n215, A => n82, S => n121, Y => n984);
   U267 : INVX1 port map( A => memory_22_2_port, Y => n215);
   U268 : MUX2X1 port map( B => n216, A => n83, S => n121, Y => n985);
   U269 : INVX1 port map( A => memory_22_1_port, Y => n216);
   U270 : MUX2X1 port map( B => n217, A => n84, S => n121, Y => n986);
   U271 : INVX1 port map( A => memory_22_0_port, Y => n217);
   U272 : MUX2X1 port map( B => n218, A => n77, S => n47, Y => n987);
   U273 : INVX1 port map( A => memory_21_7_port, Y => n218);
   U274 : MUX2X1 port map( B => n219, A => n78, S => n47, Y => n988);
   U275 : INVX1 port map( A => memory_21_6_port, Y => n219);
   U276 : MUX2X1 port map( B => n220, A => n79, S => n47, Y => n989);
   U277 : INVX1 port map( A => memory_21_5_port, Y => n220);
   U278 : MUX2X1 port map( B => n221, A => n80, S => n47, Y => n990);
   U279 : INVX1 port map( A => memory_21_4_port, Y => n221);
   U280 : MUX2X1 port map( B => n222, A => n81, S => n47, Y => n991);
   U281 : INVX1 port map( A => memory_21_3_port, Y => n222);
   U282 : MUX2X1 port map( B => n223, A => n82, S => n47, Y => n992);
   U283 : INVX1 port map( A => memory_21_2_port, Y => n223);
   U284 : MUX2X1 port map( B => n224, A => n83, S => n47, Y => n993);
   U285 : INVX1 port map( A => memory_21_1_port, Y => n224);
   U286 : MUX2X1 port map( B => n225, A => n84, S => n47, Y => n994);
   U287 : INVX1 port map( A => memory_21_0_port, Y => n225);
   U288 : MUX2X1 port map( B => n227, A => n77, S => n48_port, Y => n995);
   U289 : INVX1 port map( A => memory_20_7_port, Y => n227);
   U290 : MUX2X1 port map( B => n228, A => n78, S => n48_port, Y => n996);
   U291 : INVX1 port map( A => memory_20_6_port, Y => n228);
   U292 : MUX2X1 port map( B => n229, A => n79, S => n48_port, Y => n997);
   U293 : INVX1 port map( A => memory_20_5_port, Y => n229);
   U294 : MUX2X1 port map( B => n230, A => n80, S => n48_port, Y => n998);
   U295 : INVX1 port map( A => memory_20_4_port, Y => n230);
   U296 : MUX2X1 port map( B => n231, A => n81, S => n48_port, Y => n999);
   U297 : INVX1 port map( A => memory_20_3_port, Y => n231);
   U298 : MUX2X1 port map( B => n232, A => n82, S => n48_port, Y => n1000);
   U299 : INVX1 port map( A => memory_20_2_port, Y => n232);
   U300 : MUX2X1 port map( B => n233, A => n83, S => n48_port, Y => n1001);
   U301 : INVX1 port map( A => memory_20_1_port, Y => n233);
   U302 : MUX2X1 port map( B => n234, A => n84, S => n48_port, Y => n1002);
   U303 : INVX1 port map( A => memory_20_0_port, Y => n234);
   U304 : MUX2X1 port map( B => n77, A => n236, S => n136, Y => n1003);
   U305 : INVX1 port map( A => memory_15_7_port, Y => n236);
   U306 : MUX2X1 port map( B => n78, A => n237, S => n136, Y => n1004);
   U307 : INVX1 port map( A => memory_15_6_port, Y => n237);
   U308 : MUX2X1 port map( B => n79, A => n238, S => n136, Y => n1005);
   U309 : INVX1 port map( A => memory_15_5_port, Y => n238);
   U310 : MUX2X1 port map( B => n80, A => n239, S => n136, Y => n1006);
   U311 : INVX1 port map( A => memory_15_4_port, Y => n239);
   U312 : MUX2X1 port map( B => n81, A => n240, S => n136, Y => n1007);
   U313 : INVX1 port map( A => memory_15_3_port, Y => n240);
   U314 : MUX2X1 port map( B => n82, A => n241, S => n136, Y => n1008);
   U315 : INVX1 port map( A => memory_15_2_port, Y => n241);
   U316 : MUX2X1 port map( B => n83, A => n242, S => n136, Y => n1009);
   U317 : INVX1 port map( A => memory_15_1_port, Y => n242);
   U318 : MUX2X1 port map( B => n84, A => n243, S => n136, Y => n1010);
   U319 : NAND2X1 port map( A => n244, B => n125, Y => n136);
   U320 : INVX1 port map( A => memory_15_0_port, Y => n243);
   U321 : MUX2X1 port map( B => n77, A => n245, S => n141, Y => n1011);
   U322 : INVX1 port map( A => memory_14_7_port, Y => n245);
   U323 : MUX2X1 port map( B => n78, A => n246, S => n141, Y => n1012);
   U324 : INVX1 port map( A => memory_14_6_port, Y => n246);
   U325 : MUX2X1 port map( B => n79, A => n247, S => n141, Y => n1013);
   U326 : INVX1 port map( A => memory_14_5_port, Y => n247);
   U327 : MUX2X1 port map( B => n80, A => n248, S => n141, Y => n1014);
   U328 : INVX1 port map( A => memory_14_4_port, Y => n248);
   U329 : MUX2X1 port map( B => n81, A => n249, S => n141, Y => n1015);
   U330 : INVX1 port map( A => memory_14_3_port, Y => n249);
   U331 : MUX2X1 port map( B => n82, A => n250, S => n141, Y => n1016);
   U332 : INVX1 port map( A => memory_14_2_port, Y => n250);
   U333 : MUX2X1 port map( B => n83, A => n251, S => n141, Y => n1017);
   U334 : INVX1 port map( A => memory_14_1_port, Y => n251);
   U335 : MUX2X1 port map( B => n84, A => n252, S => n141, Y => n1018);
   U336 : NAND2X1 port map( A => n244, B => n130, Y => n141);
   U337 : INVX1 port map( A => memory_14_0_port, Y => n252);
   U338 : MUX2X1 port map( B => n77, A => n253, S => n147, Y => n1019);
   U339 : INVX1 port map( A => memory_13_7_port, Y => n253);
   U340 : MUX2X1 port map( B => n78, A => n254, S => n147, Y => n1020);
   U341 : INVX1 port map( A => memory_13_6_port, Y => n254);
   U342 : MUX2X1 port map( B => n79, A => n255, S => n147, Y => n1021);
   U343 : INVX1 port map( A => memory_13_5_port, Y => n255);
   U344 : MUX2X1 port map( B => n80, A => n256, S => n147, Y => n1022);
   U345 : INVX1 port map( A => memory_13_4_port, Y => n256);
   U346 : MUX2X1 port map( B => n81, A => n257, S => n147, Y => n1023);
   U347 : INVX1 port map( A => memory_13_3_port, Y => n257);
   U348 : MUX2X1 port map( B => n82, A => n258, S => n147, Y => n1024);
   U349 : INVX1 port map( A => memory_13_2_port, Y => n258);
   U350 : MUX2X1 port map( B => n83, A => n259, S => n147, Y => n1025);
   U351 : INVX1 port map( A => memory_13_1_port, Y => n259);
   U352 : MUX2X1 port map( B => n84, A => n260, S => n147, Y => n1026);
   U353 : NAND2X1 port map( A => n244, B => n95, Y => n147);
   U354 : INVX1 port map( A => memory_13_0_port, Y => n260);
   U355 : MUX2X1 port map( B => n77, A => n261, S => n152, Y => n1027);
   U356 : INVX1 port map( A => memory_12_7_port, Y => n261);
   U357 : MUX2X1 port map( B => n78, A => n262, S => n152, Y => n1028);
   U358 : INVX1 port map( A => memory_12_6_port, Y => n262);
   U359 : MUX2X1 port map( B => n79, A => n263, S => n152, Y => n1029);
   U360 : INVX1 port map( A => memory_12_5_port, Y => n263);
   U361 : MUX2X1 port map( B => n80, A => n264, S => n152, Y => n1064);
   U362 : INVX1 port map( A => memory_12_4_port, Y => n264);
   U363 : MUX2X1 port map( B => n81, A => n265, S => n152, Y => n1065);
   U364 : INVX1 port map( A => memory_12_3_port, Y => n265);
   U365 : MUX2X1 port map( B => n82, A => n266, S => n152, Y => n1066);
   U366 : INVX1 port map( A => memory_12_2_port, Y => n266);
   U367 : MUX2X1 port map( B => n83, A => n267, S => n152, Y => n1067);
   U368 : INVX1 port map( A => memory_12_1_port, Y => n267);
   U369 : MUX2X1 port map( B => n84, A => n268, S => n152, Y => n1068);
   U370 : NAND2X1 port map( A => n244, B => n100, Y => n152);
   U371 : INVX1 port map( A => memory_12_0_port, Y => n268);
   U372 : MUX2X1 port map( B => n269, A => n84, S => n49_port, Y => n1069);
   U373 : MUX2X1 port map( B => n270, A => n83, S => n49_port, Y => n1070);
   U374 : MUX2X1 port map( B => n271, A => n82, S => n49_port, Y => n1071);
   U375 : MUX2X1 port map( B => n272, A => n81, S => n49_port, Y => n1168);
   U376 : MUX2X1 port map( B => n273, A => n80, S => n49_port, Y => n1169);
   U377 : MUX2X1 port map( B => n274, A => n79, S => n49_port, Y => n1170);
   U378 : MUX2X1 port map( B => n275, A => n78, S => n49_port, Y => n1171);
   U379 : MUX2X1 port map( B => n276, A => n77, S => n49_port, Y => n1172);
   U380 : MUX2X1 port map( B => n278, A => n84, S => n50_port, Y => n1173);
   U381 : MUX2X1 port map( B => n279, A => n83, S => n50_port, Y => n1174);
   U382 : MUX2X1 port map( B => n280, A => n82, S => n50_port, Y => n1175);
   U383 : MUX2X1 port map( B => n281, A => n81, S => n50_port, Y => n1176);
   U384 : MUX2X1 port map( B => n282, A => n80, S => n50_port, Y => n1177);
   U385 : MUX2X1 port map( B => n283, A => n79, S => n50_port, Y => n1178);
   U386 : MUX2X1 port map( B => n284, A => n78, S => n50_port, Y => n1179);
   U387 : MUX2X1 port map( B => n285, A => n77, S => n50_port, Y => n1180);
   U388 : MUX2X1 port map( B => n286, A => n84, S => n51_port, Y => n1181);
   U389 : MUX2X1 port map( B => n287, A => n83, S => n51_port, Y => n1182);
   U390 : MUX2X1 port map( B => n288, A => n82, S => n51_port, Y => n1183);
   U391 : MUX2X1 port map( B => n289, A => n81, S => n51_port, Y => n1184);
   U392 : MUX2X1 port map( B => n290, A => n80, S => n51_port, Y => n1185);
   U393 : MUX2X1 port map( B => n291, A => n79, S => n51_port, Y => n1186);
   U394 : MUX2X1 port map( B => n292, A => n78, S => n51_port, Y => n1187);
   U395 : MUX2X1 port map( B => n293, A => n77, S => n51_port, Y => n1188);
   U396 : MUX2X1 port map( B => n294, A => n84, S => n52, Y => n1189);
   U397 : MUX2X1 port map( B => n295, A => n83, S => n52, Y => n1190);
   U398 : MUX2X1 port map( B => n296, A => n82, S => n52, Y => n1191);
   U399 : MUX2X1 port map( B => n297, A => n81, S => n52, Y => n1192);
   U400 : MUX2X1 port map( B => n298, A => n80, S => n52, Y => n1193);
   U401 : MUX2X1 port map( B => n299, A => n79, S => n52, Y => n1194);
   U402 : MUX2X1 port map( B => n300, A => n78, S => n52, Y => n1195);
   U403 : MUX2X1 port map( B => n301, A => n77, S => n52, Y => n1196);
   U404 : MUX2X1 port map( B => n302, A => n303, S => RST, Y => n1197);
   U405 : INVX1 port map( A => FULL_port, Y => n303);
   U406 : MUX2X1 port map( B => n304, A => n305, S => RST, Y => n1198);
   U407 : INVX1 port map( A => EMPTY_port, Y => n305);
   U408 : MUX2X1 port map( B => n76, A => n306, S => n307, Y => n908);
   U409 : INVX1 port map( A => opcode_7_0_port, Y => n306);
   U410 : MUX2X1 port map( B => n73, A => n308, S => n307, Y => n907);
   U411 : AOI21X1 port map( A => n115, B => n309, C => n53, Y => n307);
   U412 : INVX1 port map( A => opcode_7_1_port, Y => n308);
   U413 : MUX2X1 port map( B => n310, A => n84, S => n53, Y => n906);
   U414 : INVX1 port map( A => memory_7_0_port, Y => n310);
   U415 : MUX2X1 port map( B => n311, A => n83, S => n53, Y => n905);
   U416 : INVX1 port map( A => memory_7_1_port, Y => n311);
   U417 : MUX2X1 port map( B => n312, A => n82, S => n53, Y => n904);
   U418 : INVX1 port map( A => memory_7_2_port, Y => n312);
   U419 : MUX2X1 port map( B => n313, A => n81, S => n53, Y => n903);
   U420 : INVX1 port map( A => memory_7_3_port, Y => n313);
   U421 : MUX2X1 port map( B => n314, A => n80, S => n53, Y => n902);
   U422 : INVX1 port map( A => memory_7_4_port, Y => n314);
   U423 : MUX2X1 port map( B => n315, A => n79, S => n53, Y => n901);
   U424 : INVX1 port map( A => memory_7_5_port, Y => n315);
   U425 : MUX2X1 port map( B => n316, A => n78, S => n53, Y => n900);
   U426 : INVX1 port map( A => memory_7_6_port, Y => n316);
   U427 : MUX2X1 port map( B => n317, A => n77, S => n53, Y => n899);
   U428 : INVX1 port map( A => memory_7_7_port, Y => n317);
   U429 : MUX2X1 port map( B => n76, A => n318, S => n319, Y => n898);
   U430 : INVX1 port map( A => opcode_6_0_port, Y => n318);
   U431 : MUX2X1 port map( B => n74, A => n320, S => n319, Y => n897);
   U432 : AOI21X1 port map( A => n120, B => n309, C => n54, Y => n319);
   U433 : INVX1 port map( A => opcode_6_1_port, Y => n320);
   U434 : MUX2X1 port map( B => n321, A => n84, S => n54, Y => n896);
   U435 : INVX1 port map( A => memory_6_0_port, Y => n321);
   U436 : MUX2X1 port map( B => n322, A => n83, S => n54, Y => n895);
   U437 : INVX1 port map( A => memory_6_1_port, Y => n322);
   U438 : MUX2X1 port map( B => n323, A => n82, S => n54, Y => n894);
   U439 : INVX1 port map( A => memory_6_2_port, Y => n323);
   U440 : MUX2X1 port map( B => n324, A => n81, S => n54, Y => n893);
   U441 : INVX1 port map( A => memory_6_3_port, Y => n324);
   U442 : MUX2X1 port map( B => n325, A => n80, S => n54, Y => n892);
   U443 : INVX1 port map( A => memory_6_4_port, Y => n325);
   U444 : MUX2X1 port map( B => n326, A => n79, S => n54, Y => n891);
   U445 : INVX1 port map( A => memory_6_5_port, Y => n326);
   U446 : MUX2X1 port map( B => n327, A => n78, S => n54, Y => n890);
   U447 : INVX1 port map( A => memory_6_6_port, Y => n327);
   U448 : MUX2X1 port map( B => n328, A => n77, S => n54, Y => n889);
   U449 : INVX1 port map( A => memory_6_7_port, Y => n328);
   U450 : MUX2X1 port map( B => n93, A => n329, S => n330, Y => n888);
   U451 : INVX1 port map( A => opcode_5_0_port, Y => n329);
   U452 : MUX2X1 port map( B => n74, A => n331, S => n330, Y => n887);
   U453 : AOI21X1 port map( A => n125, B => n156, C => n55, Y => n330);
   U454 : INVX1 port map( A => opcode_5_1_port, Y => n331);
   U455 : MUX2X1 port map( B => n332, A => n84, S => n55, Y => n886);
   U456 : INVX1 port map( A => memory_5_0_port, Y => n332);
   U457 : MUX2X1 port map( B => n333_port, A => n83, S => n55, Y => n885);
   U458 : INVX1 port map( A => memory_5_1_port, Y => n333_port);
   U459 : MUX2X1 port map( B => n334_port, A => n82, S => n55, Y => n884);
   U460 : INVX1 port map( A => memory_5_2_port, Y => n334_port);
   U461 : MUX2X1 port map( B => n335_port, A => n81, S => n55, Y => n883);
   U462 : INVX1 port map( A => memory_5_3_port, Y => n335_port);
   U463 : MUX2X1 port map( B => n336_port, A => n80, S => n55, Y => n882);
   U464 : INVX1 port map( A => memory_5_4_port, Y => n336_port);
   U465 : MUX2X1 port map( B => n337_port, A => n79, S => n55, Y => n881);
   U466 : INVX1 port map( A => memory_5_5_port, Y => n337_port);
   U467 : MUX2X1 port map( B => n338_port, A => n78, S => n55, Y => n880);
   U468 : INVX1 port map( A => memory_5_6_port, Y => n338_port);
   U469 : MUX2X1 port map( B => n339_port, A => n77, S => n55, Y => n879);
   U470 : INVX1 port map( A => memory_5_7_port, Y => n339_port);
   U471 : MUX2X1 port map( B => n76, A => n340_port, S => n341_port, Y => n878)
                           ;
   U472 : INVX1 port map( A => opcode_4_0_port, Y => n340_port);
   U473 : MUX2X1 port map( B => n74, A => n342_port, S => n341_port, Y => n877)
                           ;
   U474 : AOI21X1 port map( A => n130, B => n156, C => n56, Y => n341_port);
   U475 : INVX1 port map( A => opcode_4_1_port, Y => n342_port);
   U476 : MUX2X1 port map( B => n343_port, A => n84, S => n56, Y => n876);
   U477 : INVX1 port map( A => memory_4_0_port, Y => n343_port);
   U478 : MUX2X1 port map( B => n344_port, A => n83, S => n56, Y => n875);
   U479 : INVX1 port map( A => memory_4_1_port, Y => n344_port);
   U480 : MUX2X1 port map( B => n345_port, A => n82, S => n56, Y => n874);
   U481 : INVX1 port map( A => memory_4_2_port, Y => n345_port);
   U482 : MUX2X1 port map( B => n346_port, A => n81, S => n56, Y => n873);
   U483 : INVX1 port map( A => memory_4_3_port, Y => n346_port);
   U484 : MUX2X1 port map( B => n347_port, A => n80, S => n56, Y => n872);
   U485 : INVX1 port map( A => memory_4_4_port, Y => n347_port);
   U486 : MUX2X1 port map( B => n348, A => n79, S => n56, Y => n871);
   U487 : INVX1 port map( A => memory_4_5_port, Y => n348);
   U488 : MUX2X1 port map( B => n349, A => n78, S => n56, Y => n870);
   U489 : INVX1 port map( A => memory_4_6_port, Y => n349);
   U490 : MUX2X1 port map( B => n350, A => n77, S => n56, Y => n869);
   U491 : NAND3X1 port map( A => n63, B => n70, C => n352, Y => n277);
   U492 : INVX1 port map( A => memory_4_7_port, Y => n350);
   U493 : OAI21X1 port map( A => n353, B => n354, C => n355, Y => n862);
   U494 : AOI22X1 port map( A => N51, B => n44_port, C => N46, D => n356, Y => 
                           n355);
   U495 : OAI21X1 port map( A => n353, B => n70, C => n357, Y => n860);
   U496 : AOI22X1 port map( A => N50, B => n44_port, C => N45, D => n356, Y => 
                           n357);
   U497 : OAI21X1 port map( A => n353, B => n358, C => n359, Y => n858);
   U498 : AOI22X1 port map( A => n358, B => n44_port, C => n358, D => n356, Y 
                           => n359);
   U499 : OAI21X1 port map( A => n353, B => n360, C => n361, Y => n856);
   U500 : AOI22X1 port map( A => N48, B => n44_port, C => N43, D => n356, Y => 
                           n361);
   U501 : OAI21X1 port map( A => n353, B => n64, C => n362, Y => n854);
   U502 : AOI22X1 port map( A => N49, B => n44_port, C => N44, D => n356, Y => 
                           n362);
   U503 : MUX2X1 port map( B => n77, A => n363, S => n364, Y => n1167);
   U504 : MUX2X1 port map( B => n78, A => n365, S => n364, Y => n1166);
   U505 : MUX2X1 port map( B => n79, A => n366, S => n364, Y => n1165);
   U506 : MUX2X1 port map( B => n80, A => n367, S => n364, Y => n1164);
   U507 : MUX2X1 port map( B => n81, A => n368, S => n364, Y => n1163);
   U508 : MUX2X1 port map( B => n82, A => n369, S => n364, Y => n1162);
   U509 : MUX2X1 port map( B => n83, A => n370, S => n364, Y => n1161);
   U510 : MUX2X1 port map( B => n84, A => n371, S => n364, Y => n1160);
   U511 : MUX2X1 port map( B => n77, A => n372, S => n373, Y => n1159);
   U512 : MUX2X1 port map( B => n78, A => n374, S => n373, Y => n1158);
   U513 : MUX2X1 port map( B => n79, A => n375, S => n373, Y => n1157);
   U514 : MUX2X1 port map( B => n80, A => n376, S => n373, Y => n1156);
   U515 : MUX2X1 port map( B => n81, A => n377, S => n373, Y => n1155);
   U516 : MUX2X1 port map( B => n82, A => n378, S => n373, Y => n1154);
   U517 : MUX2X1 port map( B => n83, A => n379, S => n373, Y => n1153);
   U518 : MUX2X1 port map( B => n84, A => n380, S => n373, Y => n1152);
   U519 : MUX2X1 port map( B => n77, A => n381, S => n382, Y => n1151);
   U520 : MUX2X1 port map( B => n78, A => n383, S => n382, Y => n1150);
   U521 : MUX2X1 port map( B => n79, A => n384, S => n382, Y => n1149);
   U522 : MUX2X1 port map( B => n80, A => n385, S => n382, Y => n1148);
   U523 : MUX2X1 port map( B => n81, A => n386, S => n382, Y => n1147);
   U524 : MUX2X1 port map( B => n82, A => n387, S => n382, Y => n1146);
   U525 : MUX2X1 port map( B => n83, A => n388, S => n382, Y => n1145);
   U526 : MUX2X1 port map( B => n84, A => n389, S => n382, Y => n1144);
   U527 : MUX2X1 port map( B => n390, A => n77, S => n391, Y => n1143);
   U528 : MUX2X1 port map( B => n392, A => n78, S => n391, Y => n1142);
   U529 : MUX2X1 port map( B => n393, A => n79, S => n391, Y => n1141);
   U530 : MUX2X1 port map( B => n394, A => n80, S => n391, Y => n1140);
   U531 : MUX2X1 port map( B => n395, A => n81, S => n391, Y => n1139);
   U532 : MUX2X1 port map( B => n396, A => n82, S => n391, Y => n1138);
   U533 : MUX2X1 port map( B => n397, A => n83, S => n391, Y => n1137);
   U534 : MUX2X1 port map( B => n398, A => n84, S => n391, Y => n1136);
   U535 : AND2X1 port map( A => n244, B => n105, Y => n391);
   U536 : MUX2X1 port map( B => n399, A => n77, S => n57, Y => n1135);
   U537 : MUX2X1 port map( B => n400, A => n78, S => n57, Y => n1134);
   U538 : MUX2X1 port map( B => n401, A => n79, S => n57, Y => n1133);
   U539 : MUX2X1 port map( B => n402, A => n80, S => n57, Y => n1132);
   U540 : MUX2X1 port map( B => n403, A => n81, S => n57, Y => n1131);
   U541 : MUX2X1 port map( B => n404, A => n82, S => n57, Y => n1130);
   U542 : MUX2X1 port map( B => n405, A => n83, S => n57, Y => n1129);
   U543 : MUX2X1 port map( B => n406, A => n84, S => n57, Y => n1128);
   U544 : MUX2X1 port map( B => n407, A => n77, S => n58, Y => n1127);
   U545 : MUX2X1 port map( B => n408, A => n78, S => n58, Y => n1126);
   U546 : MUX2X1 port map( B => n409, A => n79, S => n58, Y => n1125);
   U547 : MUX2X1 port map( B => n410, A => n80, S => n58, Y => n1124);
   U548 : MUX2X1 port map( B => n411, A => n81, S => n58, Y => n1123);
   U549 : MUX2X1 port map( B => n412, A => n82, S => n58, Y => n1122);
   U550 : MUX2X1 port map( B => n413, A => n83, S => n58, Y => n1121);
   U551 : MUX2X1 port map( B => n414, A => n84, S => n58, Y => n1120);
   U552 : MUX2X1 port map( B => n415, A => n77, S => n59, Y => n1119);
   U553 : MUX2X1 port map( B => n416, A => n78, S => n59, Y => n1118);
   U554 : MUX2X1 port map( B => n417, A => n79, S => n59, Y => n1117);
   U555 : MUX2X1 port map( B => n418, A => n80, S => n59, Y => n1116);
   U556 : MUX2X1 port map( B => n419, A => n81, S => n59, Y => n1115);
   U557 : MUX2X1 port map( B => n420, A => n82, S => n59, Y => n1114);
   U558 : MUX2X1 port map( B => n421, A => n83, S => n59, Y => n1113);
   U559 : MUX2X1 port map( B => n422, A => n84, S => n59, Y => n1112);
   U560 : MUX2X1 port map( B => n423, A => n77, S => n60, Y => n1111);
   U561 : MUX2X1 port map( B => n424, A => n78, S => n60, Y => n1110);
   U562 : MUX2X1 port map( B => n425, A => n79, S => n60, Y => n1109);
   U563 : MUX2X1 port map( B => n426, A => n80, S => n60, Y => n1108);
   U564 : MUX2X1 port map( B => n427, A => n81, S => n60, Y => n1107);
   U565 : MUX2X1 port map( B => n428, A => n82, S => n60, Y => n1106);
   U566 : MUX2X1 port map( B => n429, A => n83, S => n60, Y => n1105);
   U567 : MUX2X1 port map( B => n430, A => n84, S => n60, Y => n1104);
   U568 : INVX1 port map( A => n431, Y => n1103);
   U569 : MUX2X1 port map( B => memory_28_7_port, A => RCV_DATA(7), S => n432, 
                           Y => n431);
   U570 : INVX1 port map( A => n433, Y => n1102);
   U571 : MUX2X1 port map( B => memory_28_6_port, A => RCV_DATA(6), S => n432, 
                           Y => n433);
   U572 : INVX1 port map( A => n434, Y => n1101);
   U573 : MUX2X1 port map( B => memory_28_5_port, A => RCV_DATA(5), S => n432, 
                           Y => n434);
   U574 : INVX1 port map( A => n435, Y => n1100);
   U575 : MUX2X1 port map( B => memory_28_4_port, A => RCV_DATA(4), S => n432, 
                           Y => n435);
   U576 : INVX1 port map( A => n436, Y => n1099);
   U577 : MUX2X1 port map( B => memory_28_3_port, A => RCV_DATA(3), S => n432, 
                           Y => n436);
   U578 : INVX1 port map( A => n437, Y => n1098);
   U579 : MUX2X1 port map( B => memory_28_2_port, A => RCV_DATA(2), S => n432, 
                           Y => n437);
   U580 : INVX1 port map( A => n438, Y => n1097);
   U581 : MUX2X1 port map( B => memory_28_1_port, A => RCV_DATA(1), S => n432, 
                           Y => n438);
   U582 : INVX1 port map( A => n439, Y => n1096);
   U583 : MUX2X1 port map( B => memory_28_0_port, A => RCV_DATA(0), S => n432, 
                           Y => n439);
   U584 : INVX1 port map( A => n440, Y => n1095);
   U585 : MUX2X1 port map( B => memory_29_7_port, A => RCV_DATA(7), S => n61, Y
                           => n440);
   U586 : INVX1 port map( A => n441, Y => n1094);
   U587 : MUX2X1 port map( B => memory_29_6_port, A => RCV_DATA(6), S => n61, Y
                           => n441);
   U588 : INVX1 port map( A => n442, Y => n1093);
   U589 : MUX2X1 port map( B => memory_29_5_port, A => RCV_DATA(5), S => n61, Y
                           => n442);
   U590 : INVX1 port map( A => n443, Y => n1092);
   U591 : MUX2X1 port map( B => memory_29_4_port, A => RCV_DATA(4), S => n61, Y
                           => n443);
   U592 : INVX1 port map( A => n444, Y => n1091);
   U593 : MUX2X1 port map( B => memory_29_3_port, A => RCV_DATA(3), S => n61, Y
                           => n444);
   U594 : INVX1 port map( A => n445, Y => n1090);
   U595 : MUX2X1 port map( B => memory_29_2_port, A => RCV_DATA(2), S => n61, Y
                           => n445);
   U596 : INVX1 port map( A => n446, Y => n1089);
   U597 : MUX2X1 port map( B => memory_29_1_port, A => RCV_DATA(1), S => n61, Y
                           => n446);
   U598 : INVX1 port map( A => n447, Y => n1088);
   U599 : MUX2X1 port map( B => memory_29_0_port, A => RCV_DATA(0), S => n61, Y
                           => n447);
   U600 : INVX1 port map( A => n448, Y => n1087);
   U601 : MUX2X1 port map( B => memory_30_7_port, A => RCV_DATA(7), S => n62, Y
                           => n448);
   U602 : INVX1 port map( A => n450, Y => n1086);
   U603 : MUX2X1 port map( B => memory_30_6_port, A => RCV_DATA(6), S => n62, Y
                           => n450);
   U604 : INVX1 port map( A => n451, Y => n1085);
   U605 : MUX2X1 port map( B => memory_30_5_port, A => RCV_DATA(5), S => n62, Y
                           => n451);
   U606 : INVX1 port map( A => n452, Y => n1084);
   U607 : MUX2X1 port map( B => memory_30_4_port, A => RCV_DATA(4), S => n62, Y
                           => n452);
   U608 : INVX1 port map( A => n453, Y => n1083);
   U609 : MUX2X1 port map( B => memory_30_3_port, A => RCV_DATA(3), S => n62, Y
                           => n453);
   U610 : INVX1 port map( A => n454, Y => n1082);
   U611 : MUX2X1 port map( B => memory_30_2_port, A => RCV_DATA(2), S => n62, Y
                           => n454);
   U612 : INVX1 port map( A => n455, Y => n1081);
   U613 : MUX2X1 port map( B => memory_30_1_port, A => RCV_DATA(1), S => n62, Y
                           => n455);
   U614 : INVX1 port map( A => n456, Y => n1080);
   U615 : MUX2X1 port map( B => memory_30_0_port, A => RCV_DATA(0), S => n62, Y
                           => n456);
   U616 : INVX1 port map( A => n457, Y => n1079);
   U617 : MUX2X1 port map( B => memory_31_7_port, A => RCV_DATA(7), S => n458, 
                           Y => n457);
   U618 : INVX1 port map( A => n459, Y => n1078);
   U619 : MUX2X1 port map( B => memory_31_6_port, A => RCV_DATA(6), S => n458, 
                           Y => n459);
   U620 : INVX1 port map( A => n460, Y => n1077);
   U621 : MUX2X1 port map( B => memory_31_5_port, A => RCV_DATA(5), S => n458, 
                           Y => n460);
   U622 : INVX1 port map( A => n461, Y => n1076);
   U623 : MUX2X1 port map( B => memory_31_4_port, A => RCV_DATA(4), S => n458, 
                           Y => n461);
   U624 : INVX1 port map( A => n462, Y => n1075);
   U625 : MUX2X1 port map( B => memory_31_3_port, A => RCV_DATA(3), S => n458, 
                           Y => n462);
   U626 : INVX1 port map( A => n463, Y => n1074);
   U627 : MUX2X1 port map( B => memory_31_2_port, A => RCV_DATA(2), S => n458, 
                           Y => n463);
   U628 : INVX1 port map( A => n464, Y => n1073);
   U629 : MUX2X1 port map( B => memory_31_1_port, A => RCV_DATA(1), S => n458, 
                           Y => n464);
   U630 : INVX1 port map( A => n465, Y => n1072);
   U631 : MUX2X1 port map( B => memory_31_0_port, A => RCV_DATA(0), S => n458, 
                           Y => n465);
   U632 : MUX2X1 port map( B => n466, A => n75, S => n467, Y => n1063);
   U633 : MUX2X1 port map( B => n468, A => n76, S => n467, Y => n1062);
   U634 : OAI21X1 port map( A => n184, B => n146, C => n364, Y => n467);
   U635 : NAND2X1 port map( A => n244, B => n120, Y => n364);
   U636 : MUX2X1 port map( B => n469, A => n75, S => n470, Y => n1061);
   U637 : MUX2X1 port map( B => n471, A => n76, S => n470, Y => n1060);
   U638 : OAI21X1 port map( A => n175, B => n146, C => n373, Y => n470);
   U639 : NAND2X1 port map( A => n244, B => n115, Y => n373);
   U640 : MUX2X1 port map( B => n472, A => n75, S => n473, Y => n1059);
   U641 : MUX2X1 port map( B => n474, A => n76, S => n473, Y => n1058);
   U642 : OAI21X1 port map( A => n235, B => n146, C => n382, Y => n473);
   U643 : NAND2X1 port map( A => n244, B => n110, Y => n382);
   U644 : NAND2X1 port map( A => n475, B => n356, Y => n146);
   U645 : MUX2X1 port map( B => n74, A => n476, S => n477, Y => n1057);
   U646 : MUX2X1 port map( B => n76, A => n478, S => n477, Y => n1056);
   U647 : NAND3X1 port map( A => n475, B => n353, C => n479, Y => n477);
   U648 : MUX2X1 port map( B => n175, A => n226, S => n480, Y => n479);
   U649 : AND2X1 port map( A => n352, B => n71, Y => n475);
   U650 : MUX2X1 port map( B => n74, A => n481, S => n482, Y => n1055);
   U651 : MUX2X1 port map( B => n76, A => n483, S => n482, Y => n1054);
   U652 : AOI21X1 port map( A => n110, B => n126, C => n57, Y => n482);
   U653 : INVX1 port map( A => n184, Y => n110);
   U654 : MUX2X1 port map( B => n74, A => n484, S => n485, Y => n1053);
   U655 : MUX2X1 port map( B => n76, A => n486, S => n485, Y => n1052);
   U656 : AOI21X1 port map( A => n105, B => n126, C => n58, Y => n485);
   U657 : INVX1 port map( A => n175, Y => n105);
   U658 : MUX2X1 port map( B => n74, A => n487, S => n488, Y => n1051);
   U659 : MUX2X1 port map( B => n76, A => n489, S => n488, Y => n1050);
   U660 : AOI21X1 port map( A => n100, B => n126, C => n59, Y => n488);
   U661 : NAND3X1 port map( A => n358, B => n64, C => n67, Y => n184);
   U662 : INVX1 port map( A => n235, Y => n100);
   U663 : MUX2X1 port map( B => n74, A => n490, S => n491, Y => n1049);
   U664 : MUX2X1 port map( B => n76, A => n492, S => n491, Y => n1048);
   U665 : AOI21X1 port map( A => n95, B => n126, C => n60, Y => n491);
   U666 : NAND3X1 port map( A => n69, B => n64, C => n67, Y => n175);
   U667 : NAND3X1 port map( A => n493, B => n70, C => n356, Y => n135);
   U668 : INVX1 port map( A => n226, Y => n95);
   U669 : MUX2X1 port map( B => n74, A => n494, S => n495, Y => n1047);
   U670 : INVX1 port map( A => opcode_28_1_port, Y => n494);
   U671 : MUX2X1 port map( B => n76, A => n496, S => n495, Y => n1046);
   U672 : AOI21X1 port map( A => n96, B => n130, C => n432, Y => n495);
   U673 : NAND3X1 port map( A => n358, B => n360, C => n65, Y => n235);
   U674 : INVX1 port map( A => n151, Y => n130);
   U675 : INVX1 port map( A => opcode_28_0_port, Y => n496);
   U676 : MUX2X1 port map( B => n74, A => n497, S => n498, Y => n1045);
   U677 : INVX1 port map( A => opcode_29_1_port, Y => n497);
   U678 : MUX2X1 port map( B => n76, A => n499, S => n498, Y => n1044);
   U679 : AOI21X1 port map( A => n96, B => n125, C => n61, Y => n498);
   U680 : NAND3X1 port map( A => n69, B => n360, C => n65, Y => n226);
   U681 : INVX1 port map( A => n145, Y => n125);
   U682 : NAND3X1 port map( A => n356, B => n493, C => n71, Y => n500);
   U683 : INVX1 port map( A => opcode_29_0_port, Y => n499);
   U684 : MUX2X1 port map( B => n74, A => n501, S => n502, Y => n1043);
   U685 : INVX1 port map( A => opcode_30_1_port, Y => n501);
   U686 : MUX2X1 port map( B => n76, A => n503, S => n502, Y => n1042);
   U687 : AOI21X1 port map( A => n120, B => n156, C => n62, Y => n502);
   U688 : NOR2X1 port map( A => n151, B => n174, Y => n449);
   U689 : NAND3X1 port map( A => n65, B => n358, C => n67, Y => n151);
   U690 : INVX1 port map( A => n140, Y => n120);
   U691 : NAND3X1 port map( A => n360, B => n64, C => n358, Y => n140);
   U692 : INVX1 port map( A => n69, Y => n358);
   U693 : INVX1 port map( A => opcode_30_0_port, Y => n503);
   U694 : MUX2X1 port map( B => n75, A => n504, S => n505, Y => n1041);
   U695 : INVX1 port map( A => opcode_31_1_port, Y => n504);
   U696 : MUX2X1 port map( B => n93, A => n506, S => n505, Y => n1040);
   U697 : AOI21X1 port map( A => n115, B => n156, C => n458, Y => n505);
   U698 : NOR2X1 port map( A => n507, B => n480, Y => n351);
   U699 : NOR2X1 port map( A => n354, B => RST, Y => n493);
   U700 : INVX1 port map( A => writeptr_4_port, Y => n354);
   U701 : NAND3X1 port map( A => n65, B => n69, C => n67, Y => n145);
   U702 : NAND3X1 port map( A => n356, B => n70, C => n352, Y => n508);
   U703 : NOR2X1 port map( A => writeptr_4_port, B => RST, Y => n352);
   U704 : NAND2X1 port map( A => W_ENABLE, B => n302, Y => n507);
   U705 : NAND3X1 port map( A => n509, B => n510, C => n511, Y => n302);
   U706 : NOR2X1 port map( A => n512, B => n513, Y => n511);
   U707 : XOR2X1 port map( A => readptr_3_port, B => N34, Y => n512);
   U708 : XOR2X1 port map( A => n514, B => N32, Y => n510);
   U709 : NOR2X1 port map( A => n515, B => n516, Y => n509);
   U710 : XOR2X1 port map( A => readptr_2_port, B => N33, Y => n515);
   U711 : INVX1 port map( A => n134, Y => n115);
   U712 : NAND3X1 port map( A => n360, B => n64, C => n69, Y => n134);
   U713 : INVX1 port map( A => n67, Y => n360);
   U714 : INVX1 port map( A => opcode_31_0_port, Y => n506);
   U715 : INVX1 port map( A => n517, Y => n1039);
   U716 : MUX2X1 port map( B => n518, A => DATA_7_port, S => n519, Y => n517);
   U717 : NAND2X1 port map( A => n520, B => n521, Y => n518);
   U718 : NOR2X1 port map( A => n522, B => n523, Y => n521);
   U719 : NAND3X1 port map( A => n524, B => n525, C => n526, Y => n523);
   U720 : NOR2X1 port map( A => n527, B => n528, Y => n526);
   U721 : OAI22X1 port map( A => n399, B => n529, C => n407, D => n530, Y => 
                           n528);
   U722 : INVX1 port map( A => memory_17_7_port, Y => n407);
   U723 : INVX1 port map( A => memory_16_7_port, Y => n399);
   U724 : OAI22X1 port map( A => n415, B => n531, C => n423, D => n532, Y => 
                           n527);
   U725 : INVX1 port map( A => memory_19_7_port, Y => n423);
   U726 : INVX1 port map( A => memory_18_7_port, Y => n415);
   U727 : AOI22X1 port map( A => n533, B => memory_23_7_port, C => n534, D => 
                           memory_22_7_port, Y => n525);
   U728 : AOI22X1 port map( A => n535, B => memory_21_7_port, C => n536, D => 
                           memory_20_7_port, Y => n524);
   U729 : NAND3X1 port map( A => n537, B => n538, C => n539, Y => n522);
   U730 : NOR2X1 port map( A => n540, B => n541, Y => n539);
   U731 : OAI22X1 port map( A => n193_port, B => n542, C => n185, D => n543, Y 
                           => n541);
   U732 : INVX1 port map( A => memory_25_7_port, Y => n185);
   U733 : INVX1 port map( A => memory_24_7_port, Y => n193_port);
   U734 : OAI22X1 port map( A => n176, B => n544, C => n166, D => n545, Y => 
                           n540);
   U735 : INVX1 port map( A => memory_27_7_port, Y => n166);
   U736 : INVX1 port map( A => memory_26_7_port, Y => n176);
   U737 : AOI22X1 port map( A => n546, B => memory_31_7_port, C => n547, D => 
                           memory_30_7_port, Y => n538);
   U738 : AOI22X1 port map( A => n548, B => memory_29_7_port, C => n549, D => 
                           memory_28_7_port, Y => n537);
   U739 : NOR2X1 port map( A => n550, B => n551, Y => n520);
   U740 : NAND3X1 port map( A => n552, B => n553, C => n554, Y => n551);
   U741 : NOR2X1 port map( A => n555, B => n556, Y => n554);
   U742 : OAI22X1 port map( A => n301, B => n557, C => n293, D => n558, Y => 
                           n556);
   U743 : INVX1 port map( A => memory_2_7_port, Y => n293);
   U744 : INVX1 port map( A => memory_3_7_port, Y => n301);
   U745 : OAI22X1 port map( A => n285, B => n559, C => n276, D => n560, Y => 
                           n555);
   U746 : INVX1 port map( A => memory_0_7_port, Y => n276);
   U747 : INVX1 port map( A => memory_1_7_port, Y => n285);
   U748 : AOI22X1 port map( A => n561, B => memory_4_7_port, C => n562, D => 
                           memory_5_7_port, Y => n553);
   U749 : AOI22X1 port map( A => n563, B => memory_6_7_port, C => n564, D => 
                           memory_7_7_port, Y => n552);
   U750 : NAND3X1 port map( A => n565, B => n566, C => n567, Y => n550);
   U751 : NOR2X1 port map( A => n568, B => n569, Y => n567);
   U752 : OAI22X1 port map( A => n363, B => n570, C => n372, D => n571, Y => 
                           n569);
   U753 : INVX1 port map( A => memory_9_7_port, Y => n372);
   U754 : INVX1 port map( A => memory_8_7_port, Y => n363);
   U755 : OAI22X1 port map( A => n381, B => n572, C => n390, D => n573, Y => 
                           n568);
   U756 : INVX1 port map( A => memory_11_7_port, Y => n390);
   U757 : INVX1 port map( A => memory_10_7_port, Y => n381);
   U758 : AOI22X1 port map( A => n574, B => memory_15_7_port, C => n575, D => 
                           memory_14_7_port, Y => n566);
   U759 : AOI22X1 port map( A => n576, B => memory_13_7_port, C => n577, D => 
                           memory_12_7_port, Y => n565);
   U760 : INVX1 port map( A => n578, Y => n1038);
   U761 : MUX2X1 port map( B => n579, A => DATA_6_port, S => n519, Y => n578);
   U762 : NAND2X1 port map( A => n580, B => n581, Y => n579);
   U763 : NOR2X1 port map( A => n582, B => n583, Y => n581);
   U764 : NAND3X1 port map( A => n584, B => n585, C => n586, Y => n583);
   U765 : NOR2X1 port map( A => n587, B => n588, Y => n586);
   U766 : OAI22X1 port map( A => n400, B => n529, C => n408, D => n530, Y => 
                           n588);
   U767 : INVX1 port map( A => memory_17_6_port, Y => n408);
   U768 : INVX1 port map( A => memory_16_6_port, Y => n400);
   U769 : OAI22X1 port map( A => n416, B => n531, C => n424, D => n532, Y => 
                           n587);
   U770 : INVX1 port map( A => memory_19_6_port, Y => n424);
   U771 : INVX1 port map( A => memory_18_6_port, Y => n416);
   U772 : AOI22X1 port map( A => n533, B => memory_23_6_port, C => n534, D => 
                           memory_22_6_port, Y => n585);
   U773 : AOI22X1 port map( A => n535, B => memory_21_6_port, C => n536, D => 
                           memory_20_6_port, Y => n584);
   U774 : NAND3X1 port map( A => n589, B => n590, C => n591, Y => n582);
   U775 : NOR2X1 port map( A => n592, B => n593, Y => n591);
   U776 : OAI22X1 port map( A => n194, B => n542, C => n186, D => n543, Y => 
                           n593);
   U777 : INVX1 port map( A => memory_25_6_port, Y => n186);
   U778 : INVX1 port map( A => memory_24_6_port, Y => n194);
   U779 : OAI22X1 port map( A => n177, B => n544, C => n167, D => n545, Y => 
                           n592);
   U780 : INVX1 port map( A => memory_27_6_port, Y => n167);
   U781 : INVX1 port map( A => memory_26_6_port, Y => n177);
   U782 : AOI22X1 port map( A => n546, B => memory_31_6_port, C => n547, D => 
                           memory_30_6_port, Y => n590);
   U783 : AOI22X1 port map( A => n548, B => memory_29_6_port, C => n549, D => 
                           memory_28_6_port, Y => n589);
   U784 : NOR2X1 port map( A => n594, B => n595, Y => n580);
   U785 : NAND3X1 port map( A => n596, B => n597, C => n598, Y => n595);
   U786 : NOR2X1 port map( A => n599, B => n600, Y => n598);
   U787 : OAI22X1 port map( A => n300, B => n557, C => n292, D => n558, Y => 
                           n600);
   U788 : INVX1 port map( A => memory_2_6_port, Y => n292);
   U789 : INVX1 port map( A => memory_3_6_port, Y => n300);
   U790 : OAI22X1 port map( A => n284, B => n559, C => n275, D => n560, Y => 
                           n599);
   U791 : INVX1 port map( A => memory_0_6_port, Y => n275);
   U792 : INVX1 port map( A => memory_1_6_port, Y => n284);
   U793 : AOI22X1 port map( A => n561, B => memory_4_6_port, C => n562, D => 
                           memory_5_6_port, Y => n597);
   U794 : AOI22X1 port map( A => n563, B => memory_6_6_port, C => n564, D => 
                           memory_7_6_port, Y => n596);
   U795 : NAND3X1 port map( A => n601, B => n602, C => n603, Y => n594);
   U796 : NOR2X1 port map( A => n604, B => n605, Y => n603);
   U797 : OAI22X1 port map( A => n365, B => n570, C => n374, D => n571, Y => 
                           n605);
   U798 : INVX1 port map( A => memory_9_6_port, Y => n374);
   U799 : INVX1 port map( A => memory_8_6_port, Y => n365);
   U800 : OAI22X1 port map( A => n383, B => n572, C => n392, D => n573, Y => 
                           n604);
   U801 : INVX1 port map( A => memory_11_6_port, Y => n392);
   U802 : INVX1 port map( A => memory_10_6_port, Y => n383);
   U803 : AOI22X1 port map( A => n574, B => memory_15_6_port, C => n575, D => 
                           memory_14_6_port, Y => n602);
   U804 : AOI22X1 port map( A => n576, B => memory_13_6_port, C => n577, D => 
                           memory_12_6_port, Y => n601);
   U805 : INVX1 port map( A => n606, Y => n1037);
   U806 : MUX2X1 port map( B => n607, A => DATA_5_port, S => n519, Y => n606);
   U807 : NAND2X1 port map( A => n608, B => n609, Y => n607);
   U808 : NOR2X1 port map( A => n610, B => n611, Y => n609);
   U809 : NAND3X1 port map( A => n612, B => n613, C => n614, Y => n611);
   U810 : NOR2X1 port map( A => n615, B => n616, Y => n614);
   U811 : OAI22X1 port map( A => n401, B => n529, C => n409, D => n530, Y => 
                           n616);
   U812 : INVX1 port map( A => memory_17_5_port, Y => n409);
   U813 : INVX1 port map( A => memory_16_5_port, Y => n401);
   U814 : OAI22X1 port map( A => n417, B => n531, C => n425, D => n532, Y => 
                           n615);
   U815 : INVX1 port map( A => memory_19_5_port, Y => n425);
   U816 : INVX1 port map( A => memory_18_5_port, Y => n417);
   U817 : AOI22X1 port map( A => n533, B => memory_23_5_port, C => n534, D => 
                           memory_22_5_port, Y => n613);
   U818 : AOI22X1 port map( A => n535, B => memory_21_5_port, C => n536, D => 
                           memory_20_5_port, Y => n612);
   U819 : NAND3X1 port map( A => n617, B => n618, C => n619, Y => n610);
   U820 : NOR2X1 port map( A => n620, B => n621, Y => n619);
   U821 : OAI22X1 port map( A => n195_port, B => n542, C => n187, D => n543, Y 
                           => n621);
   U822 : INVX1 port map( A => memory_25_5_port, Y => n187);
   U823 : INVX1 port map( A => memory_24_5_port, Y => n195_port);
   U824 : OAI22X1 port map( A => n178, B => n544, C => n168, D => n545, Y => 
                           n620);
   U825 : INVX1 port map( A => memory_27_5_port, Y => n168);
   U826 : INVX1 port map( A => memory_26_5_port, Y => n178);
   U827 : AOI22X1 port map( A => n546, B => memory_31_5_port, C => n547, D => 
                           memory_30_5_port, Y => n618);
   U828 : AOI22X1 port map( A => n548, B => memory_29_5_port, C => n549, D => 
                           memory_28_5_port, Y => n617);
   U829 : NOR2X1 port map( A => n622, B => n623, Y => n608);
   U830 : NAND3X1 port map( A => n624, B => n625, C => n626, Y => n623);
   U831 : NOR2X1 port map( A => n627, B => n628, Y => n626);
   U832 : OAI22X1 port map( A => n299, B => n557, C => n291, D => n558, Y => 
                           n628);
   U833 : INVX1 port map( A => memory_2_5_port, Y => n291);
   U834 : INVX1 port map( A => memory_3_5_port, Y => n299);
   U835 : OAI22X1 port map( A => n283, B => n559, C => n274, D => n560, Y => 
                           n627);
   U836 : INVX1 port map( A => memory_0_5_port, Y => n274);
   U837 : INVX1 port map( A => memory_1_5_port, Y => n283);
   U838 : AOI22X1 port map( A => n561, B => memory_4_5_port, C => n562, D => 
                           memory_5_5_port, Y => n625);
   U839 : AOI22X1 port map( A => n563, B => memory_6_5_port, C => n564, D => 
                           memory_7_5_port, Y => n624);
   U840 : NAND3X1 port map( A => n629, B => n630, C => n631, Y => n622);
   U841 : NOR2X1 port map( A => n632, B => n633, Y => n631);
   U842 : OAI22X1 port map( A => n366, B => n570, C => n375, D => n571, Y => 
                           n633);
   U843 : INVX1 port map( A => memory_9_5_port, Y => n375);
   U844 : INVX1 port map( A => memory_8_5_port, Y => n366);
   U845 : OAI22X1 port map( A => n384, B => n572, C => n393, D => n573, Y => 
                           n632);
   U846 : INVX1 port map( A => memory_11_5_port, Y => n393);
   U847 : INVX1 port map( A => memory_10_5_port, Y => n384);
   U848 : AOI22X1 port map( A => n574, B => memory_15_5_port, C => n575, D => 
                           memory_14_5_port, Y => n630);
   U849 : AOI22X1 port map( A => n576, B => memory_13_5_port, C => n577, D => 
                           memory_12_5_port, Y => n629);
   U850 : INVX1 port map( A => n634, Y => n1036);
   U851 : MUX2X1 port map( B => n635, A => DATA_4_port, S => n519, Y => n634);
   U852 : NAND2X1 port map( A => n636, B => n637, Y => n635);
   U853 : NOR2X1 port map( A => n638, B => n639, Y => n637);
   U854 : NAND3X1 port map( A => n640, B => n641, C => n642, Y => n639);
   U855 : NOR2X1 port map( A => n643, B => n644, Y => n642);
   U856 : OAI22X1 port map( A => n402, B => n529, C => n410, D => n530, Y => 
                           n644);
   U857 : INVX1 port map( A => memory_17_4_port, Y => n410);
   U858 : INVX1 port map( A => memory_16_4_port, Y => n402);
   U859 : OAI22X1 port map( A => n418, B => n531, C => n426, D => n532, Y => 
                           n643);
   U860 : INVX1 port map( A => memory_19_4_port, Y => n426);
   U861 : INVX1 port map( A => memory_18_4_port, Y => n418);
   U862 : AOI22X1 port map( A => n533, B => memory_23_4_port, C => n534, D => 
                           memory_22_4_port, Y => n641);
   U863 : AOI22X1 port map( A => n535, B => memory_21_4_port, C => n536, D => 
                           memory_20_4_port, Y => n640);
   U864 : NAND3X1 port map( A => n645, B => n646, C => n647, Y => n638);
   U865 : NOR2X1 port map( A => n648, B => n649, Y => n647);
   U866 : OAI22X1 port map( A => n196, B => n542, C => n188, D => n543, Y => 
                           n649);
   U867 : INVX1 port map( A => memory_25_4_port, Y => n188);
   U868 : INVX1 port map( A => memory_24_4_port, Y => n196);
   U869 : OAI22X1 port map( A => n179, B => n544, C => n169, D => n545, Y => 
                           n648);
   U870 : INVX1 port map( A => memory_27_4_port, Y => n169);
   U871 : INVX1 port map( A => memory_26_4_port, Y => n179);
   U872 : AOI22X1 port map( A => n546, B => memory_31_4_port, C => n547, D => 
                           memory_30_4_port, Y => n646);
   U873 : AOI22X1 port map( A => n548, B => memory_29_4_port, C => n549, D => 
                           memory_28_4_port, Y => n645);
   U874 : NOR2X1 port map( A => n650, B => n651, Y => n636);
   U875 : NAND3X1 port map( A => n652, B => n653, C => n654, Y => n651);
   U876 : NOR2X1 port map( A => n655, B => n656, Y => n654);
   U877 : OAI22X1 port map( A => n298, B => n557, C => n290, D => n558, Y => 
                           n656);
   U878 : INVX1 port map( A => memory_2_4_port, Y => n290);
   U879 : INVX1 port map( A => memory_3_4_port, Y => n298);
   U880 : OAI22X1 port map( A => n282, B => n559, C => n273, D => n560, Y => 
                           n655);
   U881 : INVX1 port map( A => memory_0_4_port, Y => n273);
   U882 : INVX1 port map( A => memory_1_4_port, Y => n282);
   U883 : AOI22X1 port map( A => n561, B => memory_4_4_port, C => n562, D => 
                           memory_5_4_port, Y => n653);
   U884 : AOI22X1 port map( A => n563, B => memory_6_4_port, C => n564, D => 
                           memory_7_4_port, Y => n652);
   U885 : NAND3X1 port map( A => n657, B => n658, C => n659, Y => n650);
   U886 : NOR2X1 port map( A => n660, B => n661, Y => n659);
   U887 : OAI22X1 port map( A => n367, B => n570, C => n376, D => n571, Y => 
                           n661);
   U888 : INVX1 port map( A => memory_9_4_port, Y => n376);
   U889 : INVX1 port map( A => memory_8_4_port, Y => n367);
   U890 : OAI22X1 port map( A => n385, B => n572, C => n394, D => n573, Y => 
                           n660);
   U891 : INVX1 port map( A => memory_11_4_port, Y => n394);
   U892 : INVX1 port map( A => memory_10_4_port, Y => n385);
   U893 : AOI22X1 port map( A => n574, B => memory_15_4_port, C => n575, D => 
                           memory_14_4_port, Y => n658);
   U894 : AOI22X1 port map( A => n576, B => memory_13_4_port, C => n577, D => 
                           memory_12_4_port, Y => n657);
   U895 : INVX1 port map( A => n662, Y => n1035);
   U896 : MUX2X1 port map( B => n663, A => DATA_3_port, S => n519, Y => n662);
   U897 : NAND2X1 port map( A => n664, B => n665, Y => n663);
   U898 : NOR2X1 port map( A => n666, B => n667, Y => n665);
   U899 : NAND3X1 port map( A => n668, B => n669, C => n670, Y => n667);
   U900 : NOR2X1 port map( A => n671, B => n672, Y => n670);
   U901 : OAI22X1 port map( A => n403, B => n529, C => n411, D => n530, Y => 
                           n672);
   U902 : INVX1 port map( A => memory_17_3_port, Y => n411);
   U903 : INVX1 port map( A => memory_16_3_port, Y => n403);
   U904 : OAI22X1 port map( A => n419, B => n531, C => n427, D => n532, Y => 
                           n671);
   U905 : INVX1 port map( A => memory_19_3_port, Y => n427);
   U906 : INVX1 port map( A => memory_18_3_port, Y => n419);
   U907 : AOI22X1 port map( A => n533, B => memory_23_3_port, C => n534, D => 
                           memory_22_3_port, Y => n669);
   U908 : AOI22X1 port map( A => n535, B => memory_21_3_port, C => n536, D => 
                           memory_20_3_port, Y => n668);
   U909 : NAND3X1 port map( A => n673, B => n674, C => n675, Y => n666);
   U910 : NOR2X1 port map( A => n676, B => n677, Y => n675);
   U911 : OAI22X1 port map( A => n197, B => n542, C => n189_port, D => n543, Y 
                           => n677);
   U912 : INVX1 port map( A => memory_25_3_port, Y => n189_port);
   U913 : INVX1 port map( A => memory_24_3_port, Y => n197);
   U914 : OAI22X1 port map( A => n180, B => n544, C => n170, D => n545, Y => 
                           n676);
   U915 : INVX1 port map( A => memory_27_3_port, Y => n170);
   U916 : INVX1 port map( A => memory_26_3_port, Y => n180);
   U917 : AOI22X1 port map( A => n546, B => memory_31_3_port, C => n547, D => 
                           memory_30_3_port, Y => n674);
   U918 : AOI22X1 port map( A => n548, B => memory_29_3_port, C => n549, D => 
                           memory_28_3_port, Y => n673);
   U919 : NOR2X1 port map( A => n678, B => n679, Y => n664);
   U920 : NAND3X1 port map( A => n680, B => n681, C => n682, Y => n679);
   U921 : NOR2X1 port map( A => n683, B => n684, Y => n682);
   U922 : OAI22X1 port map( A => n297, B => n557, C => n289, D => n558, Y => 
                           n684);
   U923 : INVX1 port map( A => memory_2_3_port, Y => n289);
   U924 : INVX1 port map( A => memory_3_3_port, Y => n297);
   U925 : OAI22X1 port map( A => n281, B => n559, C => n272, D => n560, Y => 
                           n683);
   U926 : INVX1 port map( A => memory_0_3_port, Y => n272);
   U927 : INVX1 port map( A => memory_1_3_port, Y => n281);
   U928 : AOI22X1 port map( A => n561, B => memory_4_3_port, C => n562, D => 
                           memory_5_3_port, Y => n681);
   U929 : AOI22X1 port map( A => n563, B => memory_6_3_port, C => n564, D => 
                           memory_7_3_port, Y => n680);
   U930 : NAND3X1 port map( A => n685, B => n686, C => n687, Y => n678);
   U931 : NOR2X1 port map( A => n688, B => n689, Y => n687);
   U932 : OAI22X1 port map( A => n368, B => n570, C => n377, D => n571, Y => 
                           n689);
   U933 : INVX1 port map( A => memory_9_3_port, Y => n377);
   U934 : INVX1 port map( A => memory_8_3_port, Y => n368);
   U935 : OAI22X1 port map( A => n386, B => n572, C => n395, D => n573, Y => 
                           n688);
   U936 : INVX1 port map( A => memory_11_3_port, Y => n395);
   U937 : INVX1 port map( A => memory_10_3_port, Y => n386);
   U938 : AOI22X1 port map( A => n574, B => memory_15_3_port, C => n575, D => 
                           memory_14_3_port, Y => n686);
   U939 : AOI22X1 port map( A => n576, B => memory_13_3_port, C => n577, D => 
                           memory_12_3_port, Y => n685);
   U940 : INVX1 port map( A => n690, Y => n1034);
   U941 : MUX2X1 port map( B => n691, A => DATA_2_port, S => n519, Y => n690);
   U942 : NAND2X1 port map( A => n692, B => n693, Y => n691);
   U943 : NOR2X1 port map( A => n694, B => n695, Y => n693);
   U944 : NAND3X1 port map( A => n696, B => n697, C => n698, Y => n695);
   U945 : NOR2X1 port map( A => n699, B => n700, Y => n698);
   U946 : OAI22X1 port map( A => n404, B => n529, C => n412, D => n530, Y => 
                           n700);
   U947 : INVX1 port map( A => memory_17_2_port, Y => n412);
   U948 : INVX1 port map( A => memory_16_2_port, Y => n404);
   U949 : OAI22X1 port map( A => n420, B => n531, C => n428, D => n532, Y => 
                           n699);
   U950 : INVX1 port map( A => memory_19_2_port, Y => n428);
   U951 : INVX1 port map( A => memory_18_2_port, Y => n420);
   U952 : AOI22X1 port map( A => n533, B => memory_23_2_port, C => n534, D => 
                           memory_22_2_port, Y => n697);
   U953 : AOI22X1 port map( A => n535, B => memory_21_2_port, C => n536, D => 
                           memory_20_2_port, Y => n696);
   U954 : NAND3X1 port map( A => n701, B => n702, C => n703, Y => n694);
   U955 : NOR2X1 port map( A => n704, B => n705, Y => n703);
   U956 : OAI22X1 port map( A => n198, B => n542, C => n190_port, D => n543, Y 
                           => n705);
   U957 : INVX1 port map( A => memory_25_2_port, Y => n190_port);
   U958 : INVX1 port map( A => memory_24_2_port, Y => n198);
   U959 : OAI22X1 port map( A => n181, B => n544, C => n171, D => n545, Y => 
                           n704);
   U960 : INVX1 port map( A => memory_27_2_port, Y => n171);
   U961 : INVX1 port map( A => memory_26_2_port, Y => n181);
   U962 : AOI22X1 port map( A => n546, B => memory_31_2_port, C => n547, D => 
                           memory_30_2_port, Y => n702);
   U963 : AOI22X1 port map( A => n548, B => memory_29_2_port, C => n549, D => 
                           memory_28_2_port, Y => n701);
   U964 : NOR2X1 port map( A => n706, B => n707, Y => n692);
   U965 : NAND3X1 port map( A => n708, B => n709, C => n710, Y => n707);
   U966 : NOR2X1 port map( A => n711, B => n712, Y => n710);
   U967 : OAI22X1 port map( A => n296, B => n557, C => n288, D => n558, Y => 
                           n712);
   U968 : INVX1 port map( A => memory_2_2_port, Y => n288);
   U969 : INVX1 port map( A => memory_3_2_port, Y => n296);
   U970 : OAI22X1 port map( A => n280, B => n559, C => n271, D => n560, Y => 
                           n711);
   U971 : INVX1 port map( A => memory_0_2_port, Y => n271);
   U972 : INVX1 port map( A => memory_1_2_port, Y => n280);
   U973 : AOI22X1 port map( A => n561, B => memory_4_2_port, C => n562, D => 
                           memory_5_2_port, Y => n709);
   U974 : AOI22X1 port map( A => n563, B => memory_6_2_port, C => n564, D => 
                           memory_7_2_port, Y => n708);
   U975 : NAND3X1 port map( A => n713, B => n714, C => n715, Y => n706);
   U976 : NOR2X1 port map( A => n716, B => n717, Y => n715);
   U977 : OAI22X1 port map( A => n369, B => n570, C => n378, D => n571, Y => 
                           n717);
   U978 : INVX1 port map( A => memory_9_2_port, Y => n378);
   U979 : INVX1 port map( A => memory_8_2_port, Y => n369);
   U980 : OAI22X1 port map( A => n387, B => n572, C => n396, D => n573, Y => 
                           n716);
   U981 : INVX1 port map( A => memory_11_2_port, Y => n396);
   U982 : INVX1 port map( A => memory_10_2_port, Y => n387);
   U983 : AOI22X1 port map( A => n574, B => memory_15_2_port, C => n575, D => 
                           memory_14_2_port, Y => n714);
   U984 : AOI22X1 port map( A => n576, B => memory_13_2_port, C => n577, D => 
                           memory_12_2_port, Y => n713);
   U985 : INVX1 port map( A => n718, Y => n1033);
   U986 : MUX2X1 port map( B => n719, A => DATA_1_port, S => n519, Y => n718);
   U987 : NAND2X1 port map( A => n720, B => n721, Y => n719);
   U988 : NOR2X1 port map( A => n722, B => n723, Y => n721);
   U989 : NAND3X1 port map( A => n724, B => n725, C => n726, Y => n723);
   U990 : NOR2X1 port map( A => n727, B => n728, Y => n726);
   U991 : OAI22X1 port map( A => n405, B => n529, C => n413, D => n530, Y => 
                           n728);
   U992 : INVX1 port map( A => memory_17_1_port, Y => n413);
   U993 : INVX1 port map( A => memory_16_1_port, Y => n405);
   U994 : OAI22X1 port map( A => n421, B => n531, C => n429, D => n532, Y => 
                           n727);
   U995 : INVX1 port map( A => memory_19_1_port, Y => n429);
   U996 : INVX1 port map( A => memory_18_1_port, Y => n421);
   U997 : AOI22X1 port map( A => n533, B => memory_23_1_port, C => n534, D => 
                           memory_22_1_port, Y => n725);
   U998 : AOI22X1 port map( A => n535, B => memory_21_1_port, C => n536, D => 
                           memory_20_1_port, Y => n724);
   U999 : NAND3X1 port map( A => n729, B => n730, C => n731, Y => n722);
   U1000 : NOR2X1 port map( A => n732, B => n733, Y => n731);
   U1001 : OAI22X1 port map( A => n199, B => n542, C => n191_port, D => n543, Y
                           => n733);
   U1002 : INVX1 port map( A => memory_25_1_port, Y => n191_port);
   U1003 : INVX1 port map( A => memory_24_1_port, Y => n199);
   U1004 : OAI22X1 port map( A => n182, B => n544, C => n172, D => n545, Y => 
                           n732);
   U1005 : INVX1 port map( A => memory_27_1_port, Y => n172);
   U1006 : INVX1 port map( A => memory_26_1_port, Y => n182);
   U1007 : AOI22X1 port map( A => n546, B => memory_31_1_port, C => n547, D => 
                           memory_30_1_port, Y => n730);
   U1008 : AOI22X1 port map( A => n548, B => memory_29_1_port, C => n549, D => 
                           memory_28_1_port, Y => n729);
   U1009 : NOR2X1 port map( A => n734, B => n735, Y => n720);
   U1010 : NAND3X1 port map( A => n736, B => n737, C => n738, Y => n735);
   U1011 : NOR2X1 port map( A => n739, B => n740, Y => n738);
   U1012 : OAI22X1 port map( A => n295, B => n557, C => n287, D => n558, Y => 
                           n740);
   U1013 : INVX1 port map( A => memory_2_1_port, Y => n287);
   U1014 : INVX1 port map( A => memory_3_1_port, Y => n295);
   U1015 : OAI22X1 port map( A => n279, B => n559, C => n270, D => n560, Y => 
                           n739);
   U1016 : INVX1 port map( A => memory_0_1_port, Y => n270);
   U1017 : INVX1 port map( A => memory_1_1_port, Y => n279);
   U1018 : AOI22X1 port map( A => n561, B => memory_4_1_port, C => n562, D => 
                           memory_5_1_port, Y => n737);
   U1019 : AOI22X1 port map( A => n563, B => memory_6_1_port, C => n564, D => 
                           memory_7_1_port, Y => n736);
   U1020 : NAND3X1 port map( A => n741, B => n742, C => n743, Y => n734);
   U1021 : NOR2X1 port map( A => n744, B => n745, Y => n743);
   U1022 : OAI22X1 port map( A => n370, B => n570, C => n379, D => n571, Y => 
                           n745);
   U1023 : INVX1 port map( A => memory_9_1_port, Y => n379);
   U1024 : INVX1 port map( A => memory_8_1_port, Y => n370);
   U1025 : OAI22X1 port map( A => n388, B => n572, C => n397, D => n573, Y => 
                           n744);
   U1026 : INVX1 port map( A => memory_11_1_port, Y => n397);
   U1027 : INVX1 port map( A => memory_10_1_port, Y => n388);
   U1028 : AOI22X1 port map( A => n574, B => memory_15_1_port, C => n575, D => 
                           memory_14_1_port, Y => n742);
   U1029 : AOI22X1 port map( A => n576, B => memory_13_1_port, C => n577, D => 
                           memory_12_1_port, Y => n741);
   U1030 : INVX1 port map( A => n746, Y => n1032);
   U1031 : MUX2X1 port map( B => n747, A => DATA_0_port, S => n519, Y => n746);
   U1032 : NAND2X1 port map( A => n748, B => n749, Y => n747);
   U1033 : NOR2X1 port map( A => n750, B => n751, Y => n749);
   U1034 : NAND3X1 port map( A => n752, B => n753, C => n754, Y => n751);
   U1035 : NOR2X1 port map( A => n755, B => n756, Y => n754);
   U1036 : OAI22X1 port map( A => n406, B => n529, C => n414, D => n530, Y => 
                           n756);
   U1037 : INVX1 port map( A => memory_17_0_port, Y => n414);
   U1038 : INVX1 port map( A => memory_16_0_port, Y => n406);
   U1039 : OAI22X1 port map( A => n422, B => n531, C => n430, D => n532, Y => 
                           n755);
   U1040 : INVX1 port map( A => memory_19_0_port, Y => n430);
   U1041 : INVX1 port map( A => memory_18_0_port, Y => n422);
   U1042 : AOI22X1 port map( A => n533, B => memory_23_0_port, C => n534, D => 
                           memory_22_0_port, Y => n753);
   U1043 : AOI22X1 port map( A => n535, B => memory_21_0_port, C => n536, D => 
                           memory_20_0_port, Y => n752);
   U1044 : NAND3X1 port map( A => n757, B => n758, C => n759, Y => n750);
   U1045 : NOR2X1 port map( A => n760, B => n761, Y => n759);
   U1046 : OAI22X1 port map( A => n200, B => n542, C => n192_port, D => n543, Y
                           => n761);
   U1047 : INVX1 port map( A => memory_25_0_port, Y => n192_port);
   U1048 : INVX1 port map( A => memory_24_0_port, Y => n200);
   U1049 : OAI22X1 port map( A => n183, B => n544, C => n173, D => n545, Y => 
                           n760);
   U1050 : INVX1 port map( A => memory_27_0_port, Y => n173);
   U1051 : INVX1 port map( A => memory_26_0_port, Y => n183);
   U1052 : AOI22X1 port map( A => n546, B => memory_31_0_port, C => n547, D => 
                           memory_30_0_port, Y => n758);
   U1053 : AOI22X1 port map( A => n548, B => memory_29_0_port, C => n549, D => 
                           memory_28_0_port, Y => n757);
   U1054 : NOR2X1 port map( A => n762, B => n763, Y => n748);
   U1055 : NAND3X1 port map( A => n764, B => n765, C => n766, Y => n763);
   U1056 : NOR2X1 port map( A => n767, B => n768, Y => n766);
   U1057 : OAI22X1 port map( A => n294, B => n557, C => n286, D => n558, Y => 
                           n768);
   U1058 : INVX1 port map( A => memory_2_0_port, Y => n286);
   U1059 : INVX1 port map( A => memory_3_0_port, Y => n294);
   U1060 : OAI22X1 port map( A => n278, B => n559, C => n269, D => n560, Y => 
                           n767);
   U1061 : INVX1 port map( A => memory_0_0_port, Y => n269);
   U1062 : INVX1 port map( A => memory_1_0_port, Y => n278);
   U1063 : AOI22X1 port map( A => n561, B => memory_4_0_port, C => n562, D => 
                           memory_5_0_port, Y => n765);
   U1064 : AOI22X1 port map( A => n563, B => memory_6_0_port, C => n564, D => 
                           memory_7_0_port, Y => n764);
   U1065 : NAND3X1 port map( A => n769, B => n770, C => n771, Y => n762);
   U1066 : NOR2X1 port map( A => n772, B => n773, Y => n771);
   U1067 : OAI22X1 port map( A => n371, B => n570, C => n380, D => n571, Y => 
                           n773);
   U1068 : INVX1 port map( A => memory_9_0_port, Y => n380);
   U1069 : INVX1 port map( A => memory_8_0_port, Y => n371);
   U1070 : OAI22X1 port map( A => n389, B => n572, C => n398, D => n573, Y => 
                           n772);
   U1071 : INVX1 port map( A => memory_11_0_port, Y => n398);
   U1072 : INVX1 port map( A => memory_10_0_port, Y => n389);
   U1073 : AOI22X1 port map( A => n574, B => memory_15_0_port, C => n575, D => 
                           memory_14_0_port, Y => n770);
   U1074 : AOI22X1 port map( A => n576, B => memory_13_0_port, C => n577, D => 
                           memory_12_0_port, Y => n769);
   U1075 : INVX1 port map( A => n774, Y => n1031);
   U1076 : MUX2X1 port map( B => n775, A => OUT_OPCODE_1_port, S => n519, Y => 
                           n774);
   U1077 : NAND2X1 port map( A => n776, B => n777, Y => n775);
   U1078 : NOR2X1 port map( A => n778, B => n779, Y => n777);
   U1079 : NAND3X1 port map( A => n780, B => n781, C => n782, Y => n779);
   U1080 : NOR2X1 port map( A => n783, B => n784, Y => n782);
   U1081 : OAI22X1 port map( A => n481, B => n529, C => n484, D => n530, Y => 
                           n784);
   U1082 : INVX1 port map( A => opcode_17_1_port, Y => n484);
   U1083 : INVX1 port map( A => opcode_16_1_port, Y => n481);
   U1084 : OAI22X1 port map( A => n487, B => n531, C => n490, D => n532, Y => 
                           n783);
   U1085 : INVX1 port map( A => opcode_19_1_port, Y => n490);
   U1086 : INVX1 port map( A => opcode_18_1_port, Y => n487);
   U1087 : AOI22X1 port map( A => n533, B => opcode_23_1_port, C => n534, D => 
                           opcode_22_1_port, Y => n781);
   U1088 : AOI22X1 port map( A => n535, B => opcode_21_1_port, C => n536, D => 
                           opcode_20_1_port, Y => n780);
   U1089 : NAND3X1 port map( A => n785, B => n786, C => n787, Y => n778);
   U1090 : NOR2X1 port map( A => n788, B => n789, Y => n787);
   U1091 : OAI22X1 port map( A => n107, B => n542, C => n102, D => n543, Y => 
                           n789);
   U1092 : INVX1 port map( A => opcode_25_1_port, Y => n102);
   U1093 : INVX1 port map( A => opcode_24_1_port, Y => n107);
   U1094 : OAI22X1 port map( A => n97, B => n544, C => n91, D => n545, Y => 
                           n788);
   U1095 : INVX1 port map( A => opcode_27_1_port, Y => n91);
   U1096 : INVX1 port map( A => opcode_26_1_port, Y => n97);
   U1097 : AOI22X1 port map( A => n546, B => opcode_31_1_port, C => n547, D => 
                           opcode_30_1_port, Y => n786);
   U1098 : AOI22X1 port map( A => n548, B => opcode_29_1_port, C => n549, D => 
                           opcode_28_1_port, Y => n785);
   U1099 : NOR2X1 port map( A => n790, B => n791, Y => n776);
   U1100 : NAND3X1 port map( A => n792, B => n793, C => n794, Y => n791);
   U1101 : NOR2X1 port map( A => n795, B => n796, Y => n794);
   U1102 : OAI22X1 port map( A => n165, B => n557, C => n162, D => n558, Y => 
                           n796);
   U1103 : INVX1 port map( A => opcode_2_1_port, Y => n162);
   U1104 : INVX1 port map( A => opcode_3_1_port, Y => n165);
   U1105 : OAI22X1 port map( A => n159, B => n559, C => n155, D => n560, Y => 
                           n795);
   U1106 : INVX1 port map( A => opcode_0_1_port, Y => n155);
   U1107 : INVX1 port map( A => opcode_1_1_port, Y => n159);
   U1108 : AOI22X1 port map( A => n561, B => opcode_4_1_port, C => n562, D => 
                           opcode_5_1_port, Y => n793);
   U1109 : AOI22X1 port map( A => n563, B => opcode_6_1_port, C => n564, D => 
                           opcode_7_1_port, Y => n792);
   U1110 : NAND3X1 port map( A => n797, B => n798, C => n799, Y => n790);
   U1111 : NOR2X1 port map( A => n800, B => n801, Y => n799);
   U1112 : OAI22X1 port map( A => n466, B => n570, C => n469, D => n571, Y => 
                           n801);
   U1113 : INVX1 port map( A => opcode_9_1_port, Y => n469);
   U1114 : INVX1 port map( A => opcode_8_1_port, Y => n466);
   U1115 : OAI22X1 port map( A => n472, B => n572, C => n476, D => n573, Y => 
                           n800);
   U1116 : INVX1 port map( A => opcode_11_1_port, Y => n476);
   U1117 : INVX1 port map( A => opcode_10_1_port, Y => n472);
   U1118 : AOI22X1 port map( A => n574, B => opcode_15_1_port, C => n575, D => 
                           opcode_14_1_port, Y => n798);
   U1119 : AOI22X1 port map( A => n576, B => opcode_13_1_port, C => n577, D => 
                           opcode_12_1_port, Y => n797);
   U1120 : INVX1 port map( A => n802, Y => n1030);
   U1121 : MUX2X1 port map( B => n803, A => OUT_OPCODE_0_port, S => n519, Y => 
                           n802);
   U1122 : NAND3X1 port map( A => N195, B => n85, C => n72, Y => n519);
   U1123 : NAND2X1 port map( A => n804, B => n805, Y => n803);
   U1124 : NOR2X1 port map( A => n806, B => n807, Y => n805);
   U1125 : NAND3X1 port map( A => n808, B => n809, C => n810, Y => n807);
   U1126 : NOR2X1 port map( A => n811, B => n812, Y => n810);
   U1127 : OAI22X1 port map( A => n483, B => n529, C => n486, D => n530, Y => 
                           n812);
   U1128 : NAND2X1 port map( A => n813, B => n814, Y => n530);
   U1129 : INVX1 port map( A => opcode_17_0_port, Y => n486);
   U1130 : NAND2X1 port map( A => n815, B => n814, Y => n529);
   U1131 : INVX1 port map( A => opcode_16_0_port, Y => n483);
   U1132 : OAI22X1 port map( A => n489, B => n531, C => n492, D => n532, Y => 
                           n811);
   U1133 : NAND2X1 port map( A => n813, B => n816, Y => n532);
   U1134 : INVX1 port map( A => opcode_19_0_port, Y => n492);
   U1135 : NAND2X1 port map( A => n815, B => n816, Y => n531);
   U1136 : INVX1 port map( A => opcode_18_0_port, Y => n489);
   U1137 : AOI22X1 port map( A => n533, B => opcode_23_0_port, C => n534, D => 
                           opcode_22_0_port, Y => n809);
   U1138 : AOI22X1 port map( A => n535, B => opcode_21_0_port, C => n536, D => 
                           opcode_20_0_port, Y => n808);
   U1139 : INVX1 port map( A => n819, Y => n815);
   U1140 : NAND3X1 port map( A => n820, B => n821, C => readptr_4_port, Y => 
                           n819);
   U1141 : INVX1 port map( A => n822, Y => n813);
   U1142 : NAND3X1 port map( A => readptr_0_port, B => n821, C => 
                           readptr_4_port, Y => n822);
   U1143 : NAND3X1 port map( A => n823, B => n824, C => n825, Y => n806);
   U1144 : NOR2X1 port map( A => n826, B => n827, Y => n825);
   U1145 : OAI22X1 port map( A => n109, B => n542, C => n104, D => n543, Y => 
                           n827);
   U1146 : NAND2X1 port map( A => n814, B => n828, Y => n543);
   U1147 : INVX1 port map( A => opcode_25_0_port, Y => n104);
   U1148 : NAND2X1 port map( A => n814, B => n829, Y => n542);
   U1149 : INVX1 port map( A => opcode_24_0_port, Y => n109);
   U1150 : OAI22X1 port map( A => n99, B => n544, C => n94, D => n545, Y => 
                           n826);
   U1151 : NAND2X1 port map( A => n816, B => n828, Y => n545);
   U1152 : INVX1 port map( A => opcode_27_0_port, Y => n94);
   U1153 : NAND2X1 port map( A => n816, B => n829, Y => n544);
   U1154 : INVX1 port map( A => opcode_26_0_port, Y => n99);
   U1155 : AOI22X1 port map( A => n546, B => opcode_31_0_port, C => n547, D => 
                           opcode_30_0_port, Y => n824);
   U1156 : AOI22X1 port map( A => n548, B => opcode_29_0_port, C => n549, D => 
                           opcode_28_0_port, Y => n823);
   U1157 : INVX1 port map( A => n830, Y => n829);
   U1158 : NAND3X1 port map( A => readptr_3_port, B => n820, C => 
                           readptr_4_port, Y => n830);
   U1159 : INVX1 port map( A => n831, Y => n828);
   U1160 : NAND3X1 port map( A => readptr_3_port, B => readptr_0_port, C => 
                           readptr_4_port, Y => n831);
   U1161 : NOR2X1 port map( A => n832, B => n833, Y => n804);
   U1162 : NAND3X1 port map( A => n834, B => n835, C => n836, Y => n833);
   U1163 : NOR2X1 port map( A => n837, B => n838, Y => n836);
   U1164 : OAI22X1 port map( A => n163, B => n557, C => n160, D => n558, Y => 
                           n838);
   U1165 : NAND2X1 port map( A => n839, B => n816, Y => n558);
   U1166 : INVX1 port map( A => opcode_2_0_port, Y => n160);
   U1167 : NAND2X1 port map( A => n840, B => n816, Y => n557);
   U1168 : INVX1 port map( A => opcode_3_0_port, Y => n163);
   U1169 : OAI22X1 port map( A => n157, B => n559, C => n153, D => n560, Y => 
                           n837);
   U1170 : NAND2X1 port map( A => n839, B => n814, Y => n560);
   U1171 : INVX1 port map( A => opcode_0_0_port, Y => n153);
   U1172 : NAND2X1 port map( A => n840, B => n814, Y => n559);
   U1173 : INVX1 port map( A => opcode_1_0_port, Y => n157);
   U1174 : AOI22X1 port map( A => n561, B => opcode_4_0_port, C => n562, D => 
                           opcode_5_0_port, Y => n835);
   U1175 : AOI22X1 port map( A => n563, B => opcode_6_0_port, C => n564, D => 
                           opcode_7_0_port, Y => n834);
   U1176 : INVX1 port map( A => n841, Y => n840);
   U1177 : NAND3X1 port map( A => n821, B => n842, C => readptr_0_port, Y => 
                           n841);
   U1178 : INVX1 port map( A => n843, Y => n839);
   U1179 : NAND3X1 port map( A => n821, B => n842, C => n820, Y => n843);
   U1180 : INVX1 port map( A => readptr_3_port, Y => n821);
   U1181 : NAND3X1 port map( A => n844, B => n845, C => n846, Y => n832);
   U1182 : NOR2X1 port map( A => n847, B => n848, Y => n846);
   U1183 : OAI22X1 port map( A => n468, B => n570, C => n471, D => n571, Y => 
                           n848);
   U1184 : NAND2X1 port map( A => n849, B => n814, Y => n571);
   U1185 : INVX1 port map( A => opcode_9_0_port, Y => n471);
   U1186 : NAND2X1 port map( A => n850, B => n814, Y => n570);
   U1187 : NOR2X1 port map( A => readptr_1_port, B => readptr_2_port, Y => n814
                           );
   U1188 : INVX1 port map( A => opcode_8_0_port, Y => n468);
   U1189 : OAI22X1 port map( A => n474, B => n572, C => n478, D => n573, Y => 
                           n847);
   U1190 : NAND2X1 port map( A => n849, B => n816, Y => n573);
   U1191 : INVX1 port map( A => opcode_11_0_port, Y => n478);
   U1192 : NAND2X1 port map( A => n850, B => n816, Y => n572);
   U1193 : NOR2X1 port map( A => n514, B => readptr_2_port, Y => n816);
   U1194 : INVX1 port map( A => opcode_10_0_port, Y => n474);
   U1195 : AOI22X1 port map( A => n574, B => opcode_15_0_port, C => n575, D => 
                           opcode_14_0_port, Y => n845);
   U1196 : NOR2X1 port map( A => n514, B => n851, Y => n817);
   U1197 : AOI22X1 port map( A => n576, B => opcode_13_0_port, C => n577, D => 
                           opcode_12_0_port, Y => n844);
   U1198 : INVX1 port map( A => n852, Y => n850);
   U1199 : NAND3X1 port map( A => n820, B => n842, C => readptr_3_port, Y => 
                           n852);
   U1200 : INVX1 port map( A => readptr_0_port, Y => n820);
   U1201 : NOR2X1 port map( A => n851, B => readptr_1_port, Y => n818);
   U1202 : INVX1 port map( A => readptr_2_port, Y => n851);
   U1203 : INVX1 port map( A => n853, Y => n849);
   U1204 : NAND3X1 port map( A => readptr_0_port, B => n842, C => 
                           readptr_3_port, Y => n853);
   U1205 : INVX1 port map( A => readptr_4_port, Y => n842);
   U1207 : AND2X1 port map( A => N337, B => n72, Y => N347);
   U1208 : AND2X1 port map( A => N336, B => n72, Y => N346);
   U1209 : AND2X1 port map( A => N335, B => n72, Y => N345);
   U1210 : AND2X1 port map( A => N334, B => n72, Y => N344);
   U1211 : AND2X1 port map( A => N333, B => n72, Y => N343);
   U1212 : AND2X1 port map( A => N193, B => n72, Y => N342);
   U1213 : AND2X1 port map( A => N192, B => n72, Y => N341);
   U1214 : AND2X1 port map( A => N191, B => n72, Y => N340);
   U1215 : AND2X1 port map( A => N190, B => n72, Y => N339);
   U1216 : AND2X1 port map( A => N189, B => n72, Y => N338);
   U1217 : AND2X1 port map( A => R_ENABLE, B => n304, Y => N195);
   U1218 : NAND3X1 port map( A => n855, B => n857, C => n859, Y => n304);
   U1219 : NOR2X1 port map( A => n861, B => n863, Y => n859);
   U1220 : XOR2X1 port map( A => writeptr_4_port, B => readptr_4_port, Y => 
                           n863);
   U1221 : XOR2X1 port map( A => n71, B => readptr_3_port, Y => n861);
   U1222 : XOR2X1 port map( A => n514, B => n67, Y => n857);
   U1223 : INVX1 port map( A => readptr_1_port, Y => n514);
   U1224 : NOR2X1 port map( A => n864, B => n865, Y => n855);
   U1225 : XOR2X1 port map( A => n69, B => readptr_0_port, Y => n865);
   U1226 : XOR2X1 port map( A => n65, B => readptr_2_port, Y => n864);

end SYN_BRFIFO;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RBUFFER_1 is

   port( CLK, RST, NEXT_BYTE : in std_logic;  DATA : in std_logic_vector (7 
         downto 0);  OPCODE : in std_logic_vector (1 downto 0);  BYTE_COUNT : 
         in std_logic_vector (4 downto 0);  EOP : in std_logic;  B_READY, 
         R_ENABLE : out std_logic;  PRGA_IN : out std_logic_vector (7 downto 0)
         ;  PRGA_OPCODE : out std_logic_vector (1 downto 0));

end RBUFFER_1;

architecture SYN_brbuffer of RBUFFER_1 is

   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal B_READY_port, R_ENABLE_port, PRGA_IN_7_port, PRGA_IN_6_port, 
      PRGA_IN_5_port, PRGA_IN_4_port, PRGA_IN_3_port, PRGA_IN_2_port, 
      PRGA_IN_1_port, PRGA_IN_0_port, PRGA_OPCODE_1_port, PRGA_OPCODE_0_port, 
      state_2_port, state_1_port, state_0_port, nextState_2_port, 
      nextState_1_port, nextState_0_port, tempData_7_port, tempData_6_port, 
      tempData_5_port, tempData_4_port, tempData_3_port, tempData_2_port, 
      tempData_1_port, tempData_0_port, tempOpcode_1_port, tempOpcode_0_port, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n97, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n86, n88, 
      n89, n90, n91 : std_logic;

begin
   B_READY <= B_READY_port;
   R_ENABLE <= R_ENABLE_port;
   PRGA_IN <= ( PRGA_IN_7_port, PRGA_IN_6_port, PRGA_IN_5_port, PRGA_IN_4_port,
      PRGA_IN_3_port, PRGA_IN_2_port, PRGA_IN_1_port, PRGA_IN_0_port );
   PRGA_OPCODE <= ( PRGA_OPCODE_1_port, PRGA_OPCODE_0_port );
   
   B_READY_reg : DFFPOSX1 port map( D => n97, CLK => CLK, Q => B_READY_port);
   tempData_reg_7_inst : DFFPOSX1 port map( D => n71, CLK => CLK, Q => 
                           tempData_7_port);
   tempData_reg_6_inst : DFFPOSX1 port map( D => n72, CLK => CLK, Q => 
                           tempData_6_port);
   tempData_reg_5_inst : DFFPOSX1 port map( D => n73, CLK => CLK, Q => 
                           tempData_5_port);
   tempData_reg_4_inst : DFFPOSX1 port map( D => n74, CLK => CLK, Q => 
                           tempData_4_port);
   tempData_reg_3_inst : DFFPOSX1 port map( D => n75, CLK => CLK, Q => 
                           tempData_3_port);
   tempData_reg_2_inst : DFFPOSX1 port map( D => n86, CLK => CLK, Q => 
                           tempData_2_port);
   tempData_reg_1_inst : DFFPOSX1 port map( D => n88, CLK => CLK, Q => 
                           tempData_1_port);
   tempData_reg_0_inst : DFFPOSX1 port map( D => n89, CLK => CLK, Q => 
                           tempData_0_port);
   tempOpcode_reg_1_inst : DFFPOSX1 port map( D => n90, CLK => CLK, Q => 
                           tempOpcode_1_port);
   PRGA_OPCODE_reg_1_inst : DFFPOSX1 port map( D => n87, CLK => CLK, Q => 
                           PRGA_OPCODE_1_port);
   tempOpcode_reg_0_inst : DFFPOSX1 port map( D => n91, CLK => CLK, Q => 
                           tempOpcode_0_port);
   PRGA_OPCODE_reg_0_inst : DFFPOSX1 port map( D => n85, CLK => CLK, Q => 
                           PRGA_OPCODE_0_port);
   R_ENABLE_reg : DFFPOSX1 port map( D => n84, CLK => CLK, Q => R_ENABLE_port);
   PRGA_IN_reg_7_inst : DFFPOSX1 port map( D => n83, CLK => CLK, Q => 
                           PRGA_IN_7_port);
   PRGA_IN_reg_6_inst : DFFPOSX1 port map( D => n82, CLK => CLK, Q => 
                           PRGA_IN_6_port);
   PRGA_IN_reg_5_inst : DFFPOSX1 port map( D => n81, CLK => CLK, Q => 
                           PRGA_IN_5_port);
   PRGA_IN_reg_4_inst : DFFPOSX1 port map( D => n80, CLK => CLK, Q => 
                           PRGA_IN_4_port);
   PRGA_IN_reg_3_inst : DFFPOSX1 port map( D => n79, CLK => CLK, Q => 
                           PRGA_IN_3_port);
   PRGA_IN_reg_2_inst : DFFPOSX1 port map( D => n78, CLK => CLK, Q => 
                           PRGA_IN_2_port);
   PRGA_IN_reg_1_inst : DFFPOSX1 port map( D => n77, CLK => CLK, Q => 
                           PRGA_IN_1_port);
   PRGA_IN_reg_0_inst : DFFPOSX1 port map( D => n76, CLK => CLK, Q => 
                           PRGA_IN_0_port);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n4, S => n3, Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n4, S => n2, Q => state_2_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n4, S => n1, Q => state_0_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   U6 : INVX2 port map( A => n44, Y => n31);
   U7 : INVX2 port map( A => RST, Y => n4);
   U8 : OR2X2 port map( A => n42, B => RST, Y => n32);
   U9 : AND2X2 port map( A => n42, B => n4, Y => n47);
   U10 : OAI21X1 port map( A => n5, B => n6, C => n7, Y => nextState_2_port);
   U11 : MUX2X1 port map( B => n8, A => n9, S => state_0_port, Y => n7);
   U12 : NOR2X1 port map( A => state_2_port, B => n10, Y => n9);
   U13 : AND2X1 port map( A => state_2_port, B => n11, Y => n8);
   U14 : OAI21X1 port map( A => NEXT_BYTE, B => n12, C => state_1_port, Y => 
                           n11);
   U15 : AND2X1 port map( A => n13, B => NEXT_BYTE, Y => n5);
   U16 : OAI21X1 port map( A => state_2_port, B => n14, C => n15, Y => 
                           nextState_1_port);
   U17 : OAI21X1 port map( A => n16, B => n17, C => n18, Y => n15);
   U18 : INVX1 port map( A => n6, Y => n17);
   U19 : OAI21X1 port map( A => state_2_port, B => n19, C => n20, Y => 
                           nextState_0_port);
   U20 : AOI22X1 port map( A => n21, B => n22, C => NEXT_BYTE, D => n23, Y => 
                           n20);
   U21 : OAI21X1 port map( A => n13, B => n6, C => n24, Y => n23);
   U22 : INVX1 port map( A => n16, Y => n24);
   U23 : NOR2X1 port map( A => n19, B => n12, Y => n16);
   U24 : NOR2X1 port map( A => n25, B => BYTE_COUNT(4), Y => n12);
   U25 : NAND3X1 port map( A => state_0_port, B => n10, C => state_2_port, Y =>
                           n6);
   U26 : AND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n13);
   U27 : OAI21X1 port map( A => n26, B => n18, C => n27, Y => n22);
   U28 : INVX1 port map( A => NEXT_BYTE, Y => n18);
   U29 : AOI21X1 port map( A => EOP, B => n25, C => BYTE_COUNT(4), Y => n26);
   U30 : NAND2X1 port map( A => n28, B => n29, Y => n25);
   U31 : NOR2X1 port map( A => BYTE_COUNT(3), B => BYTE_COUNT(2), Y => n29);
   U32 : NOR2X1 port map( A => BYTE_COUNT(1), B => BYTE_COUNT(0), Y => n28);
   U33 : NOR2X1 port map( A => state_1_port, B => state_0_port, Y => n21);
   U34 : INVX1 port map( A => n30, Y => n71);
   U35 : AOI22X1 port map( A => n31, B => DATA(7), C => n32, D => 
                           tempData_7_port, Y => n30);
   U36 : INVX1 port map( A => n33, Y => n72);
   U37 : AOI22X1 port map( A => n31, B => DATA(6), C => n32, D => 
                           tempData_6_port, Y => n33);
   U38 : INVX1 port map( A => n34, Y => n73);
   U39 : AOI22X1 port map( A => n31, B => DATA(5), C => n32, D => 
                           tempData_5_port, Y => n34);
   U40 : INVX1 port map( A => n35, Y => n74);
   U41 : AOI22X1 port map( A => n31, B => DATA(4), C => n32, D => 
                           tempData_4_port, Y => n35);
   U42 : INVX1 port map( A => n36, Y => n75);
   U43 : AOI22X1 port map( A => n31, B => DATA(3), C => n32, D => 
                           tempData_3_port, Y => n36);
   U44 : INVX1 port map( A => n37, Y => n86);
   U45 : AOI22X1 port map( A => n31, B => DATA(2), C => n32, D => 
                           tempData_2_port, Y => n37);
   U46 : INVX1 port map( A => n38, Y => n88);
   U47 : AOI22X1 port map( A => n31, B => DATA(1), C => n32, D => 
                           tempData_1_port, Y => n38);
   U48 : INVX1 port map( A => n39, Y => n89);
   U49 : AOI22X1 port map( A => n31, B => DATA(0), C => n32, D => 
                           tempData_0_port, Y => n39);
   U50 : INVX1 port map( A => n40, Y => n90);
   U51 : AOI22X1 port map( A => OPCODE(1), B => n31, C => n32, D => 
                           tempOpcode_1_port, Y => n40);
   U52 : INVX1 port map( A => n41, Y => n91);
   U53 : AOI22X1 port map( A => OPCODE(0), B => n31, C => n32, D => 
                           tempOpcode_0_port, Y => n41);
   U54 : OAI21X1 port map( A => n4, B => n43, C => n44, Y => n97);
   U55 : INVX1 port map( A => B_READY_port, Y => n43);
   U56 : OAI21X1 port map( A => n4, B => n45, C => n46, Y => n87);
   U57 : AOI22X1 port map( A => n31, B => OPCODE(1), C => n47, D => 
                           tempOpcode_1_port, Y => n46);
   U58 : INVX1 port map( A => PRGA_OPCODE_1_port, Y => n45);
   U59 : OAI21X1 port map( A => n4, B => n48, C => n49, Y => n85);
   U60 : AOI22X1 port map( A => n31, B => OPCODE(0), C => n47, D => 
                           tempOpcode_0_port, Y => n49);
   U61 : INVX1 port map( A => PRGA_OPCODE_0_port, Y => n48);
   U62 : MUX2X1 port map( B => n50, A => n51, S => RST, Y => n84);
   U63 : INVX1 port map( A => R_ENABLE_port, Y => n51);
   U64 : NAND3X1 port map( A => n10, B => n27, C => state_0_port, Y => n50);
   U65 : OAI21X1 port map( A => n4, B => n52, C => n53, Y => n83);
   U66 : AOI22X1 port map( A => DATA(7), B => n31, C => n47, D => 
                           tempData_7_port, Y => n53);
   U67 : INVX1 port map( A => PRGA_IN_7_port, Y => n52);
   U68 : OAI21X1 port map( A => n4, B => n54, C => n55, Y => n82);
   U69 : AOI22X1 port map( A => DATA(6), B => n31, C => n47, D => 
                           tempData_6_port, Y => n55);
   U70 : INVX1 port map( A => PRGA_IN_6_port, Y => n54);
   U71 : OAI21X1 port map( A => n4, B => n56, C => n57, Y => n81);
   U72 : AOI22X1 port map( A => DATA(5), B => n31, C => n47, D => 
                           tempData_5_port, Y => n57);
   U73 : INVX1 port map( A => PRGA_IN_5_port, Y => n56);
   U74 : OAI21X1 port map( A => n4, B => n58, C => n59, Y => n80);
   U75 : AOI22X1 port map( A => DATA(4), B => n31, C => n47, D => 
                           tempData_4_port, Y => n59);
   U76 : INVX1 port map( A => PRGA_IN_4_port, Y => n58);
   U77 : OAI21X1 port map( A => n4, B => n60, C => n61, Y => n79);
   U78 : AOI22X1 port map( A => DATA(3), B => n31, C => n47, D => 
                           tempData_3_port, Y => n61);
   U79 : INVX1 port map( A => PRGA_IN_3_port, Y => n60);
   U80 : OAI21X1 port map( A => n4, B => n62, C => n63, Y => n78);
   U81 : AOI22X1 port map( A => DATA(2), B => n31, C => n47, D => 
                           tempData_2_port, Y => n63);
   U82 : INVX1 port map( A => PRGA_IN_2_port, Y => n62);
   U83 : OAI21X1 port map( A => n4, B => n64, C => n65, Y => n77);
   U84 : AOI22X1 port map( A => DATA(1), B => n31, C => n47, D => 
                           tempData_1_port, Y => n65);
   U85 : INVX1 port map( A => PRGA_IN_1_port, Y => n64);
   U86 : OAI21X1 port map( A => n4, B => n66, C => n67, Y => n76);
   U87 : AOI22X1 port map( A => DATA(0), B => n31, C => n47, D => 
                           tempData_0_port, Y => n67);
   U88 : NAND2X1 port map( A => n14, B => state_2_port, Y => n42);
   U89 : INVX1 port map( A => n68, Y => n14);
   U90 : OAI21X1 port map( A => state_1_port, B => n69, C => n19, Y => n68);
   U91 : NAND2X1 port map( A => state_1_port, B => n69, Y => n19);
   U92 : NAND3X1 port map( A => n69, B => n10, C => n70, Y => n44);
   U93 : NOR2X1 port map( A => RST, B => n27, Y => n70);
   U94 : INVX1 port map( A => state_2_port, Y => n27);
   U95 : INVX1 port map( A => state_1_port, Y => n10);
   U96 : INVX1 port map( A => state_0_port, Y => n69);
   U97 : INVX1 port map( A => PRGA_IN_0_port, Y => n66);

end SYN_brbuffer;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity uart_rcv_block_1 is

   port( CLK, RST, SERIAL_IN : in std_logic;  KEY_ERROR, PROG_ERROR : out 
         std_logic;  PLAINKEY : out std_logic_vector (63 downto 0);  RBUF_FULL,
         PARITY_ERROR : out std_logic);

end uart_rcv_block_1;

architecture SYN_struct1 of uart_rcv_block_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component uart_timer_1
      port( CLK, RST, TIMER_TRIG : in std_logic;  STOP_RCVING, SHIFT_STROBE : 
            out std_logic);
   end component;
   
   component keyreg_1
      port( CLK, RST, SBE, OE, RBUF_FULL : in std_logic;  RCV_DATA : in 
            std_logic_vector (7 downto 0);  PLAINKEY : out std_logic_vector (63
            downto 0);  KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR : out 
            std_logic);
   end component;
   
   component uart_sr_10bit_1
      port( CLK, RST, SHIFT_STROBE, SERIAL_IN : in std_logic;  LOAD_DATA : out 
            std_logic_vector (7 downto 0);  STOP_DATA : out std_logic_vector (1
            downto 0));
   end component;
   
   component uart_sb_check_1
      port( RST, CLK, SBC_CLR, SBC_EN : in std_logic;  STOP_DATA : in 
            std_logic_vector (1 downto 0);  SB_DETECT, SBE : out std_logic);
   end component;
   
   component uart_rcv_buf_full_1
      port( CLK, RST, CLR_RBUF, SET_RBUF_FULL : in std_logic;  RBUF_FULL : out 
            std_logic);
   end component;
   
   component uart_rcv_buf_1
      port( CLK, RST, LOAD_RBUF : in std_logic;  LOAD_DATA : in 
            std_logic_vector (7 downto 0);  RCV_DATA : out std_logic_vector (7 
            downto 0));
   end component;
   
   component uart_rcu_1
      port( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT : in std_logic;  
            RBUF_LOAD, TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR : 
            out std_logic);
   end component;
   
   component uart_error_1
      port( RST, CLK, RBUF_FULL, CHK_ERROR : in std_logic;  OE : out std_logic
            );
   end component;
   
   component uart_edge_detector_1
      port( CLK, RST, SERIAL_IN : in std_logic;  START_BIT : out std_logic);
   end component;
   
   signal RBUF_FULL_port, START_BIT, CHK_ERROR, OE, SB_DETECT, STOP_RCVING, 
      RBUF_LOAD, SBC_CLR, SBC_EN, SET_RBUF_FULL, TIMER_TRIG, LOAD_DATA_7_port, 
      LOAD_DATA_6_port, LOAD_DATA_5_port, LOAD_DATA_4_port, LOAD_DATA_3_port, 
      LOAD_DATA_2_port, LOAD_DATA_1_port, LOAD_DATA_0_port, RCV_DATA_7_port, 
      RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, RCV_DATA_3_port, 
      RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, CLR_RBUF, 
      STOP_DATA_1_port, STOP_DATA_0_port, SBE, SHIFT_STROBE, n1, n2 : std_logic
      ;

begin
   RBUF_FULL <= RBUF_FULL_port;
   
   U_0 : uart_edge_detector_1 port map( CLK => CLK, RST => n1, SERIAL_IN => 
                           SERIAL_IN, START_BIT => START_BIT);
   U_1 : uart_error_1 port map( RST => n1, CLK => CLK, RBUF_FULL => 
                           RBUF_FULL_port, CHK_ERROR => CHK_ERROR, OE => OE);
   U_2 : uart_rcu_1 port map( CLK => CLK, RST => n1, START_BIT => START_BIT, 
                           STOP_RCVING => STOP_RCVING, SB_DETECT => SB_DETECT, 
                           RBUF_LOAD => RBUF_LOAD, TIMER_TRIG => TIMER_TRIG, 
                           CHK_ERROR => CHK_ERROR, SET_RBUF_FULL => 
                           SET_RBUF_FULL, SBC_EN => SBC_EN, SBC_CLR => SBC_CLR)
                           ;
   U_3 : uart_rcv_buf_1 port map( CLK => CLK, RST => n1, LOAD_RBUF => RBUF_LOAD
                           , LOAD_DATA(7) => LOAD_DATA_7_port, LOAD_DATA(6) => 
                           LOAD_DATA_6_port, LOAD_DATA(5) => LOAD_DATA_5_port, 
                           LOAD_DATA(4) => LOAD_DATA_4_port, LOAD_DATA(3) => 
                           LOAD_DATA_3_port, LOAD_DATA(2) => LOAD_DATA_2_port, 
                           LOAD_DATA(1) => LOAD_DATA_1_port, LOAD_DATA(0) => 
                           LOAD_DATA_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port);
   U_4 : uart_rcv_buf_full_1 port map( CLK => CLK, RST => n1, CLR_RBUF => 
                           CLR_RBUF, SET_RBUF_FULL => SET_RBUF_FULL, RBUF_FULL 
                           => RBUF_FULL_port);
   U_5 : uart_sb_check_1 port map( RST => n1, CLK => CLK, SBC_CLR => SBC_CLR, 
                           SBC_EN => SBC_EN, STOP_DATA(1) => STOP_DATA_1_port, 
                           STOP_DATA(0) => STOP_DATA_0_port, SB_DETECT => 
                           SB_DETECT, SBE => SBE);
   U_6 : uart_sr_10bit_1 port map( CLK => CLK, RST => n1, SHIFT_STROBE => 
                           SHIFT_STROBE, SERIAL_IN => SERIAL_IN, LOAD_DATA(7) 
                           => LOAD_DATA_7_port, LOAD_DATA(6) => 
                           LOAD_DATA_6_port, LOAD_DATA(5) => LOAD_DATA_5_port, 
                           LOAD_DATA(4) => LOAD_DATA_4_port, LOAD_DATA(3) => 
                           LOAD_DATA_3_port, LOAD_DATA(2) => LOAD_DATA_2_port, 
                           LOAD_DATA(1) => LOAD_DATA_1_port, LOAD_DATA(0) => 
                           LOAD_DATA_0_port, STOP_DATA(1) => STOP_DATA_1_port, 
                           STOP_DATA(0) => STOP_DATA_0_port);
   U_8 : keyreg_1 port map( CLK => CLK, RST => n1, SBE => SBE, OE => OE, 
                           RBUF_FULL => RBUF_FULL_port, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           PLAINKEY(63) => PLAINKEY(63), PLAINKEY(62) => 
                           PLAINKEY(62), PLAINKEY(61) => PLAINKEY(61), 
                           PLAINKEY(60) => PLAINKEY(60), PLAINKEY(59) => 
                           PLAINKEY(59), PLAINKEY(58) => PLAINKEY(58), 
                           PLAINKEY(57) => PLAINKEY(57), PLAINKEY(56) => 
                           PLAINKEY(56), PLAINKEY(55) => PLAINKEY(55), 
                           PLAINKEY(54) => PLAINKEY(54), PLAINKEY(53) => 
                           PLAINKEY(53), PLAINKEY(52) => PLAINKEY(52), 
                           PLAINKEY(51) => PLAINKEY(51), PLAINKEY(50) => 
                           PLAINKEY(50), PLAINKEY(49) => PLAINKEY(49), 
                           PLAINKEY(48) => PLAINKEY(48), PLAINKEY(47) => 
                           PLAINKEY(47), PLAINKEY(46) => PLAINKEY(46), 
                           PLAINKEY(45) => PLAINKEY(45), PLAINKEY(44) => 
                           PLAINKEY(44), PLAINKEY(43) => PLAINKEY(43), 
                           PLAINKEY(42) => PLAINKEY(42), PLAINKEY(41) => 
                           PLAINKEY(41), PLAINKEY(40) => PLAINKEY(40), 
                           PLAINKEY(39) => PLAINKEY(39), PLAINKEY(38) => 
                           PLAINKEY(38), PLAINKEY(37) => PLAINKEY(37), 
                           PLAINKEY(36) => PLAINKEY(36), PLAINKEY(35) => 
                           PLAINKEY(35), PLAINKEY(34) => PLAINKEY(34), 
                           PLAINKEY(33) => PLAINKEY(33), PLAINKEY(32) => 
                           PLAINKEY(32), PLAINKEY(31) => PLAINKEY(31), 
                           PLAINKEY(30) => PLAINKEY(30), PLAINKEY(29) => 
                           PLAINKEY(29), PLAINKEY(28) => PLAINKEY(28), 
                           PLAINKEY(27) => PLAINKEY(27), PLAINKEY(26) => 
                           PLAINKEY(26), PLAINKEY(25) => PLAINKEY(25), 
                           PLAINKEY(24) => PLAINKEY(24), PLAINKEY(23) => 
                           PLAINKEY(23), PLAINKEY(22) => PLAINKEY(22), 
                           PLAINKEY(21) => PLAINKEY(21), PLAINKEY(20) => 
                           PLAINKEY(20), PLAINKEY(19) => PLAINKEY(19), 
                           PLAINKEY(18) => PLAINKEY(18), PLAINKEY(17) => 
                           PLAINKEY(17), PLAINKEY(16) => PLAINKEY(16), 
                           PLAINKEY(15) => PLAINKEY(15), PLAINKEY(14) => 
                           PLAINKEY(14), PLAINKEY(13) => PLAINKEY(13), 
                           PLAINKEY(12) => PLAINKEY(12), PLAINKEY(11) => 
                           PLAINKEY(11), PLAINKEY(10) => PLAINKEY(10), 
                           PLAINKEY(9) => PLAINKEY(9), PLAINKEY(8) => 
                           PLAINKEY(8), PLAINKEY(7) => PLAINKEY(7), PLAINKEY(6)
                           => PLAINKEY(6), PLAINKEY(5) => PLAINKEY(5), 
                           PLAINKEY(4) => PLAINKEY(4), PLAINKEY(3) => 
                           PLAINKEY(3), PLAINKEY(2) => PLAINKEY(2), PLAINKEY(1)
                           => PLAINKEY(1), PLAINKEY(0) => PLAINKEY(0), 
                           KEY_ERROR => KEY_ERROR, PROG_ERROR => PROG_ERROR, 
                           CLR_RBUFF => CLR_RBUF, PARITY_ERROR => PARITY_ERROR)
                           ;
   U_7 : uart_timer_1 port map( CLK => CLK, RST => n1, TIMER_TRIG => TIMER_TRIG
                           , STOP_RCVING => STOP_RCVING, SHIFT_STROBE => 
                           SHIFT_STROBE);
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct1;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity KSA_1 is

   port( KEY : in std_logic_vector (63 downto 0);  CLK, RST, KEY_ERROR, 
         BYTE_READY : in std_logic;  BYTE : in std_logic_vector (7 downto 0);  
         OPCODE : in std_logic_vector (1 downto 0);  DATA_IN : in 
         std_logic_vector (7 downto 0);  PROCESSED_DATA : out std_logic_vector 
         (7 downto 0);  PDATA_READY, W_ENABLE, R_ENABLE : out std_logic;  ADDR,
         DATA : out std_logic_vector (7 downto 0));

end KSA_1;

architecture SYN_bksa of KSA_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUFX1
      port( A, EN : in std_logic;  Y : out std_logic);
   end component;
   
   component KSA_1_DW01_add_2
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_1_DW01_add_3
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_1_DW01_inc_2
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_1_DW01_inc_1
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_1_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component KSA_1_DW01_add_1
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component KSA_1_DW01_add_0
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, PROCESSED_DATA_5_port, 
      PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, PROCESSED_DATA_2_port, 
      PROCESSED_DATA_1_port, PROCESSED_DATA_0_port, W_ENABLE_port, 
      R_ENABLE_port, ADDR_7_port, ADDR_6_port, ADDR_5_port, ADDR_4_port, 
      ADDR_3_port, ADDR_2_port, ADDR_1_port, ADDR_0_port, DATA_7_port, 
      DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, DATA_2_port, 
      DATA_1_port, DATA_0_port, state_4_port, state_3_port, state_2_port, 
      state_1_port, state_0_port, si_7_port, si_6_port, si_5_port, si_4_port, 
      si_3_port, si_2_port, si_1_port, si_0_port, sj_7_port, sj_6_port, 
      sj_5_port, sj_4_port, sj_3_port, sj_2_port, sj_1_port, sj_0_port, 
      currentProcessedData_7_port, currentProcessedData_6_port, 
      currentProcessedData_5_port, currentProcessedData_4_port, 
      currentProcessedData_3_port, currentProcessedData_2_port, 
      currentProcessedData_1_port, currentProcessedData_0_port, 
      nextState_4_port, nextState_3_port, nextState_2_port, nextState_1_port, 
      nextState_0_port, inti_7_port, inti_6_port, inti_5_port, inti_4_port, 
      inti_3_port, inti_2_port, inti_1_port, inti_0_port, intj_7_port, 
      intj_6_port, intj_5_port, intj_4_port, intj_3_port, intj_2_port, 
      intj_1_port, intj_0_port, keyi_2_port, keyi_1_port, keyi_0_port, 
      permuteComplete, temp_7_port, temp_6_port, temp_5_port, temp_4_port, 
      temp_3_port, temp_2_port, temp_1_port, temp_0_port, extratemp_7_port, 
      extratemp_6_port, extratemp_5_port, extratemp_4_port, extratemp_3_port, 
      extratemp_2_port, extratemp_1_port, extratemp_0_port, 
      nextProcessedData_7_port, nextProcessedData_6_port, 
      nextProcessedData_5_port, nextProcessedData_4_port, 
      nextProcessedData_3_port, nextProcessedData_2_port, 
      nextProcessedData_1_port, nextProcessedData_0_port, keyTable_0_7_port, 
      keyTable_0_6_port, keyTable_0_5_port, keyTable_0_4_port, 
      keyTable_0_3_port, keyTable_0_2_port, keyTable_0_1_port, 
      keyTable_0_0_port, keyTable_1_7_port, keyTable_1_6_port, 
      keyTable_1_5_port, keyTable_1_4_port, keyTable_1_3_port, 
      keyTable_1_2_port, keyTable_1_1_port, keyTable_1_0_port, 
      keyTable_2_7_port, keyTable_2_6_port, keyTable_2_5_port, 
      keyTable_2_4_port, keyTable_2_3_port, keyTable_2_2_port, 
      keyTable_2_1_port, keyTable_2_0_port, keyTable_3_7_port, 
      keyTable_3_6_port, keyTable_3_5_port, keyTable_3_4_port, 
      keyTable_3_3_port, keyTable_3_2_port, keyTable_3_1_port, 
      keyTable_3_0_port, keyTable_4_7_port, keyTable_4_6_port, 
      keyTable_4_5_port, keyTable_4_4_port, keyTable_4_3_port, 
      keyTable_4_2_port, keyTable_4_1_port, keyTable_4_0_port, 
      keyTable_5_7_port, keyTable_5_6_port, keyTable_5_5_port, 
      keyTable_5_4_port, keyTable_5_3_port, keyTable_5_2_port, 
      keyTable_5_1_port, keyTable_5_0_port, keyTable_6_7_port, 
      keyTable_6_6_port, keyTable_6_5_port, keyTable_6_4_port, 
      keyTable_6_3_port, keyTable_6_2_port, keyTable_6_1_port, 
      keyTable_6_0_port, keyTable_7_7_port, keyTable_7_6_port, 
      keyTable_7_5_port, keyTable_7_4_port, keyTable_7_3_port, 
      keyTable_7_2_port, keyTable_7_1_port, keyTable_7_0_port, delaydata_7_port
      , delaydata_6_port, delaydata_5_port, delaydata_4_port, delaydata_3_port,
      delaydata_2_port, delaydata_1_port, delaydata_0_port, 
      prefillCounter_7_port, prefillCounter_6_port, prefillCounter_5_port, 
      prefillCounter_4_port, prefillCounter_3_port, prefillCounter_2_port, 
      prefillCounter_1_port, prefillCounter_0_port, faddr_7_port, faddr_6_port,
      faddr_5_port, faddr_4_port, faddr_3_port, faddr_2_port, faddr_1_port, 
      faddr_0_port, nfaddr_7_port, nfaddr_6_port, nfaddr_5_port, nfaddr_4_port,
      nfaddr_3_port, nfaddr_2_port, nfaddr_1_port, nfaddr_0_port, fdata_7_port,
      fdata_6_port, fdata_5_port, fdata_4_port, fdata_3_port, fdata_2_port, 
      fdata_1_port, fdata_0_port, nfdata_7_port, nfdata_6_port, nfdata_5_port, 
      nfdata_4_port, nfdata_3_port, nfdata_2_port, nfdata_1_port, nfdata_0_port
      , fw_enable, fr_enable, N407, N408, N409, N410, N411, N412, N413, N414, 
      N424, N425, N426, N427, N428, N429, N430, N431, N442, N443, N444, N445, 
      N446, N447, N448, N472, N473, N474, N475, N476, N477, N478, N479, N480, 
      N481, N482, N483, N484, N485, N486, N487, N496, N497, N498, N499, N500, 
      N501, N502, N503, N512, N513, N514, N515, N516, N517, N518, N519, N520, 
      N521, N522, N523, N524, N525, N526, N527, n1, n2, n11, n13, n18, n21, n23
      , n25, n26, n28, n30, n31, n33, n35, n36, n38, n40, n41, n43, n45, n46, 
      n48, n50, n51, n53, n55, n56, n57, n58, n59, n60, n61, n63, n65, n66, n67
      , n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n118, n119, n120, n123, n124, 
      n125, n126, n127, n128, n130, n132, n133, n134, n137, n138, n139, n140, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n152, n153, n154, 
      n155, n156, n157, n158, n159, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n173, n174, n176, n178, n179, n181, n182, n183, n184, 
      n186, n189, n190, n191, n192, n193, n194, n195, n197, n198, n199, n200, 
      n202, n204, n205, n207, n209, n211, n213, n215, n217, n219, n221, n222, 
      n223, n224, n225, n226, n227, n229, n231, n232, n233, n234, n236, n242, 
      n243, n245, n248, n251, n254, n257, n260, n263, n266, n269, n272, n273, 
      n274, n276, n278, n279, n281, n283, n284, n286, n288, n289, n291, n293, 
      n294, n296, n298, n299, n301, n303, n304, n306, n308, n309, n310, n312, 
      n313, n314, n315, n316, n319, n320, n321, n322, n323, n324, n325, n328, 
      n330, n332, n334, n336, n338, n340, n342, n344, n346, n348, n350, n352, 
      n354, n356, n358, n360, n362, n364, n366, n368, n370, n372, n374, n376, 
      n378, n380, n382, n384, n386, n388, n390, n392, n394, n396, n398, n400, 
      n402, n404, n406, n408_port, n410_port, n412_port, n414_port, n416, n418,
      n420, n422, n424_port, n426_port, n428_port, n430_port, n432, n434, n436,
      n438, n440, n442_port, n444_port, n446_port, n448_port, n450, n452, n454,
      n456, n457, n460, n464, n466, n468, n470, n472_port, n474_port, n476_port
      , n477_port, n478_port, n479_port, n481_port, n483_port, n484_port, 
      n485_port, n486_port, n487_port, n489, n490, n491, n492, n493, n494, n495
      , n496_port, n497_port, n499_port, n502_port, n508, n510, n511, n513_port
      , n515_port, n517_port, n519_port, n521_port, n523_port, n525_port, 
      n526_port, n527_port, n529, n530, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n544, n546, n548, n550, n552, n554, n556, n558, n559, 
      n560, n561, n563, n564, n565, n566, n567, n568, n570, n573, n574, n576, 
      n578, n580, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n593, n595, n596, n597, n598, n599, n601, n602, n603, n607, n608, n609, 
      n611, n613, n615, n617, n619, n620, n621, n622, n623, n625, n627, n628, 
      n631, n633, n634, n635, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n693, n694, n695, n696, n697, n698, n699, 
      n700, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n747, n749, n751, 
      n753, n755, n757, n759, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, N456_port, N455, N454_port, N453, N452_port, N451
      , N450_port, N449, n3, n4, n5, n6, n7, n8, n9, n10, n12, n14, n15, n16, 
      n17, n19, n20, n22, n24, n27, n29, n32, n34, n37, n39, n42, n44, n47, n49
      , n52, n54, n62, n64, n69, n117, n121, n122, n129, n131, n135, n136, n141
      , n151, n160, n161, n172, n175, n177, n180, n185, n187, n188, n196, n201,
      n203, n206, n208, n210, n212, n214, n216, n218, n220, n228, n230, n235, 
      n237, n238, n239, n240, n241, n244, n246, n247, n249, n250, n252, n253, 
      n255, n256, n258, n259, n261, n262, n264, n265, n267, n268, n270, n271, 
      n275, n277, n280, n282, n285, n287, n290, n292, n295, n297, n300, n302, 
      n305, n307, n311, n317, n318, n326, n327, n329, n331, n333, n335, n337, 
      n339, n341, n343, n345, n347, n349, n351, n353, n355, n357, n359, n361, 
      n363, n365, n367, n369, n371, n373, n375, n377, n379, n381, n383, n385, 
      n387, n389, n391, n393, n395, n397, n399, n401, n403, n405, n407_port, 
      n409_port, n411_port, n413_port, n415, n417, n419, n421, n423, n425_port,
      n427_port, n429_port, n431_port, n433, n435, n437, n439, n441, n443_port,
      n445_port, n447_port, n449_port, n451_port, n453_port, n455_port, n458, 
      n459, n461, n462, n463, n465, n467, n469, n471, n473_port, n475_port, 
      n480_port, n482_port, n488, n498_port, n500_port, n501_port, n503_port, 
      n504, n505, n506, n507, n509, n512_port, n514_port, n516_port, n518_port,
      n520_port, n522_port, n524_port, n528, n540, n541, n542, n543, n545, n547
      , n549, n551, n553, n555, n557, n562, n569, n571, n572, n575, n577, n579,
      n581, n592, n594, n600, n604, n605, n606, n610, n612, n614, n616, n618, 
      n624, n626, n629, n630, n632, n636, n637, n638, n648, n649, n650, n651, 
      n692, n701, n746, n748, n750, n752, n754, n756, n758, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n864, n865, n866, n867, n868, n869, n870, 
      n871, n883, n884, n885, n886, n887, n888, n889, n890, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n_1026,
      n_1027, n_1028, n_1029 : std_logic;

begin
   PROCESSED_DATA <= ( PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, 
      PROCESSED_DATA_5_port, PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, 
      PROCESSED_DATA_2_port, PROCESSED_DATA_1_port, PROCESSED_DATA_0_port );
   W_ENABLE <= W_ENABLE_port;
   R_ENABLE <= R_ENABLE_port;
   ADDR <= ( ADDR_7_port, ADDR_6_port, ADDR_5_port, ADDR_4_port, ADDR_3_port, 
      ADDR_2_port, ADDR_1_port, ADDR_0_port );
   DATA <= ( DATA_7_port, DATA_6_port, DATA_5_port, DATA_4_port, DATA_3_port, 
      DATA_2_port, DATA_1_port, DATA_0_port );
   
   n1 <= '0';
   n2 <= '0';
   prefillCounter_reg_0_inst : DFFPOSX1 port map( D => n915, CLK => CLK, Q => 
                           prefillCounter_0_port);
   permuteComplete_reg : DFFPOSX1 port map( D => n899, CLK => CLK, Q => 
                           permuteComplete);
   extratemp_reg_7_inst : DFFPOSX1 port map( D => n465, CLK => CLK, Q => 
                           extratemp_7_port);
   extratemp_reg_6_inst : DFFPOSX1 port map( D => n463, CLK => CLK, Q => 
                           extratemp_6_port);
   extratemp_reg_5_inst : DFFPOSX1 port map( D => n462, CLK => CLK, Q => 
                           extratemp_5_port);
   extratemp_reg_4_inst : DFFPOSX1 port map( D => n461, CLK => CLK, Q => 
                           extratemp_4_port);
   extratemp_reg_3_inst : DFFPOSX1 port map( D => n459, CLK => CLK, Q => 
                           extratemp_3_port);
   extratemp_reg_2_inst : DFFPOSX1 port map( D => n458, CLK => CLK, Q => 
                           extratemp_2_port);
   extratemp_reg_1_inst : DFFPOSX1 port map( D => n455_port, CLK => CLK, Q => 
                           extratemp_1_port);
   extratemp_reg_0_inst : DFFPOSX1 port map( D => n453_port, CLK => CLK, Q => 
                           extratemp_0_port);
   keyTable_reg_7_0_inst : DFFPOSX1 port map( D => n792, CLK => CLK, Q => 
                           keyTable_7_0_port);
   keyTable_reg_7_1_inst : DFFPOSX1 port map( D => n793, CLK => CLK, Q => 
                           keyTable_7_1_port);
   keyTable_reg_7_2_inst : DFFPOSX1 port map( D => n794, CLK => CLK, Q => 
                           keyTable_7_2_port);
   keyTable_reg_7_3_inst : DFFPOSX1 port map( D => n795, CLK => CLK, Q => 
                           keyTable_7_3_port);
   keyTable_reg_7_4_inst : DFFPOSX1 port map( D => n796, CLK => CLK, Q => 
                           keyTable_7_4_port);
   keyTable_reg_7_5_inst : DFFPOSX1 port map( D => n797, CLK => CLK, Q => 
                           keyTable_7_5_port);
   keyTable_reg_7_6_inst : DFFPOSX1 port map( D => n798, CLK => CLK, Q => 
                           keyTable_7_6_port);
   keyTable_reg_7_7_inst : DFFPOSX1 port map( D => n799, CLK => CLK, Q => 
                           keyTable_7_7_port);
   keyTable_reg_6_0_inst : DFFPOSX1 port map( D => n800, CLK => CLK, Q => 
                           keyTable_6_0_port);
   keyTable_reg_6_1_inst : DFFPOSX1 port map( D => n801, CLK => CLK, Q => 
                           keyTable_6_1_port);
   keyTable_reg_6_2_inst : DFFPOSX1 port map( D => n802, CLK => CLK, Q => 
                           keyTable_6_2_port);
   keyTable_reg_6_3_inst : DFFPOSX1 port map( D => n803, CLK => CLK, Q => 
                           keyTable_6_3_port);
   keyTable_reg_6_4_inst : DFFPOSX1 port map( D => n804, CLK => CLK, Q => 
                           keyTable_6_4_port);
   keyTable_reg_6_5_inst : DFFPOSX1 port map( D => n805, CLK => CLK, Q => 
                           keyTable_6_5_port);
   keyTable_reg_6_6_inst : DFFPOSX1 port map( D => n806, CLK => CLK, Q => 
                           keyTable_6_6_port);
   keyTable_reg_6_7_inst : DFFPOSX1 port map( D => n807, CLK => CLK, Q => 
                           keyTable_6_7_port);
   keyTable_reg_5_0_inst : DFFPOSX1 port map( D => n808, CLK => CLK, Q => 
                           keyTable_5_0_port);
   keyTable_reg_5_1_inst : DFFPOSX1 port map( D => n809, CLK => CLK, Q => 
                           keyTable_5_1_port);
   keyTable_reg_5_2_inst : DFFPOSX1 port map( D => n810, CLK => CLK, Q => 
                           keyTable_5_2_port);
   keyTable_reg_5_3_inst : DFFPOSX1 port map( D => n811, CLK => CLK, Q => 
                           keyTable_5_3_port);
   keyTable_reg_5_4_inst : DFFPOSX1 port map( D => n812, CLK => CLK, Q => 
                           keyTable_5_4_port);
   keyTable_reg_5_5_inst : DFFPOSX1 port map( D => n813, CLK => CLK, Q => 
                           keyTable_5_5_port);
   keyTable_reg_5_6_inst : DFFPOSX1 port map( D => n814, CLK => CLK, Q => 
                           keyTable_5_6_port);
   keyTable_reg_5_7_inst : DFFPOSX1 port map( D => n815, CLK => CLK, Q => 
                           keyTable_5_7_port);
   keyTable_reg_4_0_inst : DFFPOSX1 port map( D => n816, CLK => CLK, Q => 
                           keyTable_4_0_port);
   keyTable_reg_4_1_inst : DFFPOSX1 port map( D => n817, CLK => CLK, Q => 
                           keyTable_4_1_port);
   keyTable_reg_4_2_inst : DFFPOSX1 port map( D => n818, CLK => CLK, Q => 
                           keyTable_4_2_port);
   keyTable_reg_4_3_inst : DFFPOSX1 port map( D => n819, CLK => CLK, Q => 
                           keyTable_4_3_port);
   keyTable_reg_4_4_inst : DFFPOSX1 port map( D => n820, CLK => CLK, Q => 
                           keyTable_4_4_port);
   keyTable_reg_4_5_inst : DFFPOSX1 port map( D => n821, CLK => CLK, Q => 
                           keyTable_4_5_port);
   keyTable_reg_4_6_inst : DFFPOSX1 port map( D => n822, CLK => CLK, Q => 
                           keyTable_4_6_port);
   keyTable_reg_4_7_inst : DFFPOSX1 port map( D => n823, CLK => CLK, Q => 
                           keyTable_4_7_port);
   keyTable_reg_3_0_inst : DFFPOSX1 port map( D => n824, CLK => CLK, Q => 
                           keyTable_3_0_port);
   keyTable_reg_3_1_inst : DFFPOSX1 port map( D => n825, CLK => CLK, Q => 
                           keyTable_3_1_port);
   keyTable_reg_3_2_inst : DFFPOSX1 port map( D => n826, CLK => CLK, Q => 
                           keyTable_3_2_port);
   keyTable_reg_3_3_inst : DFFPOSX1 port map( D => n827, CLK => CLK, Q => 
                           keyTable_3_3_port);
   keyTable_reg_3_4_inst : DFFPOSX1 port map( D => n828, CLK => CLK, Q => 
                           keyTable_3_4_port);
   keyTable_reg_3_5_inst : DFFPOSX1 port map( D => n829, CLK => CLK, Q => 
                           keyTable_3_5_port);
   keyTable_reg_3_6_inst : DFFPOSX1 port map( D => n830, CLK => CLK, Q => 
                           keyTable_3_6_port);
   keyTable_reg_3_7_inst : DFFPOSX1 port map( D => n831, CLK => CLK, Q => 
                           keyTable_3_7_port);
   keyTable_reg_2_0_inst : DFFPOSX1 port map( D => n832, CLK => CLK, Q => 
                           keyTable_2_0_port);
   keyTable_reg_2_1_inst : DFFPOSX1 port map( D => n833, CLK => CLK, Q => 
                           keyTable_2_1_port);
   keyTable_reg_2_2_inst : DFFPOSX1 port map( D => n834, CLK => CLK, Q => 
                           keyTable_2_2_port);
   keyTable_reg_2_3_inst : DFFPOSX1 port map( D => n835, CLK => CLK, Q => 
                           keyTable_2_3_port);
   keyTable_reg_2_4_inst : DFFPOSX1 port map( D => n836, CLK => CLK, Q => 
                           keyTable_2_4_port);
   keyTable_reg_2_5_inst : DFFPOSX1 port map( D => n837, CLK => CLK, Q => 
                           keyTable_2_5_port);
   keyTable_reg_2_6_inst : DFFPOSX1 port map( D => n838, CLK => CLK, Q => 
                           keyTable_2_6_port);
   keyTable_reg_2_7_inst : DFFPOSX1 port map( D => n839, CLK => CLK, Q => 
                           keyTable_2_7_port);
   keyTable_reg_1_0_inst : DFFPOSX1 port map( D => n840, CLK => CLK, Q => 
                           keyTable_1_0_port);
   keyTable_reg_1_1_inst : DFFPOSX1 port map( D => n841, CLK => CLK, Q => 
                           keyTable_1_1_port);
   keyTable_reg_1_2_inst : DFFPOSX1 port map( D => n842, CLK => CLK, Q => 
                           keyTable_1_2_port);
   keyTable_reg_1_3_inst : DFFPOSX1 port map( D => n843, CLK => CLK, Q => 
                           keyTable_1_3_port);
   keyTable_reg_1_4_inst : DFFPOSX1 port map( D => n844, CLK => CLK, Q => 
                           keyTable_1_4_port);
   keyTable_reg_1_5_inst : DFFPOSX1 port map( D => n845, CLK => CLK, Q => 
                           keyTable_1_5_port);
   keyTable_reg_1_6_inst : DFFPOSX1 port map( D => n846, CLK => CLK, Q => 
                           keyTable_1_6_port);
   keyTable_reg_0_6_inst : DFFPOSX1 port map( D => n847, CLK => CLK, Q => 
                           keyTable_0_6_port);
   keyTable_reg_0_5_inst : DFFPOSX1 port map( D => n848, CLK => CLK, Q => 
                           keyTable_0_5_port);
   keyTable_reg_0_4_inst : DFFPOSX1 port map( D => n849, CLK => CLK, Q => 
                           keyTable_0_4_port);
   keyTable_reg_0_3_inst : DFFPOSX1 port map( D => n850, CLK => CLK, Q => 
                           keyTable_0_3_port);
   keyTable_reg_0_2_inst : DFFPOSX1 port map( D => n851, CLK => CLK, Q => 
                           keyTable_0_2_port);
   keyTable_reg_0_1_inst : DFFPOSX1 port map( D => n852, CLK => CLK, Q => 
                           keyTable_0_1_port);
   keyTable_reg_0_0_inst : DFFPOSX1 port map( D => n853, CLK => CLK, Q => 
                           keyTable_0_0_port);
   keyTable_reg_1_7_inst : DFFPOSX1 port map( D => n854, CLK => CLK, Q => 
                           keyTable_1_7_port);
   keyTable_reg_0_7_inst : DFFPOSX1 port map( D => n855, CLK => CLK, Q => 
                           keyTable_0_7_port);
   prefillCounter_reg_7_inst : DFFPOSX1 port map( D => n914, CLK => CLK, Q => 
                           prefillCounter_7_port);
   prefillCounter_reg_1_inst : DFFPOSX1 port map( D => n913, CLK => CLK, Q => 
                           prefillCounter_1_port);
   prefillCounter_reg_2_inst : DFFPOSX1 port map( D => n912, CLK => CLK, Q => 
                           prefillCounter_2_port);
   prefillCounter_reg_3_inst : DFFPOSX1 port map( D => n911, CLK => CLK, Q => 
                           prefillCounter_3_port);
   prefillCounter_reg_4_inst : DFFPOSX1 port map( D => n910, CLK => CLK, Q => 
                           prefillCounter_4_port);
   prefillCounter_reg_5_inst : DFFPOSX1 port map( D => n909, CLK => CLK, Q => 
                           prefillCounter_5_port);
   prefillCounter_reg_6_inst : DFFPOSX1 port map( D => n908, CLK => CLK, Q => 
                           prefillCounter_6_port);
   temp_reg_7_inst : DFFPOSX1 port map( D => n856, CLK => CLK, Q => temp_7_port
                           );
   temp_reg_0_inst : DFFPOSX1 port map( D => n863, CLK => CLK, Q => temp_0_port
                           );
   temp_reg_1_inst : DFFPOSX1 port map( D => n862, CLK => CLK, Q => temp_1_port
                           );
   temp_reg_2_inst : DFFPOSX1 port map( D => n861, CLK => CLK, Q => temp_2_port
                           );
   temp_reg_3_inst : DFFPOSX1 port map( D => n860, CLK => CLK, Q => temp_3_port
                           );
   temp_reg_4_inst : DFFPOSX1 port map( D => n859, CLK => CLK, Q => temp_4_port
                           );
   temp_reg_5_inst : DFFPOSX1 port map( D => n858, CLK => CLK, Q => temp_5_port
                           );
   temp_reg_6_inst : DFFPOSX1 port map( D => n857, CLK => CLK, Q => temp_6_port
                           );
   delaydata_reg_7_inst : DFFPOSX1 port map( D => n371, CLK => CLK, Q => 
                           delaydata_7_port);
   delaydata_reg_0_inst : DFFPOSX1 port map( D => n399, CLK => CLK, Q => 
                           delaydata_0_port);
   delaydata_reg_1_inst : DFFPOSX1 port map( D => n395, CLK => CLK, Q => 
                           delaydata_1_port);
   delaydata_reg_2_inst : DFFPOSX1 port map( D => n391, CLK => CLK, Q => 
                           delaydata_2_port);
   delaydata_reg_3_inst : DFFPOSX1 port map( D => n387, CLK => CLK, Q => 
                           delaydata_3_port);
   delaydata_reg_4_inst : DFFPOSX1 port map( D => n383, CLK => CLK, Q => 
                           delaydata_4_port);
   delaydata_reg_5_inst : DFFPOSX1 port map( D => n379, CLK => CLK, Q => 
                           delaydata_5_port);
   delaydata_reg_6_inst : DFFPOSX1 port map( D => n375, CLK => CLK, Q => 
                           delaydata_6_port);
   intj_reg_7_inst : DFFPOSX1 port map( D => n875, CLK => CLK, Q => intj_7_port
                           );
   intj_reg_0_inst : DFFPOSX1 port map( D => n882, CLK => CLK, Q => intj_0_port
                           );
   intj_reg_1_inst : DFFPOSX1 port map( D => n881, CLK => CLK, Q => intj_1_port
                           );
   intj_reg_2_inst : DFFPOSX1 port map( D => n880, CLK => CLK, Q => intj_2_port
                           );
   intj_reg_3_inst : DFFPOSX1 port map( D => n879, CLK => CLK, Q => intj_3_port
                           );
   intj_reg_4_inst : DFFPOSX1 port map( D => n878, CLK => CLK, Q => intj_4_port
                           );
   intj_reg_5_inst : DFFPOSX1 port map( D => n877, CLK => CLK, Q => intj_5_port
                           );
   intj_reg_6_inst : DFFPOSX1 port map( D => n876, CLK => CLK, Q => intj_6_port
                           );
   keyi_reg_2_inst : DFFPOSX1 port map( D => n874, CLK => CLK, Q => keyi_2_port
                           );
   keyi_reg_1_inst : DFFPOSX1 port map( D => n873, CLK => CLK, Q => keyi_1_port
                           );
   keyi_reg_0_inst : DFFPOSX1 port map( D => n872, CLK => CLK, Q => keyi_0_port
                           );
   inti_reg_7_inst : DFFPOSX1 port map( D => n425_port, CLK => CLK, Q => 
                           inti_7_port);
   inti_reg_0_inst : DFFPOSX1 port map( D => n411_port, CLK => CLK, Q => 
                           inti_0_port);
   inti_reg_1_inst : DFFPOSX1 port map( D => n413_port, CLK => CLK, Q => 
                           inti_1_port);
   inti_reg_2_inst : DFFPOSX1 port map( D => n415, CLK => CLK, Q => inti_2_port
                           );
   inti_reg_3_inst : DFFPOSX1 port map( D => n417, CLK => CLK, Q => inti_3_port
                           );
   inti_reg_4_inst : DFFPOSX1 port map( D => n419, CLK => CLK, Q => inti_4_port
                           );
   inti_reg_5_inst : DFFPOSX1 port map( D => n421, CLK => CLK, Q => inti_5_port
                           );
   inti_reg_6_inst : DFFPOSX1 port map( D => n423, CLK => CLK, Q => inti_6_port
                           );
   PROCESSED_DATA_reg_0_inst : DFFPOSX1 port map( D => n759, CLK => CLK, Q => 
                           PROCESSED_DATA_0_port);
   PROCESSED_DATA_reg_1_inst : DFFPOSX1 port map( D => n757, CLK => CLK, Q => 
                           PROCESSED_DATA_1_port);
   PROCESSED_DATA_reg_2_inst : DFFPOSX1 port map( D => n755, CLK => CLK, Q => 
                           PROCESSED_DATA_2_port);
   PROCESSED_DATA_reg_3_inst : DFFPOSX1 port map( D => n753, CLK => CLK, Q => 
                           PROCESSED_DATA_3_port);
   PROCESSED_DATA_reg_4_inst : DFFPOSX1 port map( D => n751, CLK => CLK, Q => 
                           PROCESSED_DATA_4_port);
   PROCESSED_DATA_reg_5_inst : DFFPOSX1 port map( D => n749, CLK => CLK, Q => 
                           PROCESSED_DATA_5_port);
   PROCESSED_DATA_reg_6_inst : DFFPOSX1 port map( D => n747, CLK => CLK, Q => 
                           PROCESSED_DATA_6_port);
   PROCESSED_DATA_reg_7_inst : DFFPOSX1 port map( D => n745, CLK => CLK, Q => 
                           PROCESSED_DATA_7_port);
   faddr_reg_7_inst : DFFPOSX1 port map( D => n744, CLK => CLK, Q => 
                           faddr_7_port);
   ADDR_reg_7_inst : DFFPOSX1 port map( D => n743, CLK => CLK, Q => ADDR_7_port
                           );
   faddr_reg_6_inst : DFFPOSX1 port map( D => n742, CLK => CLK, Q => 
                           faddr_6_port);
   ADDR_reg_6_inst : DFFPOSX1 port map( D => n741, CLK => CLK, Q => ADDR_6_port
                           );
   faddr_reg_5_inst : DFFPOSX1 port map( D => n740, CLK => CLK, Q => 
                           faddr_5_port);
   ADDR_reg_5_inst : DFFPOSX1 port map( D => n739, CLK => CLK, Q => ADDR_5_port
                           );
   faddr_reg_4_inst : DFFPOSX1 port map( D => n738, CLK => CLK, Q => 
                           faddr_4_port);
   ADDR_reg_4_inst : DFFPOSX1 port map( D => n737, CLK => CLK, Q => ADDR_4_port
                           );
   faddr_reg_3_inst : DFFPOSX1 port map( D => n736, CLK => CLK, Q => 
                           faddr_3_port);
   ADDR_reg_3_inst : DFFPOSX1 port map( D => n735, CLK => CLK, Q => ADDR_3_port
                           );
   faddr_reg_2_inst : DFFPOSX1 port map( D => n734, CLK => CLK, Q => 
                           faddr_2_port);
   ADDR_reg_2_inst : DFFPOSX1 port map( D => n733, CLK => CLK, Q => ADDR_2_port
                           );
   faddr_reg_1_inst : DFFPOSX1 port map( D => n732, CLK => CLK, Q => 
                           faddr_1_port);
   ADDR_reg_1_inst : DFFPOSX1 port map( D => n731, CLK => CLK, Q => ADDR_1_port
                           );
   faddr_reg_0_inst : DFFPOSX1 port map( D => n730, CLK => CLK, Q => 
                           faddr_0_port);
   ADDR_reg_0_inst : DFFPOSX1 port map( D => n729, CLK => CLK, Q => ADDR_0_port
                           );
   fdata_reg_7_inst : DFFPOSX1 port map( D => n728, CLK => CLK, Q => 
                           fdata_7_port);
   fdata_reg_6_inst : DFFPOSX1 port map( D => n727, CLK => CLK, Q => 
                           fdata_6_port);
   fdata_reg_5_inst : DFFPOSX1 port map( D => n726, CLK => CLK, Q => 
                           fdata_5_port);
   fdata_reg_4_inst : DFFPOSX1 port map( D => n725, CLK => CLK, Q => 
                           fdata_4_port);
   fdata_reg_3_inst : DFFPOSX1 port map( D => n724, CLK => CLK, Q => 
                           fdata_3_port);
   fdata_reg_2_inst : DFFPOSX1 port map( D => n723, CLK => CLK, Q => 
                           fdata_2_port);
   fdata_reg_1_inst : DFFPOSX1 port map( D => n722, CLK => CLK, Q => 
                           fdata_1_port);
   fdata_reg_0_inst : DFFPOSX1 port map( D => n721, CLK => CLK, Q => 
                           fdata_0_port);
   fw_enable_reg : DFFPOSX1 port map( D => n720, CLK => CLK, Q => fw_enable);
   fr_enable_reg : DFFPOSX1 port map( D => n719, CLK => CLK, Q => fr_enable);
   W_ENABLE_reg : DFFPOSX1 port map( D => n718, CLK => CLK, Q => W_ENABLE_port)
                           ;
   R_ENABLE_reg : DFFPOSX1 port map( D => n717, CLK => CLK, Q => R_ENABLE_port)
                           ;
   DATA_reg_7_inst : DFFPOSX1 port map( D => n716, CLK => CLK, Q => DATA_7_port
                           );
   DATA_reg_6_inst : DFFPOSX1 port map( D => n715, CLK => CLK, Q => DATA_6_port
                           );
   DATA_reg_5_inst : DFFPOSX1 port map( D => n714, CLK => CLK, Q => DATA_5_port
                           );
   DATA_reg_4_inst : DFFPOSX1 port map( D => n713, CLK => CLK, Q => DATA_4_port
                           );
   DATA_reg_3_inst : DFFPOSX1 port map( D => n712, CLK => CLK, Q => DATA_3_port
                           );
   DATA_reg_2_inst : DFFPOSX1 port map( D => n711, CLK => CLK, Q => DATA_2_port
                           );
   DATA_reg_1_inst : DFFPOSX1 port map( D => n710, CLK => CLK, Q => DATA_1_port
                           );
   DATA_reg_0_inst : DFFPOSX1 port map( D => n709, CLK => CLK, Q => DATA_0_port
                           );
   U3 : NOR2X1 port map( A => n11, B => n553, Y => n691);
   U7 : AOI22X1 port map( A => n246, B => extratemp_7_port, C => n572, D => 
                           temp_7_port, Y => n13);
   U8 : OAI21X1 port map( A => n451_port, B => n968, C => n18, Y => n11);
   U9 : AOI22X1 port map( A => DATA_IN(7), B => n244, C => 
                           prefillCounter_7_port, D => n247, Y => n18);
   U10 : NOR2X1 port map( A => n21, B => n551, Y => n693);
   U12 : AOI22X1 port map( A => n246, B => extratemp_6_port, C => n572, D => 
                           temp_6_port, Y => n23);
   U13 : OAI21X1 port map( A => n451_port, B => n969, C => n25, Y => n21);
   U14 : AOI22X1 port map( A => DATA_IN(6), B => n244, C => 
                           prefillCounter_6_port, D => n247, Y => n25);
   U15 : NOR2X1 port map( A => n26, B => n549, Y => n694);
   U17 : AOI22X1 port map( A => n246, B => extratemp_5_port, C => n572, D => 
                           temp_5_port, Y => n28);
   U18 : OAI21X1 port map( A => n451_port, B => n970, C => n30, Y => n26);
   U19 : AOI22X1 port map( A => DATA_IN(5), B => n244, C => 
                           prefillCounter_5_port, D => n247, Y => n30);
   U20 : NOR2X1 port map( A => n31, B => n547, Y => n695);
   U22 : AOI22X1 port map( A => n246, B => extratemp_4_port, C => n572, D => 
                           temp_4_port, Y => n33);
   U23 : OAI21X1 port map( A => n451_port, B => n971, C => n35, Y => n31);
   U24 : AOI22X1 port map( A => DATA_IN(4), B => n244, C => 
                           prefillCounter_4_port, D => n247, Y => n35);
   U25 : NOR2X1 port map( A => n36, B => n545, Y => n696);
   U27 : AOI22X1 port map( A => n246, B => extratemp_3_port, C => n572, D => 
                           temp_3_port, Y => n38);
   U28 : OAI21X1 port map( A => n451_port, B => n972, C => n40, Y => n36);
   U29 : AOI22X1 port map( A => DATA_IN(3), B => n244, C => 
                           prefillCounter_3_port, D => n247, Y => n40);
   U30 : NOR2X1 port map( A => n41, B => n543, Y => n697);
   U32 : AOI22X1 port map( A => n246, B => extratemp_2_port, C => n572, D => 
                           temp_2_port, Y => n43);
   U33 : OAI21X1 port map( A => n451_port, B => n973, C => n45, Y => n41);
   U34 : AOI22X1 port map( A => DATA_IN(2), B => n244, C => 
                           prefillCounter_2_port, D => n247, Y => n45);
   U35 : NOR2X1 port map( A => n46, B => n542, Y => n698);
   U37 : AOI22X1 port map( A => n246, B => extratemp_1_port, C => n572, D => 
                           temp_1_port, Y => n48);
   U38 : OAI21X1 port map( A => n451_port, B => n974, C => n50, Y => n46);
   U39 : AOI22X1 port map( A => DATA_IN(1), B => n244, C => 
                           prefillCounter_1_port, D => n247, Y => n50);
   U40 : NOR2X1 port map( A => n51, B => n541, Y => n699);
   U42 : AOI22X1 port map( A => n246, B => extratemp_0_port, C => n572, D => 
                           temp_0_port, Y => n53);
   U43 : OAI21X1 port map( A => n451_port, B => n975, C => n55, Y => n51);
   U44 : AOI22X1 port map( A => DATA_IN(0), B => n244, C => 
                           prefillCounter_0_port, D => n247, Y => n55);
   U46 : NOR2X1 port map( A => n57, B => n58, Y => n700);
   U47 : NAND2X1 port map( A => n59, B => n60, Y => n58);
   U48 : AOI22X1 port map( A => sj_7_port, B => n61, C => N448, D => n252, Y =>
                           n60);
   U49 : AOI22X1 port map( A => intj_7_port, B => n250, C => N503, D => n241, Y
                           => n59);
   U50 : NAND2X1 port map( A => n65, B => n66, Y => n57);
   U51 : AOI22X1 port map( A => temp_7_port, B => n240, C => inti_7_port, D => 
                           n68, Y => n66);
   U52 : AOI22X1 port map( A => prefillCounter_7_port, B => n247, C => 
                           faddr_7_port, D => n261, Y => n65);
   U53 : NOR2X1 port map( A => n70, B => n71, Y => n702);
   U54 : NAND2X1 port map( A => n72, B => n73, Y => n71);
   U55 : AOI22X1 port map( A => sj_6_port, B => n61, C => N447, D => n252, Y =>
                           n73);
   U56 : AOI22X1 port map( A => intj_6_port, B => n250, C => N502, D => n241, Y
                           => n72);
   U57 : NAND2X1 port map( A => n74, B => n75, Y => n70);
   U58 : AOI22X1 port map( A => temp_6_port, B => n240, C => inti_6_port, D => 
                           n68, Y => n75);
   U59 : AOI22X1 port map( A => prefillCounter_6_port, B => n247, C => 
                           faddr_6_port, D => n261, Y => n74);
   U60 : NOR2X1 port map( A => n76, B => n77, Y => n703);
   U61 : NAND2X1 port map( A => n78, B => n79, Y => n77);
   U62 : AOI22X1 port map( A => sj_5_port, B => n61, C => N446, D => n252, Y =>
                           n79);
   U63 : AOI22X1 port map( A => intj_5_port, B => n250, C => N501, D => n241, Y
                           => n78);
   U64 : NAND2X1 port map( A => n80, B => n81, Y => n76);
   U65 : AOI22X1 port map( A => temp_5_port, B => n240, C => inti_5_port, D => 
                           n68, Y => n81);
   U66 : AOI22X1 port map( A => prefillCounter_5_port, B => n247, C => 
                           faddr_5_port, D => n261, Y => n80);
   U67 : NOR2X1 port map( A => n82, B => n83, Y => n704);
   U68 : NAND2X1 port map( A => n84, B => n85, Y => n83);
   U69 : AOI22X1 port map( A => sj_4_port, B => n61, C => N445, D => n252, Y =>
                           n85);
   U70 : AOI22X1 port map( A => intj_4_port, B => n250, C => N500, D => n241, Y
                           => n84);
   U71 : NAND2X1 port map( A => n86, B => n87, Y => n82);
   U72 : AOI22X1 port map( A => temp_4_port, B => n240, C => inti_4_port, D => 
                           n68, Y => n87);
   U73 : AOI22X1 port map( A => prefillCounter_4_port, B => n247, C => 
                           faddr_4_port, D => n261, Y => n86);
   U74 : NOR2X1 port map( A => n88, B => n89, Y => n705);
   U75 : NAND2X1 port map( A => n90, B => n91, Y => n89);
   U76 : AOI22X1 port map( A => sj_3_port, B => n61, C => N444, D => n252, Y =>
                           n91);
   U77 : AOI22X1 port map( A => intj_3_port, B => n250, C => N499, D => n241, Y
                           => n90);
   U78 : NAND2X1 port map( A => n92, B => n93, Y => n88);
   U79 : AOI22X1 port map( A => temp_3_port, B => n240, C => inti_3_port, D => 
                           n68, Y => n93);
   U80 : AOI22X1 port map( A => prefillCounter_3_port, B => n247, C => 
                           faddr_3_port, D => n261, Y => n92);
   U81 : NOR2X1 port map( A => n94, B => n95, Y => n706);
   U82 : NAND2X1 port map( A => n96, B => n97, Y => n95);
   U83 : AOI22X1 port map( A => sj_2_port, B => n61, C => N443, D => n252, Y =>
                           n97);
   U84 : AOI22X1 port map( A => intj_2_port, B => n250, C => N498, D => n241, Y
                           => n96);
   U85 : NAND2X1 port map( A => n98, B => n99, Y => n94);
   U86 : AOI22X1 port map( A => temp_2_port, B => n240, C => inti_2_port, D => 
                           n68, Y => n99);
   U87 : AOI22X1 port map( A => prefillCounter_2_port, B => n247, C => 
                           faddr_2_port, D => n261, Y => n98);
   U88 : NOR2X1 port map( A => n100, B => n101, Y => n707);
   U89 : NAND2X1 port map( A => n102, B => n103, Y => n101);
   U90 : AOI22X1 port map( A => sj_1_port, B => n61, C => N442, D => n252, Y =>
                           n103);
   U91 : AOI22X1 port map( A => intj_1_port, B => n250, C => N497, D => n241, Y
                           => n102);
   U92 : NAND2X1 port map( A => n104, B => n105, Y => n100);
   U93 : AOI22X1 port map( A => temp_1_port, B => n240, C => inti_1_port, D => 
                           n68, Y => n105);
   U94 : AOI22X1 port map( A => prefillCounter_1_port, B => n247, C => 
                           faddr_1_port, D => n261, Y => n104);
   U95 : NOR2X1 port map( A => n106, B => n107, Y => n708);
   U96 : NAND2X1 port map( A => n108, B => n109, Y => n107);
   U97 : AOI22X1 port map( A => sj_0_port, B => n61, C => n924, D => n252, Y =>
                           n109);
   U98 : OAI21X1 port map( A => n110, B => n111, C => n112, Y => n61);
   U99 : AOI22X1 port map( A => intj_0_port, B => n250, C => N496, D => n241, Y
                           => n108);
   U100 : NAND2X1 port map( A => n113, B => n114, Y => n106);
   U101 : AOI22X1 port map( A => temp_0_port, B => n240, C => inti_0_port, D =>
                           n68, Y => n114);
   U102 : OAI21X1 port map( A => n115, B => n116, C => n503_port, Y => n68);
   U104 : AOI22X1 port map( A => prefillCounter_0_port, B => n247, C => 
                           faddr_0_port, D => n261, Y => n113);
   U106 : OAI21X1 port map( A => n218, B => n188, C => n249, Y => n120);
   U108 : OAI21X1 port map( A => n123, B => n124, C => n125, Y => n119);
   U109 : AOI21X1 port map( A => n126, B => n127, C => n540, Y => n125);
   U110 : NOR2X1 port map( A => KEY_ERROR, B => n128, Y => n126);
   U111 : OAI21X1 port map( A => n361, B => n130, C => n359, Y => n124);
   U112 : NAND3X1 port map( A => n132, B => n133, C => n134, Y => 
                           nextState_3_port);
   U113 : AOI21X1 port map( A => n571, B => n606, C => n137, Y => n134);
   U114 : NAND2X1 port map( A => n138, B => n139, Y => n137);
   U115 : AOI22X1 port map( A => n140, B => n359, C => n522_port, D => n142, Y 
                           => n132);
   U116 : NAND3X1 port map( A => n143, B => n144, C => n145, Y => 
                           nextState_2_port);
   U117 : NOR2X1 port map( A => n146, B => n147, Y => n145);
   U118 : OAI21X1 port map( A => n148, B => n110, C => n133, Y => n147);
   U119 : AOI21X1 port map( A => n149, B => permuteComplete, C => n150, Y => 
                           n133);
   U120 : NAND2X1 port map( A => n507, B => n152, Y => n150);
   U121 : OAI22X1 port map( A => n116, B => n153, C => KEY_ERROR, D => n154, Y 
                           => n146);
   U122 : AOI22X1 port map( A => n155, B => n156, C => n157, D => n158, Y => 
                           n154);
   U123 : NOR2X1 port map( A => n159, B => n361, Y => n155);
   U124 : NOR2X1 port map( A => n246, B => n600, Y => n144);
   U125 : NOR2X1 port map( A => n594, B => n162, Y => n143);
   U126 : NAND3X1 port map( A => n163, B => n164, C => n165, Y => 
                           nextState_1_port);
   U127 : NOR2X1 port map( A => n166, B => n167, Y => n165);
   U128 : OAI21X1 port map( A => n168, B => n169, C => n170, Y => n167);
   U129 : NAND3X1 port map( A => n171, B => n401, C => n173, Y => n169);
   U130 : NOR2X1 port map( A => prefillCounter_2_port, B => 
                           prefillCounter_1_port, Y => n173);
   U131 : NAND3X1 port map( A => n174, B => n889, C => n176, Y => n168);
   U132 : NOR2X1 port map( A => prefillCounter_4_port, B => 
                           prefillCounter_3_port, Y => n176);
   U133 : NOR2X1 port map( A => prefillCounter_7_port, B => 
                           prefillCounter_6_port, Y => n174);
   U135 : AOI22X1 port map( A => n178, B => state_0_port, C => n179, D => n359,
                           Y => n163);
   U137 : OAI21X1 port map( A => n518_port, B => n158, C => n181, Y => n179);
   U138 : NAND2X1 port map( A => n142, B => n182, Y => n181);
   U139 : OAI21X1 port map( A => n183, B => n158, C => n184, Y => n182);
   U140 : OAI21X1 port map( A => n159, B => n361, C => n569, Y => n184);
   U143 : NAND3X1 port map( A => n367, B => n365, C => BYTE_READY, Y => n158);
   U145 : NOR2X1 port map( A => state_1_port, B => n116, Y => n178);
   U146 : NAND3X1 port map( A => n189, B => n190, C => n191, Y => 
                           nextState_0_port);
   U147 : NOR2X1 port map( A => n252, B => n192, Y => n191);
   U148 : OAI21X1 port map( A => KEY_ERROR, B => n193, C => n164, Y => n192);
   U149 : NOR2X1 port map( A => n194, B => n195, Y => n164);
   U150 : OAI21X1 port map( A => permuteComplete, B => n562, C => n197, Y => 
                           n195);
   U151 : NAND3X1 port map( A => n152, B => n198, C => n199, Y => n194);
   U152 : AOI21X1 port map( A => n156, B => n128, C => n200, Y => n193);
   U153 : OAI21X1 port map( A => n218, B => n201, C => n202, Y => n200);
   U154 : NAND3X1 port map( A => BYTE_READY, B => n157, C => n363, Y => n202);
   U156 : NAND2X1 port map( A => OPCODE(0), B => n365, Y => n130);
   U158 : NAND2X1 port map( A => BYTE_READY, B => n204, Y => n128);
   U159 : OAI21X1 port map( A => OPCODE(0), B => OPCODE(1), C => n186, Y => 
                           n204);
   U160 : NAND2X1 port map( A => OPCODE(1), B => OPCODE(0), Y => n186);
   U161 : NOR2X1 port map( A => n540, B => n246, Y => n190);
   U162 : NOR2X1 port map( A => n171, B => n205, Y => n189);
   U163 : OAI21X1 port map( A => n300, B => n403, C => n207, Y => n709);
   U164 : NAND2X1 port map( A => DATA_0_port, B => n290, Y => n207);
   U165 : OAI21X1 port map( A => n302, B => n449_port, C => n209, Y => n710);
   U166 : NAND2X1 port map( A => DATA_1_port, B => n305, Y => n209);
   U167 : OAI21X1 port map( A => n302, B => n447_port, C => n211, Y => n711);
   U168 : NAND2X1 port map( A => DATA_2_port, B => n305, Y => n211);
   U169 : OAI21X1 port map( A => n302, B => n445_port, C => n213, Y => n712);
   U170 : NAND2X1 port map( A => DATA_3_port, B => n305, Y => n213);
   U171 : OAI21X1 port map( A => n302, B => n443_port, C => n215, Y => n713);
   U172 : NAND2X1 port map( A => DATA_4_port, B => RST, Y => n215);
   U173 : OAI21X1 port map( A => n302, B => n441, C => n217, Y => n714);
   U174 : NAND2X1 port map( A => DATA_5_port, B => n305, Y => n217);
   U175 : OAI21X1 port map( A => n302, B => n439, C => n219, Y => n715);
   U176 : NAND2X1 port map( A => DATA_6_port, B => n305, Y => n219);
   U177 : OAI21X1 port map( A => n302, B => n437, C => n221, Y => n716);
   U178 : NAND2X1 port map( A => DATA_7_port, B => n305, Y => n221);
   U179 : OAI21X1 port map( A => n302, B => n222, C => n223, Y => n717);
   U180 : NAND2X1 port map( A => R_ENABLE_port, B => n305, Y => n223);
   U181 : AOI21X1 port map( A => fr_enable, B => n224, C => n225, Y => n222);
   U182 : OAI21X1 port map( A => n300, B => n226, C => n227, Y => n718);
   U183 : NAND2X1 port map( A => W_ENABLE_port, B => n302, Y => n227);
   U184 : AOI21X1 port map( A => fw_enable, B => n185, C => n229, Y => n226);
   U185 : OAI21X1 port map( A => n300, B => n504, C => n231, Y => n719);
   U186 : OAI21X1 port map( A => n300, B => n224, C => fr_enable, Y => n231);
   U187 : NAND3X1 port map( A => n3, B => n233, C => n234, Y => n224);
   U188 : NOR2X1 port map( A => n577, B => n236, Y => n234);
   U189 : NAND2X1 port map( A => n210, B => n10, Y => n236);
   U191 : NAND2X1 port map( A => n579, B => n604, Y => n112);
   U192 : OAI21X1 port map( A => n300, B => n514_port, C => n242, Y => n720);
   U193 : OAI21X1 port map( A => n300, B => n185, C => fw_enable, Y => n242);
   U195 : NAND3X1 port map( A => n210, B => n10, C => n243, Y => n229);
   U196 : NOR2X1 port map( A => n244, B => n572, Y => n243);
   U197 : OAI22X1 port map( A => n331, B => n975, C => n297, D => n403, Y => 
                           n721);
   U200 : OAI22X1 port map( A => n331, B => n974, C => n295, D => n449_port, Y 
                           => n722);
   U203 : OAI22X1 port map( A => n331, B => n973, C => n297, D => n447_port, Y 
                           => n723);
   U206 : OAI22X1 port map( A => n331, B => n972, C => n295, D => n445_port, Y 
                           => n724);
   U209 : OAI22X1 port map( A => n333, B => n971, C => n297, D => n443_port, Y 
                           => n725);
   U212 : OAI22X1 port map( A => n329, B => n970, C => n295, D => n441, Y => 
                           n726);
   U215 : OAI22X1 port map( A => n329, B => n969, C => n297, D => n439, Y => 
                           n727);
   U218 : OAI22X1 port map( A => n329, B => n968, C => n295, D => n437, Y => 
                           n728);
   U221 : OAI21X1 port map( A => n300, B => n405, C => n245, Y => n729);
   U222 : NAND2X1 port map( A => ADDR_0_port, B => n302, Y => n245);
   U223 : OAI22X1 port map( A => n326, B => n967, C => n295, D => n405, Y => 
                           n730);
   U226 : OAI21X1 port map( A => n300, B => n471, C => n248, Y => n731);
   U227 : NAND2X1 port map( A => ADDR_1_port, B => n305, Y => n248);
   U228 : OAI22X1 port map( A => n335, B => n966, C => n295, D => n471, Y => 
                           n732);
   U231 : OAI21X1 port map( A => n300, B => n473_port, C => n251, Y => n733);
   U232 : NAND2X1 port map( A => ADDR_2_port, B => n302, Y => n251);
   U233 : OAI22X1 port map( A => n337, B => n965, C => n295, D => n473_port, Y 
                           => n734);
   U236 : OAI21X1 port map( A => n300, B => n475_port, C => n254, Y => n735);
   U237 : NAND2X1 port map( A => ADDR_3_port, B => n305, Y => n254);
   U238 : OAI22X1 port map( A => n327, B => n964, C => n295, D => n475_port, Y 
                           => n736);
   U241 : OAI21X1 port map( A => n300, B => n480_port, C => n257, Y => n737);
   U242 : NAND2X1 port map( A => ADDR_4_port, B => n305, Y => n257);
   U243 : OAI22X1 port map( A => n307, B => n963, C => n295, D => n480_port, Y 
                           => n738);
   U246 : OAI21X1 port map( A => n300, B => n482_port, C => n260, Y => n739);
   U247 : NAND2X1 port map( A => ADDR_5_port, B => n305, Y => n260);
   U248 : OAI22X1 port map( A => n318, B => n962, C => n295, D => n482_port, Y 
                           => n740);
   U251 : OAI21X1 port map( A => n297, B => n488, C => n263, Y => n741);
   U252 : NAND2X1 port map( A => ADDR_6_port, B => n305, Y => n263);
   U253 : OAI22X1 port map( A => n317, B => n961, C => n295, D => n488, Y => 
                           n742);
   U256 : OAI21X1 port map( A => n297, B => n498_port, C => n266, Y => n743);
   U257 : NAND2X1 port map( A => ADDR_7_port, B => n305, Y => n266);
   U258 : OAI22X1 port map( A => n311, B => n960, C => n295, D => n498_port, Y 
                           => n744);
   U261 : OAI21X1 port map( A => n297, B => n369, C => n269, Y => n745);
   U262 : NAND2X1 port map( A => PROCESSED_DATA_7_port, B => n305, Y => n269);
   U264 : OAI21X1 port map( A => n500_port, B => n959, C => n272, Y => 
                           nextProcessedData_7_port);
   U265 : AOI22X1 port map( A => n273, B => n274, C => BYTE(7), D => n575, Y =>
                           n272);
   U266 : XOR2X1 port map( A => temp_7_port, B => delaydata_7_port, Y => n274);
   U268 : OAI21X1 port map( A => n297, B => n373, C => n276, Y => n747);
   U269 : NAND2X1 port map( A => PROCESSED_DATA_6_port, B => n305, Y => n276);
   U271 : OAI21X1 port map( A => n500_port, B => n958, C => n278, Y => 
                           nextProcessedData_6_port);
   U272 : AOI22X1 port map( A => n273, B => n279, C => BYTE(6), D => n575, Y =>
                           n278);
   U273 : XOR2X1 port map( A => temp_6_port, B => delaydata_6_port, Y => n279);
   U275 : OAI21X1 port map( A => n297, B => n377, C => n281, Y => n749);
   U276 : NAND2X1 port map( A => PROCESSED_DATA_5_port, B => n305, Y => n281);
   U278 : OAI21X1 port map( A => n500_port, B => n957, C => n283, Y => 
                           nextProcessedData_5_port);
   U279 : AOI22X1 port map( A => n273, B => n284, C => BYTE(5), D => n575, Y =>
                           n283);
   U280 : XOR2X1 port map( A => temp_5_port, B => delaydata_5_port, Y => n284);
   U282 : OAI21X1 port map( A => n297, B => n381, C => n286, Y => n751);
   U283 : NAND2X1 port map( A => PROCESSED_DATA_4_port, B => n305, Y => n286);
   U285 : OAI21X1 port map( A => n500_port, B => n956, C => n288, Y => 
                           nextProcessedData_4_port);
   U286 : AOI22X1 port map( A => n273, B => n289, C => BYTE(4), D => n575, Y =>
                           n288);
   U287 : XOR2X1 port map( A => temp_4_port, B => delaydata_4_port, Y => n289);
   U289 : OAI21X1 port map( A => n300, B => n385, C => n291, Y => n753);
   U290 : NAND2X1 port map( A => PROCESSED_DATA_3_port, B => n305, Y => n291);
   U292 : OAI21X1 port map( A => n500_port, B => n955, C => n293, Y => 
                           nextProcessedData_3_port);
   U293 : AOI22X1 port map( A => n273, B => n294, C => BYTE(3), D => n575, Y =>
                           n293);
   U294 : XOR2X1 port map( A => temp_3_port, B => delaydata_3_port, Y => n294);
   U296 : OAI21X1 port map( A => n297, B => n389, C => n296, Y => n755);
   U297 : NAND2X1 port map( A => PROCESSED_DATA_2_port, B => n305, Y => n296);
   U299 : OAI21X1 port map( A => n500_port, B => n954, C => n298, Y => 
                           nextProcessedData_2_port);
   U300 : AOI22X1 port map( A => n273, B => n299, C => BYTE(2), D => n575, Y =>
                           n298);
   U301 : XOR2X1 port map( A => temp_2_port, B => delaydata_2_port, Y => n299);
   U303 : OAI21X1 port map( A => n297, B => n393, C => n301, Y => n757);
   U304 : NAND2X1 port map( A => PROCESSED_DATA_1_port, B => RST, Y => n301);
   U306 : OAI21X1 port map( A => n500_port, B => n953, C => n303, Y => 
                           nextProcessedData_1_port);
   U307 : AOI22X1 port map( A => n273, B => n304, C => BYTE(1), D => n575, Y =>
                           n303);
   U308 : XOR2X1 port map( A => temp_1_port, B => delaydata_1_port, Y => n304);
   U310 : OAI21X1 port map( A => n297, B => n397, C => n306, Y => n759);
   U311 : NAND2X1 port map( A => PROCESSED_DATA_0_port, B => RST, Y => n306);
   U313 : OAI21X1 port map( A => n500_port, B => n952, C => n308, Y => 
                           nextProcessedData_0_port);
   U314 : AOI22X1 port map( A => n273, B => n309, C => BYTE(0), D => n575, Y =>
                           n308);
   U315 : XOR2X1 port map( A => temp_0_port, B => delaydata_0_port, Y => n309);
   U318 : NAND3X1 port map( A => n253, B => n505, C => n312, Y => n310);
   U319 : NOR2X1 port map( A => n313, B => n314, Y => n312);
   U322 : AOI22X1 port map( A => BYTE(7), B => n6, C => n262, D => 
                           delaydata_7_port, Y => n316);
   U324 : AOI22X1 port map( A => BYTE(0), B => n6, C => n262, D => 
                           delaydata_0_port, Y => n319);
   U326 : AOI22X1 port map( A => BYTE(1), B => n6, C => n262, D => 
                           delaydata_1_port, Y => n320);
   U328 : AOI22X1 port map( A => BYTE(2), B => n6, C => n262, D => 
                           delaydata_2_port, Y => n321);
   U330 : AOI22X1 port map( A => BYTE(3), B => n6, C => n262, D => 
                           delaydata_3_port, Y => n322);
   U332 : AOI22X1 port map( A => BYTE(4), B => n6, C => n262, D => 
                           delaydata_4_port, Y => n323);
   U334 : AOI22X1 port map( A => BYTE(5), B => n6, C => n262, D => 
                           delaydata_5_port, Y => n324);
   U336 : AOI22X1 port map( A => BYTE(6), B => n6, C => n262, D => 
                           delaydata_6_port, Y => n325);
   U339 : OAI21X1 port map( A => n271, B => n616, C => n330, Y => n792);
   U340 : NAND2X1 port map( A => KEY(56), B => n287, Y => n330);
   U342 : OAI21X1 port map( A => n268, B => n618, C => n332, Y => n793);
   U343 : NAND2X1 port map( A => KEY(57), B => n287, Y => n332);
   U345 : OAI21X1 port map( A => n268, B => n624, C => n334, Y => n794);
   U346 : NAND2X1 port map( A => KEY(58), B => n287, Y => n334);
   U348 : OAI21X1 port map( A => n268, B => n626, C => n336, Y => n795);
   U349 : NAND2X1 port map( A => KEY(59), B => n287, Y => n336);
   U351 : OAI21X1 port map( A => n268, B => n629, C => n338, Y => n796);
   U352 : NAND2X1 port map( A => KEY(60), B => n287, Y => n338);
   U354 : OAI21X1 port map( A => n268, B => n630, C => n340, Y => n797);
   U355 : NAND2X1 port map( A => KEY(61), B => n285, Y => n340);
   U357 : OAI21X1 port map( A => n268, B => n632, C => n342, Y => n798);
   U358 : NAND2X1 port map( A => KEY(62), B => n285, Y => n342);
   U360 : OAI21X1 port map( A => n268, B => n636, C => n344, Y => n799);
   U361 : NAND2X1 port map( A => KEY(63), B => n285, Y => n344);
   U363 : OAI21X1 port map( A => n268, B => n637, C => n346, Y => n800);
   U364 : NAND2X1 port map( A => KEY(48), B => n285, Y => n346);
   U366 : OAI21X1 port map( A => n268, B => n638, C => n348, Y => n801);
   U367 : NAND2X1 port map( A => KEY(49), B => n285, Y => n348);
   U369 : OAI21X1 port map( A => n268, B => n648, C => n350, Y => n802);
   U370 : NAND2X1 port map( A => KEY(50), B => n285, Y => n350);
   U372 : OAI21X1 port map( A => n268, B => n649, C => n352, Y => n803);
   U373 : NAND2X1 port map( A => KEY(51), B => n285, Y => n352);
   U375 : OAI21X1 port map( A => n268, B => n650, C => n354, Y => n804);
   U376 : NAND2X1 port map( A => KEY(52), B => n285, Y => n354);
   U378 : OAI21X1 port map( A => n268, B => n651, C => n356, Y => n805);
   U379 : NAND2X1 port map( A => KEY(53), B => n285, Y => n356);
   U381 : OAI21X1 port map( A => n270, B => n692, C => n358, Y => n806);
   U382 : NAND2X1 port map( A => KEY(54), B => n285, Y => n358);
   U384 : OAI21X1 port map( A => n270, B => n701, C => n360, Y => n807);
   U385 : NAND2X1 port map( A => KEY(55), B => n282, Y => n360);
   U387 : OAI21X1 port map( A => n270, B => n746, C => n362, Y => n808);
   U388 : NAND2X1 port map( A => KEY(40), B => n285, Y => n362);
   U390 : OAI21X1 port map( A => n270, B => n748, C => n364, Y => n809);
   U391 : NAND2X1 port map( A => KEY(41), B => n285, Y => n364);
   U393 : OAI21X1 port map( A => n270, B => n750, C => n366, Y => n810);
   U394 : NAND2X1 port map( A => KEY(42), B => n282, Y => n366);
   U396 : OAI21X1 port map( A => n270, B => n752, C => n368, Y => n811);
   U397 : NAND2X1 port map( A => KEY(43), B => n285, Y => n368);
   U399 : OAI21X1 port map( A => n270, B => n754, C => n370, Y => n812);
   U400 : NAND2X1 port map( A => KEY(44), B => n282, Y => n370);
   U402 : OAI21X1 port map( A => n270, B => n756, C => n372, Y => n813);
   U403 : NAND2X1 port map( A => KEY(45), B => n282, Y => n372);
   U405 : OAI21X1 port map( A => n270, B => n758, C => n374, Y => n814);
   U406 : NAND2X1 port map( A => KEY(46), B => n282, Y => n374);
   U408 : OAI21X1 port map( A => n270, B => n760, C => n376, Y => n815);
   U409 : NAND2X1 port map( A => KEY(47), B => n282, Y => n376);
   U411 : OAI21X1 port map( A => n270, B => n761, C => n378, Y => n816);
   U412 : NAND2X1 port map( A => KEY(32), B => n282, Y => n378);
   U414 : OAI21X1 port map( A => n270, B => n762, C => n380, Y => n817);
   U415 : NAND2X1 port map( A => KEY(33), B => n282, Y => n380);
   U417 : OAI21X1 port map( A => n270, B => n763, C => n382, Y => n818);
   U418 : NAND2X1 port map( A => KEY(34), B => n280, Y => n382);
   U420 : OAI21X1 port map( A => n271, B => n764, C => n384, Y => n819);
   U421 : NAND2X1 port map( A => KEY(35), B => n280, Y => n384);
   U423 : OAI21X1 port map( A => n271, B => n765, C => n386, Y => n820);
   U424 : NAND2X1 port map( A => KEY(36), B => n282, Y => n386);
   U426 : OAI21X1 port map( A => n271, B => n766, C => n388, Y => n821);
   U427 : NAND2X1 port map( A => KEY(37), B => n280, Y => n388);
   U429 : OAI21X1 port map( A => n271, B => n767, C => n390, Y => n822);
   U430 : NAND2X1 port map( A => KEY(38), B => n280, Y => n390);
   U432 : OAI21X1 port map( A => n271, B => n768, C => n392, Y => n823);
   U433 : NAND2X1 port map( A => KEY(39), B => n282, Y => n392);
   U435 : OAI21X1 port map( A => n275, B => n769, C => n394, Y => n824);
   U436 : NAND2X1 port map( A => KEY(24), B => n280, Y => n394);
   U437 : OAI21X1 port map( A => n271, B => n770, C => n396, Y => n825);
   U438 : NAND2X1 port map( A => KEY(25), B => n280, Y => n396);
   U439 : OAI21X1 port map( A => n271, B => n771, C => n398, Y => n826);
   U440 : NAND2X1 port map( A => KEY(26), B => n280, Y => n398);
   U441 : OAI21X1 port map( A => n271, B => n772, C => n400, Y => n827);
   U442 : NAND2X1 port map( A => KEY(27), B => n280, Y => n400);
   U443 : OAI21X1 port map( A => n271, B => n773, C => n402, Y => n828);
   U444 : NAND2X1 port map( A => KEY(28), B => n280, Y => n402);
   U445 : OAI21X1 port map( A => n271, B => n774, C => n404, Y => n829);
   U446 : NAND2X1 port map( A => KEY(29), B => n280, Y => n404);
   U447 : OAI21X1 port map( A => n271, B => n775, C => n406, Y => n830);
   U448 : NAND2X1 port map( A => KEY(30), B => n280, Y => n406);
   U449 : OAI21X1 port map( A => n271, B => n776, C => n408_port, Y => n831);
   U450 : NAND2X1 port map( A => KEY(31), B => n280, Y => n408_port);
   U451 : OAI21X1 port map( A => n275, B => n777, C => n410_port, Y => n832);
   U452 : NAND2X1 port map( A => KEY(16), B => n280, Y => n410_port);
   U453 : OAI21X1 port map( A => n275, B => n778, C => n412_port, Y => n833);
   U454 : NAND2X1 port map( A => KEY(17), B => n277, Y => n412_port);
   U455 : OAI21X1 port map( A => n275, B => n779, C => n414_port, Y => n834);
   U456 : NAND2X1 port map( A => KEY(18), B => n280, Y => n414_port);
   U457 : OAI21X1 port map( A => n275, B => n780, C => n416, Y => n835);
   U458 : NAND2X1 port map( A => KEY(19), B => n280, Y => n416);
   U459 : OAI21X1 port map( A => n275, B => n781, C => n418, Y => n836);
   U460 : NAND2X1 port map( A => KEY(20), B => n282, Y => n418);
   U461 : OAI21X1 port map( A => n275, B => n782, C => n420, Y => n837);
   U462 : NAND2X1 port map( A => KEY(21), B => n280, Y => n420);
   U463 : OAI21X1 port map( A => n275, B => n783, C => n422, Y => n838);
   U464 : NAND2X1 port map( A => KEY(22), B => n282, Y => n422);
   U465 : OAI21X1 port map( A => n275, B => n784, C => n424_port, Y => n839);
   U466 : NAND2X1 port map( A => KEY(23), B => n280, Y => n424_port);
   U467 : OAI21X1 port map( A => n277, B => n785, C => n426_port, Y => n840);
   U468 : NAND2X1 port map( A => KEY(8), B => n282, Y => n426_port);
   U469 : OAI21X1 port map( A => n277, B => n786, C => n428_port, Y => n841);
   U470 : NAND2X1 port map( A => KEY(9), B => n282, Y => n428_port);
   U471 : OAI21X1 port map( A => n275, B => n787, C => n430_port, Y => n842);
   U472 : NAND2X1 port map( A => KEY(10), B => n280, Y => n430_port);
   U473 : OAI21X1 port map( A => n277, B => n788, C => n432, Y => n843);
   U474 : NAND2X1 port map( A => KEY(11), B => n282, Y => n432);
   U475 : OAI21X1 port map( A => n277, B => n789, C => n434, Y => n844);
   U476 : NAND2X1 port map( A => KEY(12), B => n282, Y => n434);
   U477 : OAI21X1 port map( A => n275, B => n790, C => n436, Y => n845);
   U478 : NAND2X1 port map( A => KEY(13), B => n282, Y => n436);
   U479 : OAI21X1 port map( A => n275, B => n791, C => n438, Y => n846);
   U480 : NAND2X1 port map( A => KEY(14), B => n285, Y => n438);
   U481 : OAI21X1 port map( A => n277, B => n864, C => n440, Y => n847);
   U482 : NAND2X1 port map( A => KEY(6), B => n282, Y => n440);
   U483 : OAI21X1 port map( A => n275, B => n865, C => n442_port, Y => n848);
   U484 : NAND2X1 port map( A => KEY(5), B => n285, Y => n442_port);
   U485 : OAI21X1 port map( A => n277, B => n866, C => n444_port, Y => n849);
   U486 : NAND2X1 port map( A => KEY(4), B => n285, Y => n444_port);
   U487 : OAI21X1 port map( A => n277, B => n867, C => n446_port, Y => n850);
   U488 : NAND2X1 port map( A => KEY(3), B => n285, Y => n446_port);
   U489 : OAI21X1 port map( A => n277, B => n868, C => n448_port, Y => n851);
   U490 : NAND2X1 port map( A => KEY(2), B => n285, Y => n448_port);
   U491 : OAI21X1 port map( A => n277, B => n869, C => n450, Y => n852);
   U492 : NAND2X1 port map( A => KEY(1), B => n287, Y => n450);
   U493 : OAI21X1 port map( A => n277, B => n870, C => n452, Y => n853);
   U494 : NAND2X1 port map( A => KEY(0), B => n287, Y => n452);
   U495 : OAI21X1 port map( A => n277, B => n871, C => n454, Y => n854);
   U496 : NAND2X1 port map( A => KEY(15), B => n287, Y => n454);
   U497 : OAI21X1 port map( A => n277, B => n883, C => n456, Y => n855);
   U498 : NAND2X1 port map( A => KEY(7), B => n287, Y => n456);
   U499 : NOR2X1 port map( A => n457, B => n313, Y => n328);
   U500 : OAI21X1 port map( A => n469, B => n916, C => n460, Y => n856);
   U501 : AOI22X1 port map( A => N527, B => n14, C => n180, D => DATA_IN(7), Y 
                           => n460);
   U503 : OAI21X1 port map( A => n469, B => n923, C => n464, Y => n857);
   U504 : AOI22X1 port map( A => N526, B => n14, C => n180, D => DATA_IN(6), Y 
                           => n464);
   U506 : OAI21X1 port map( A => n469, B => n922, C => n466, Y => n858);
   U507 : AOI22X1 port map( A => N525, B => n14, C => n180, D => DATA_IN(5), Y 
                           => n466);
   U509 : OAI21X1 port map( A => n469, B => n921, C => n468, Y => n859);
   U510 : AOI22X1 port map( A => N524, B => n14, C => n180, D => DATA_IN(4), Y 
                           => n468);
   U512 : OAI21X1 port map( A => n469, B => n920, C => n470, Y => n860);
   U513 : AOI22X1 port map( A => N523, B => n14, C => n180, D => DATA_IN(3), Y 
                           => n470);
   U515 : OAI21X1 port map( A => n469, B => n919, C => n472_port, Y => n861);
   U516 : AOI22X1 port map( A => N522, B => n14, C => n180, D => DATA_IN(2), Y 
                           => n472_port);
   U518 : OAI21X1 port map( A => n469, B => n918, C => n474_port, Y => n862);
   U519 : AOI22X1 port map( A => N521, B => n14, C => n180, D => DATA_IN(1), Y 
                           => n474_port);
   U521 : OAI21X1 port map( A => n469, B => n917, C => n476_port, Y => n863);
   U522 : AOI22X1 port map( A => N520, B => n14, C => n180, D => DATA_IN(0), Y 
                           => n476_port);
   U527 : NAND3X1 port map( A => n479_port, B => n509, C => n481_port, Y => 
                           n477_port);
   U528 : NOR2X1 port map( A => n315, B => n261, Y => n481_port);
   U530 : NAND3X1 port map( A => n483_port, B => n210, C => n484_port, Y => 
                           n315);
   U532 : NOR2X1 port map( A => n302, B => n171, Y => n479_port);
   U534 : AOI22X1 port map( A => n259, B => extratemp_0_port, C => DATA_IN(0), 
                           D => n258, Y => n486_port);
   U536 : AOI22X1 port map( A => n259, B => extratemp_1_port, C => DATA_IN(1), 
                           D => n258, Y => n489);
   U538 : AOI22X1 port map( A => n259, B => extratemp_2_port, C => DATA_IN(2), 
                           D => n258, Y => n490);
   U540 : AOI22X1 port map( A => n259, B => extratemp_3_port, C => DATA_IN(3), 
                           D => n258, Y => n491);
   U542 : AOI22X1 port map( A => n259, B => extratemp_4_port, C => DATA_IN(4), 
                           D => n258, Y => n492);
   U544 : AOI22X1 port map( A => n259, B => extratemp_5_port, C => DATA_IN(5), 
                           D => n258, Y => n493);
   U546 : AOI22X1 port map( A => n259, B => extratemp_6_port, C => DATA_IN(6), 
                           D => n258, Y => n494);
   U548 : AOI22X1 port map( A => n259, B => extratemp_7_port, C => DATA_IN(7), 
                           D => n258, Y => n495);
   U550 : NAND3X1 port map( A => n138, B => n210, C => n496_port, Y => 
                           n487_port);
   U551 : NOR2X1 port map( A => n497_port, B => n56, Y => n496_port);
   U552 : NAND3X1 port map( A => n5, B => n520_port, C => n3, Y => n56);
   U553 : NAND2X1 port map( A => n579, B => n142, Y => n138);
   U555 : OAI22X1 port map( A => n429_port, B => n924, C => n502_port, D => 
                           n951, Y => n872);
   U556 : OAI22X1 port map( A => n429_port, B => n357, C => n502_port, D => 
                           n228, Y => n873);
   U557 : OAI22X1 port map( A => n429_port, B => n925, C => n502_port, D => 
                           n945, Y => n874);
   U559 : NOR2X1 port map( A => n508, B => n313, Y => n502_port);
   U560 : OAI21X1 port map( A => n409_port, B => n930, C => n510, Y => n875);
   U561 : NAND2X1 port map( A => N519, B => n511, Y => n510);
   U563 : OAI21X1 port map( A => n409_port, B => n937, C => n513_port, Y => 
                           n876);
   U564 : NAND2X1 port map( A => N518, B => n511, Y => n513_port);
   U566 : OAI21X1 port map( A => n409_port, B => n936, C => n515_port, Y => 
                           n877);
   U567 : NAND2X1 port map( A => N517, B => n511, Y => n515_port);
   U569 : OAI21X1 port map( A => n409_port, B => n935, C => n517_port, Y => 
                           n878);
   U570 : NAND2X1 port map( A => N516, B => n511, Y => n517_port);
   U572 : OAI21X1 port map( A => n409_port, B => n934, C => n519_port, Y => 
                           n879);
   U573 : NAND2X1 port map( A => N515, B => n511, Y => n519_port);
   U575 : OAI21X1 port map( A => n409_port, B => n933, C => n521_port, Y => 
                           n880);
   U576 : NAND2X1 port map( A => N514, B => n511, Y => n521_port);
   U578 : OAI21X1 port map( A => n409_port, B => n932, C => n523_port, Y => 
                           n881);
   U579 : NAND2X1 port map( A => N513, B => n511, Y => n523_port);
   U581 : OAI21X1 port map( A => n409_port, B => n931, C => n525_port, Y => 
                           n882);
   U582 : NAND2X1 port map( A => N512, B => n511, Y => n525_port);
   U583 : NOR2X1 port map( A => n152, B => n526_port, Y => n511);
   U587 : NOR2X1 port map( A => n302, B => n594, Y => n529);
   U589 : AOI22X1 port map( A => n256, B => inti_7_port, C => N503, D => n216, 
                           Y => n530);
   U591 : AOI22X1 port map( A => n256, B => inti_6_port, C => N502, D => n216, 
                           Y => n533);
   U593 : AOI22X1 port map( A => n256, B => inti_5_port, C => N501, D => n216, 
                           Y => n534);
   U595 : AOI22X1 port map( A => n256, B => inti_4_port, C => N500, D => n216, 
                           Y => n535);
   U597 : AOI22X1 port map( A => n256, B => inti_3_port, C => N499, D => n214, 
                           Y => n536);
   U599 : AOI22X1 port map( A => n256, B => inti_2_port, C => N498, D => n214, 
                           Y => n537);
   U601 : AOI22X1 port map( A => n256, B => inti_1_port, C => N497, D => n214, 
                           Y => n538);
   U603 : AOI22X1 port map( A => n256, B => inti_0_port, C => N496, D => n214, 
                           Y => n539);
   U604 : NOR2X1 port map( A => n256, B => n507, Y => n532);
   U605 : NAND3X1 port map( A => n557, B => n520_port, C => n431_port, Y => 
                           n531);
   U606 : OAI21X1 port map( A => n407_port, B => n220, C => n544, Y => n891);
   U607 : NAND2X1 port map( A => N480, B => n594, Y => n544);
   U609 : OAI21X1 port map( A => n407_port, B => n944, C => n546, Y => n892);
   U610 : NAND2X1 port map( A => N481, B => n594, Y => n546);
   U612 : OAI21X1 port map( A => n407_port, B => n943, C => n548, Y => n893);
   U613 : NAND2X1 port map( A => N482, B => n594, Y => n548);
   U615 : OAI21X1 port map( A => n407_port, B => n942, C => n550, Y => n894);
   U616 : NAND2X1 port map( A => N483, B => n594, Y => n550);
   U618 : OAI21X1 port map( A => n407_port, B => n941, C => n552, Y => n895);
   U619 : NAND2X1 port map( A => N484, B => n594, Y => n552);
   U621 : OAI21X1 port map( A => n407_port, B => n940, C => n554, Y => n896);
   U622 : NAND2X1 port map( A => N485, B => n594, Y => n554);
   U624 : OAI21X1 port map( A => n407_port, B => n939, C => n556, Y => n897);
   U625 : NAND2X1 port map( A => N486, B => n594, Y => n556);
   U628 : NAND2X1 port map( A => N487, B => n594, Y => n558);
   U631 : NAND3X1 port map( A => n528, B => n152, C => n527_port, Y => n559);
   U632 : NOR2X1 port map( A => n560, B => n561, Y => n527_port);
   U633 : NAND3X1 port map( A => n3, B => n557, C => n435, Y => n561);
   U634 : NAND3X1 port map( A => n581, B => n520_port, C => n563, Y => n560);
   U637 : OAI21X1 port map( A => n557, B => n565, C => n566, Y => n899);
   U638 : OAI21X1 port map( A => n567, B => n508, C => permuteComplete, Y => 
                           n566);
   U639 : NAND2X1 port map( A => n568, B => n427_port, Y => n565);
   U641 : NAND3X1 port map( A => n172, B => n507, C => n431_port, Y => n508);
   U643 : NAND3X1 port map( A => n253, B => n329, C => n435, Y => n570);
   U646 : OAI21X1 port map( A => n433, B => n929, C => n573, Y => n900);
   U647 : NAND2X1 port map( A => N431, B => n574, Y => n573);
   U649 : OAI21X1 port map( A => n433, B => n928, C => n576, Y => n901);
   U650 : NAND2X1 port map( A => N430, B => n574, Y => n576);
   U652 : OAI21X1 port map( A => n433, B => n927, C => n578, Y => n902);
   U653 : NAND2X1 port map( A => N429, B => n574, Y => n578);
   U654 : OAI21X1 port map( A => n433, B => n926, C => n580, Y => n903);
   U655 : NAND2X1 port map( A => N428, B => n574, Y => n580);
   U656 : OAI21X1 port map( A => n433, B => n355, C => n582, Y => n904);
   U657 : NAND2X1 port map( A => N427, B => n574, Y => n582);
   U659 : OAI21X1 port map( A => n433, B => n925, C => n583, Y => n905);
   U660 : NAND2X1 port map( A => N426, B => n574, Y => n583);
   U662 : OAI21X1 port map( A => n433, B => n357, C => n584, Y => n906);
   U663 : NAND2X1 port map( A => N425, B => n574, Y => n584);
   U664 : OAI21X1 port map( A => n433, B => n924, C => n585, Y => n907);
   U665 : NAND2X1 port map( A => N424, B => n574, Y => n585);
   U666 : NOR2X1 port map( A => n557, B => n568, Y => n574);
   U667 : NOR2X1 port map( A => n586, B => n587, Y => n568);
   U668 : NAND3X1 port map( A => si_7_port, B => si_6_port, C => n588, Y => 
                           n587);
   U669 : NOR2X1 port map( A => n926, B => n927, Y => n588);
   U672 : NAND3X1 port map( A => si_3_port, B => si_2_port, C => n589, Y => 
                           n586);
   U673 : NOR2X1 port map( A => n924, B => n357, Y => n589);
   U677 : NAND3X1 port map( A => n435, B => n253, C => n591, Y => n590);
   U678 : NOR2X1 port map( A => n241, B => n313, Y => n591);
   U679 : NOR2X1 port map( A => n203, B => n116, Y => n313);
   U681 : OAI21X1 port map( A => n218, B => n499_port, C => n524_port, Y => 
                           n593);
   U684 : NAND3X1 port map( A => n123, B => n484_port, C => n597, Y => n596);
   U685 : NOR2X1 port map( A => n598, B => n599, Y => n597);
   U686 : OAI21X1 port map( A => n218, B => n170, C => n139, Y => n599);
   U690 : OAI21X1 port map( A => n111, B => n602, C => n10, Y => n63);
   U693 : OAI21X1 port map( A => n467, B => n890, C => n607, Y => n908);
   U694 : NAND2X1 port map( A => N413, B => n608, Y => n607);
   U696 : OAI21X1 port map( A => n467, B => n889, C => n609, Y => n909);
   U697 : NAND2X1 port map( A => N412, B => n608, Y => n609);
   U699 : OAI21X1 port map( A => n467, B => n888, C => n611, Y => n910);
   U700 : NAND2X1 port map( A => N411, B => n608, Y => n611);
   U702 : OAI21X1 port map( A => n467, B => n887, C => n613, Y => n911);
   U703 : NAND2X1 port map( A => N410, B => n608, Y => n613);
   U705 : OAI21X1 port map( A => n467, B => n886, C => n615, Y => n912);
   U706 : NAND2X1 port map( A => N409, B => n608, Y => n615);
   U708 : OAI21X1 port map( A => n467, B => n885, C => n617, Y => n913);
   U709 : NAND2X1 port map( A => N408, B => n608, Y => n617);
   U711 : OAI21X1 port map( A => n467, B => n884, C => n619, Y => n914);
   U712 : NAND2X1 port map( A => N414, B => n608, Y => n619);
   U714 : OAI21X1 port map( A => n467, B => n401, C => n620, Y => n915);
   U715 : NAND2X1 port map( A => N407, B => n608, Y => n620);
   U716 : NOR2X1 port map( A => n457, B => n210, Y => n608);
   U721 : NAND3X1 port map( A => n5, B => n197, C => n621, Y => n457);
   U722 : NOR2X1 port map( A => n506, B => n497_port, Y => n621);
   U723 : NAND3X1 port map( A => n8, B => n581, C => n622, Y => n497_port);
   U724 : NOR2X1 port map( A => n302, B => n246, Y => n622);
   U727 : NOR2X1 port map( A => n116, B => n499_port, Y => n171);
   U731 : NOR2X1 port map( A => n485_port, B => n162, Y => n232);
   U732 : NOR2X1 port map( A => n183, B => n110, Y => n162);
   U733 : OAI21X1 port map( A => n116, B => n625, C => n512_port, Y => 
                           n485_port);
   U735 : OAI21X1 port map( A => n170, B => n605, C => n562, Y => n627);
   U737 : NOR2X1 port map( A => n111, B => n605, Y => n149);
   U738 : NAND3X1 port map( A => n628, B => n604, C => n592, Y => n197);
   U739 : XOR2X1 port map( A => n4, B => n218, Y => n628);
   U743 : NAND2X1 port map( A => n483_port, B => n516_port, Y => n225);
   U745 : OAI21X1 port map( A => n111, B => n602, C => n601, Y => n631);
   U746 : NAND2X1 port map( A => n606, B => n177, Y => n601);
   U748 : NOR2X1 port map( A => n598, B => n241, Y => n483_port);
   U750 : OAI21X1 port map( A => n110, B => n111, C => n633, Y => n598);
   U751 : NOR2X1 port map( A => n600, B => n118, Y => n633);
   U752 : NOR2X1 port map( A => n183, B => n116, Y => n118);
   U754 : NAND2X1 port map( A => n67, B => n4, Y => n198);
   U755 : NOR2X1 port map( A => n314, B => n540, Y => n233);
   U757 : NOR2X1 port map( A => n273, B => n575, Y => n139);
   U759 : NAND3X1 port map( A => n142, B => n592, C => n4, Y => n634);
   U760 : NOR2X1 port map( A => n623, B => n605, Y => n273);
   U762 : OAI21X1 port map( A => n170, B => n110, C => n557, Y => n635);
   U764 : NOR2X1 port map( A => n111, B => n116, Y => n567);
   U765 : NAND2X1 port map( A => n571, B => n610, Y => n111);
   U766 : NAND2X1 port map( A => state_0_port, B => n522_port, Y => n170);
   U767 : NAND2X1 port map( A => n518_port, B => n501_port, Y => n140);
   U769 : AOI21X1 port map( A => n183, B => n625, C => n605, Y => n156);
   U771 : NOR2X1 port map( A => n614, B => state_2_port, Y => n142);
   U772 : NAND3X1 port map( A => n4, B => n555, C => state_0_port, Y => n183);
   U774 : NAND2X1 port map( A => n172, B => n603, Y => n157);
   U780 : NAND2X1 port map( A => n555, B => n161, Y => n148);
   U781 : NOR2X1 port map( A => n595, B => n594, Y => n478_port);
   U783 : NAND2X1 port map( A => n240, B => n188, Y => n199);
   U784 : NOR2X1 port map( A => n110, B => n115, Y => n67);
   U785 : NAND3X1 port map( A => n152, B => n564, C => n528, Y => n595);
   U787 : NOR2X1 port map( A => n116, B => n623, Y => n205);
   U788 : NAND3X1 port map( A => n612, B => n555, C => n4, Y => n623);
   U790 : NAND2X1 port map( A => n604, B => n614, Y => n116);
   U792 : NAND2X1 port map( A => n569, B => n606, Y => n564);
   U794 : NAND2X1 port map( A => state_2_port, B => n614, Y => n110);
   U797 : NAND2X1 port map( A => n571, B => n4, Y => n625);
   U799 : NAND2X1 port map( A => state_0_port, B => state_1_port, Y => n153);
   U801 : NAND2X1 port map( A => n592, B => n188, Y => n499_port);
   U804 : NAND2X1 port map( A => state_1_port, B => n612, Y => n115);
   U806 : NAND2X1 port map( A => state_2_port, B => n218, Y => n602);
   U807 : NAND3X1 port map( A => n639, B => n641, C => n640, Y => N479);
   U808 : NOR2X1 port map( A => n643, B => n642, Y => n641);
   U809 : OAI22X1 port map( A => n785, B => n212, C => n870, D => n645, Y => 
                           n643);
   U812 : OAI22X1 port map( A => n769, B => n646, C => n777, D => n647, Y => 
                           n642);
   U815 : AOI22X1 port map( A => n947, B => keyTable_5_0_port, C => n946, D => 
                           keyTable_4_0_port, Y => n640);
   U816 : AOI22X1 port map( A => n949, B => keyTable_7_0_port, C => 
                           keyTable_6_0_port, D => n948, Y => n639);
   U817 : NAND3X1 port map( A => n652, B => n653, C => n654, Y => N478);
   U818 : NOR2X1 port map( A => n655, B => n656, Y => n654);
   U819 : OAI22X1 port map( A => n786, B => n212, C => n869, D => n645, Y => 
                           n656);
   U822 : OAI22X1 port map( A => n770, B => n646, C => n778, D => n647, Y => 
                           n655);
   U825 : AOI22X1 port map( A => n947, B => keyTable_5_1_port, C => n946, D => 
                           keyTable_4_1_port, Y => n653);
   U826 : AOI22X1 port map( A => n949, B => keyTable_7_1_port, C => n948, D => 
                           keyTable_6_1_port, Y => n652);
   U827 : NAND3X1 port map( A => n657, B => n658, C => n659, Y => N477);
   U828 : NOR2X1 port map( A => n660, B => n661, Y => n659);
   U829 : OAI22X1 port map( A => n787, B => n212, C => n868, D => n645, Y => 
                           n661);
   U832 : OAI22X1 port map( A => n771, B => n646, C => n779, D => n647, Y => 
                           n660);
   U835 : AOI22X1 port map( A => n947, B => keyTable_5_2_port, C => n946, D => 
                           keyTable_4_2_port, Y => n658);
   U836 : AOI22X1 port map( A => n949, B => keyTable_7_2_port, C => n948, D => 
                           keyTable_6_2_port, Y => n657);
   U837 : NAND3X1 port map( A => n662, B => n663, C => n664, Y => N476);
   U838 : NOR2X1 port map( A => n665, B => n666, Y => n664);
   U839 : OAI22X1 port map( A => n788, B => n212, C => n867, D => n645, Y => 
                           n666);
   U842 : OAI22X1 port map( A => n772, B => n646, C => n780, D => n647, Y => 
                           n665);
   U845 : AOI22X1 port map( A => n947, B => keyTable_5_3_port, C => n946, D => 
                           keyTable_4_3_port, Y => n663);
   U846 : AOI22X1 port map( A => n949, B => keyTable_7_3_port, C => n948, D => 
                           keyTable_6_3_port, Y => n662);
   U847 : NAND3X1 port map( A => n667, B => n668, C => n669, Y => N475);
   U848 : NOR2X1 port map( A => n670, B => n671, Y => n669);
   U849 : OAI22X1 port map( A => n789, B => n212, C => n866, D => n645, Y => 
                           n671);
   U852 : OAI22X1 port map( A => n773, B => n646, C => n781, D => n647, Y => 
                           n670);
   U855 : AOI22X1 port map( A => n947, B => keyTable_5_4_port, C => n946, D => 
                           keyTable_4_4_port, Y => n668);
   U856 : AOI22X1 port map( A => n949, B => keyTable_7_4_port, C => n948, D => 
                           keyTable_6_4_port, Y => n667);
   U857 : NAND3X1 port map( A => n672, B => n673, C => n674, Y => N474);
   U858 : NOR2X1 port map( A => n675, B => n676, Y => n674);
   U859 : OAI22X1 port map( A => n790, B => n212, C => n865, D => n645, Y => 
                           n676);
   U862 : OAI22X1 port map( A => n774, B => n646, C => n782, D => n647, Y => 
                           n675);
   U865 : AOI22X1 port map( A => n947, B => keyTable_5_5_port, C => n946, D => 
                           keyTable_4_5_port, Y => n673);
   U866 : AOI22X1 port map( A => n949, B => keyTable_7_5_port, C => n948, D => 
                           keyTable_6_5_port, Y => n672);
   U867 : NAND3X1 port map( A => n677, B => n678, C => n679, Y => N473);
   U868 : NOR2X1 port map( A => n680, B => n681, Y => n679);
   U869 : OAI22X1 port map( A => n791, B => n212, C => n864, D => n645, Y => 
                           n681);
   U872 : OAI22X1 port map( A => n775, B => n237, C => n783, D => n647, Y => 
                           n680);
   U875 : AOI22X1 port map( A => n947, B => keyTable_5_6_port, C => n946, D => 
                           keyTable_4_6_port, Y => n678);
   U876 : AOI22X1 port map( A => n949, B => keyTable_7_6_port, C => n948, D => 
                           keyTable_6_6_port, Y => n677);
   U877 : NAND3X1 port map( A => n682, B => n683, C => n684, Y => N472);
   U878 : NOR2X1 port map( A => n685, B => n686, Y => n684);
   U879 : OAI22X1 port map( A => n871, B => n212, C => n883, D => n645, Y => 
                           n686);
   U880 : NAND3X1 port map( A => n950, B => n945, C => n951, Y => n645);
   U882 : NAND3X1 port map( A => n950, B => keyi_0_port, C => n945, Y => n644);
   U884 : OAI22X1 port map( A => n776, B => n237, C => n784, D => n647, Y => 
                           n685);
   U885 : NAND3X1 port map( A => n951, B => n945, C => keyi_1_port, Y => n647);
   U887 : NAND3X1 port map( A => keyi_1_port, B => n230, C => n945, Y => n646);
   U890 : AOI22X1 port map( A => n947, B => keyTable_5_7_port, C => n946, D => 
                           keyTable_4_7_port, Y => n683);
   U892 : NAND3X1 port map( A => n951, B => n228, C => n235, Y => n687);
   U894 : NAND3X1 port map( A => n228, B => n230, C => n235, Y => n688);
   U896 : AOI22X1 port map( A => n949, B => keyTable_7_7_port, C => n948, D => 
                           keyTable_6_7_port, Y => n682);
   U898 : NAND3X1 port map( A => n951, B => keyi_1_port, C => n235, Y => n689);
   U901 : NAND3X1 port map( A => keyi_1_port, B => n230, C => n235, Y => n690);
   U105 : OR2X2 port map( A => n119, B => n120, Y => nextState_4_port);
   U134 : OR2X2 port map( A => n162, B => n575, Y => n166);
   U142 : AND2X2 port map( A => n130, B => n186, Y => n159);
   U635 : AND2X2 port map( A => n507, B => n564, Y => n563);
   U692 : AND2X2 port map( A => n603, B => n501_port, Y => n123);
   U761 : OR2X2 port map( A => n140, B => n635, Y => n314);
   U775 : OR2X2 port map( A => n602, B => n623, Y => n603);
   U800 : OR2X2 port map( A => n602, B => n499_port, Y => n152);
   add_377 : KSA_1_DW01_add_0 port map( A(7) => temp_7_port, A(6) => 
                           temp_6_port, A(5) => temp_5_port, A(4) => 
                           temp_4_port, A(3) => temp_3_port, A(2) => 
                           temp_2_port, A(1) => temp_1_port, A(0) => 
                           temp_0_port, B(7) => extratemp_7_port, B(6) => 
                           extratemp_6_port, B(5) => extratemp_5_port, B(4) => 
                           extratemp_4_port, B(3) => extratemp_3_port, B(2) => 
                           extratemp_2_port, B(1) => extratemp_1_port, B(0) => 
                           extratemp_0_port, CI => n1, SUM(7) => N527, SUM(6) 
                           => N526, SUM(5) => N525, SUM(4) => N524, SUM(3) => 
                           N523, SUM(2) => N522, SUM(1) => N521, SUM(0) => N520
                           , CO => n_1026);
   add_337 : KSA_1_DW01_add_1 port map( A(7) => intj_7_port, A(6) => 
                           intj_6_port, A(5) => intj_5_port, A(4) => 
                           intj_4_port, A(3) => intj_3_port, A(2) => 
                           intj_2_port, A(1) => intj_1_port, A(0) => 
                           intj_0_port, B(7) => DATA_IN(7), B(6) => DATA_IN(6),
                           B(5) => DATA_IN(5), B(4) => DATA_IN(4), B(3) => 
                           DATA_IN(3), B(2) => DATA_IN(2), B(1) => DATA_IN(1), 
                           B(0) => DATA_IN(0), CI => n2, SUM(7) => N519, SUM(6)
                           => N518, SUM(5) => N517, SUM(4) => N516, SUM(3) => 
                           N515, SUM(2) => N514, SUM(1) => N513, SUM(0) => N512
                           , CO => n_1027);
   add_289 : KSA_1_DW01_inc_0 port map( A(7) => si_7_port, A(6) => si_6_port, 
                           A(5) => si_5_port, A(4) => si_4_port, A(3) => 
                           si_3_port, A(2) => si_2_port, A(1) => si_1_port, 
                           A(0) => si_0_port, SUM(7) => N431, SUM(6) => N430, 
                           SUM(5) => N429, SUM(4) => N428, SUM(3) => N427, 
                           SUM(2) => N426, SUM(1) => N425, SUM(0) => N424);
   add_263 : KSA_1_DW01_inc_1 port map( A(7) => prefillCounter_7_port, A(6) => 
                           prefillCounter_6_port, A(5) => prefillCounter_5_port
                           , A(4) => prefillCounter_4_port, A(3) => 
                           prefillCounter_3_port, A(2) => prefillCounter_2_port
                           , A(1) => prefillCounter_1_port, A(0) => 
                           prefillCounter_0_port, SUM(7) => N414, SUM(6) => 
                           N413, SUM(5) => N412, SUM(4) => N411, SUM(3) => N410
                           , SUM(2) => N409, SUM(1) => N408, SUM(0) => N407);
   r126 : KSA_1_DW01_inc_2 port map( A(7) => inti_7_port, A(6) => inti_6_port, 
                           A(5) => inti_5_port, A(4) => inti_4_port, A(3) => 
                           inti_3_port, A(2) => inti_2_port, A(1) => 
                           inti_1_port, A(0) => inti_0_port, SUM(7) => N503, 
                           SUM(6) => N502, SUM(5) => N501, SUM(4) => N500, 
                           SUM(3) => N499, SUM(2) => N498, SUM(1) => N497, 
                           SUM(0) => N496);
   add_1_root_add_0_root_add_302_2 : KSA_1_DW01_add_3 port map( A(7) => 
                           DATA_IN(7), A(6) => DATA_IN(6), A(5) => DATA_IN(5), 
                           A(4) => DATA_IN(4), A(3) => DATA_IN(3), A(2) => 
                           DATA_IN(2), A(1) => DATA_IN(1), A(0) => DATA_IN(0), 
                           B(7) => sj_7_port, B(6) => sj_6_port, B(5) => 
                           sj_5_port, B(4) => sj_4_port, B(3) => sj_3_port, 
                           B(2) => sj_2_port, B(1) => sj_1_port, B(0) => 
                           sj_0_port, CI => n976, SUM(7) => N456_port, SUM(6) 
                           => N455, SUM(5) => N454_port, SUM(4) => N453, SUM(3)
                           => N452_port, SUM(2) => N451, SUM(1) => N450_port, 
                           SUM(0) => N449, CO => n_1028);
   add_0_root_add_0_root_add_302_2 : KSA_1_DW01_add_2 port map( A(7) => N472, 
                           A(6) => N473, A(5) => N474, A(4) => N475, A(3) => 
                           N476, A(2) => N477, A(1) => N478, A(0) => N479, B(7)
                           => N456_port, B(6) => N455, B(5) => N454_port, B(4) 
                           => N453, B(3) => N452_port, B(2) => N451, B(1) => 
                           N450_port, B(0) => N449, CI => n977, SUM(7) => N487,
                           SUM(6) => N486, SUM(5) => N485, SUM(4) => N484, 
                           SUM(3) => N483, SUM(2) => N482, SUM(1) => N481, 
                           SUM(0) => N480, CO => n_1029);
   nfaddr_tri_5_inst : TBUFX1 port map( A => n703, EN => n253, Y => 
                           nfaddr_5_port);
   nfaddr_tri_0_inst : TBUFX1 port map( A => n708, EN => n253, Y => 
                           nfaddr_0_port);
   nfaddr_tri_1_inst : TBUFX1 port map( A => n707, EN => n253, Y => 
                           nfaddr_1_port);
   nfaddr_tri_2_inst : TBUFX1 port map( A => n706, EN => n253, Y => 
                           nfaddr_2_port);
   nfaddr_tri_3_inst : TBUFX1 port map( A => n705, EN => n253, Y => 
                           nfaddr_3_port);
   nfaddr_tri_4_inst : TBUFX1 port map( A => n704, EN => n253, Y => 
                           nfaddr_4_port);
   nfaddr_tri_6_inst : TBUFX1 port map( A => n702, EN => n253, Y => 
                           nfaddr_6_port);
   nfaddr_tri_7_inst : TBUFX1 port map( A => n700, EN => n253, Y => 
                           nfaddr_7_port);
   nfdata_tri_0_inst : TBUFX1 port map( A => n699, EN => n581, Y => 
                           nfdata_0_port);
   nfdata_tri_1_inst : TBUFX1 port map( A => n698, EN => n581, Y => 
                           nfdata_1_port);
   nfdata_tri_2_inst : TBUFX1 port map( A => n697, EN => n581, Y => 
                           nfdata_2_port);
   nfdata_tri_3_inst : TBUFX1 port map( A => n696, EN => n581, Y => 
                           nfdata_3_port);
   nfdata_tri_4_inst : TBUFX1 port map( A => n695, EN => n581, Y => 
                           nfdata_4_port);
   nfdata_tri_5_inst : TBUFX1 port map( A => n694, EN => n581, Y => 
                           nfdata_5_port);
   nfdata_tri_6_inst : TBUFX1 port map( A => n693, EN => n581, Y => 
                           nfdata_6_port);
   nfdata_tri_7_inst : TBUFX1 port map( A => n691, EN => n581, Y => 
                           nfdata_7_port);
   PDATA_READY_reg : DFFSR port map( D => n540, CLK => CLK, R => n292, S => 
                           n160, Q => PDATA_READY);
   state_reg_1_inst : DFFSR port map( D => nextState_1_port, CLK => CLK, R => 
                           n292, S => n151, Q => state_1_port);
   state_reg_4_inst : DFFSR port map( D => nextState_4_port, CLK => CLK, R => 
                           n292, S => n141, Q => state_4_port);
   state_reg_3_inst : DFFSR port map( D => nextState_3_port, CLK => CLK, R => 
                           n292, S => n136, Q => state_3_port);
   state_reg_2_inst : DFFSR port map( D => nextState_2_port, CLK => CLK, R => 
                           n292, S => n135, Q => state_2_port);
   state_reg_0_inst : DFFSR port map( D => nextState_0_port, CLK => CLK, R => 
                           n292, S => n131, Q => state_0_port);
   si_reg_7_inst : DFFSR port map( D => n900, CLK => CLK, R => n292, S => n129,
                           Q => si_7_port);
   si_reg_6_inst : DFFSR port map( D => n901, CLK => CLK, R => n292, S => n122,
                           Q => si_6_port);
   si_reg_5_inst : DFFSR port map( D => n902, CLK => CLK, R => n292, S => n121,
                           Q => si_5_port);
   si_reg_4_inst : DFFSR port map( D => n903, CLK => CLK, R => n292, S => n117,
                           Q => si_4_port);
   si_reg_3_inst : DFFSR port map( D => n904, CLK => CLK, R => n292, S => n69, 
                           Q => si_3_port);
   si_reg_2_inst : DFFSR port map( D => n905, CLK => CLK, R => n292, S => n64, 
                           Q => si_2_port);
   si_reg_1_inst : DFFSR port map( D => n906, CLK => CLK, R => n292, S => n62, 
                           Q => si_1_port);
   si_reg_0_inst : DFFSR port map( D => n907, CLK => CLK, R => n292, S => n54, 
                           Q => si_0_port);
   sj_reg_4_inst : DFFSR port map( D => n895, CLK => CLK, R => n292, S => n52, 
                           Q => sj_4_port);
   sj_reg_3_inst : DFFSR port map( D => n894, CLK => CLK, R => n292, S => n49, 
                           Q => sj_3_port);
   sj_reg_2_inst : DFFSR port map( D => n893, CLK => CLK, R => n292, S => n47, 
                           Q => sj_2_port);
   sj_reg_1_inst : DFFSR port map( D => n892, CLK => CLK, R => n292, S => n44, 
                           Q => sj_1_port);
   sj_reg_0_inst : DFFSR port map( D => n891, CLK => CLK, R => n292, S => n42, 
                           Q => sj_0_port);
   sj_reg_5_inst : DFFSR port map( D => n896, CLK => CLK, R => n292, S => n39, 
                           Q => sj_5_port);
   currentProcessedData_reg_7_inst : DFFSR port map( D => 
                           nextProcessedData_7_port, CLK => CLK, R => n292, S 
                           => n37, Q => currentProcessedData_7_port);
   currentProcessedData_reg_6_inst : DFFSR port map( D => 
                           nextProcessedData_6_port, CLK => CLK, R => n292, S 
                           => n34, Q => currentProcessedData_6_port);
   currentProcessedData_reg_5_inst : DFFSR port map( D => 
                           nextProcessedData_5_port, CLK => CLK, R => n292, S 
                           => n32, Q => currentProcessedData_5_port);
   currentProcessedData_reg_4_inst : DFFSR port map( D => 
                           nextProcessedData_4_port, CLK => CLK, R => n292, S 
                           => n29, Q => currentProcessedData_4_port);
   currentProcessedData_reg_3_inst : DFFSR port map( D => 
                           nextProcessedData_3_port, CLK => CLK, R => n292, S 
                           => n27, Q => currentProcessedData_3_port);
   currentProcessedData_reg_2_inst : DFFSR port map( D => 
                           nextProcessedData_2_port, CLK => CLK, R => n292, S 
                           => n24, Q => currentProcessedData_2_port);
   currentProcessedData_reg_1_inst : DFFSR port map( D => 
                           nextProcessedData_1_port, CLK => CLK, R => n292, S 
                           => n22, Q => currentProcessedData_1_port);
   currentProcessedData_reg_0_inst : DFFSR port map( D => 
                           nextProcessedData_0_port, CLK => CLK, R => n292, S 
                           => n20, Q => currentProcessedData_0_port);
   sj_reg_6_inst : DFFSR port map( D => n897, CLK => CLK, R => n292, S => n19, 
                           Q => sj_6_port);
   sj_reg_7_inst : DFFSR port map( D => n898, CLK => CLK, R => n292, S => n17, 
                           Q => sj_7_port);
   U4 : BUFX4 port map( A => n232, Y => n3);
   U11 : OR2X1 port map( A => n602, B => n170, Y => n12);
   U16 : INVX4 port map( A => n7, Y => n261);
   U21 : INVX2 port map( A => n688, Y => n947);
   U26 : INVX2 port map( A => n687, Y => n946);
   U31 : INVX2 port map( A => n602, Y => n175);
   U36 : INVX2 port map( A => n12, Y => n241);
   U41 : INVX2 port map( A => n255, Y => n256);
   U45 : INVX2 port map( A => n477_port, Y => n469);
   U103 : BUFX2 port map( A => state_4_port, Y => n4);
   U107 : AND2X2 port map( A => n233, B => n9, Y => n5);
   U136 : AND2X2 port map( A => n409_port, B => n172, Y => n6);
   U141 : AND2X2 port map( A => n233, B => n520_port, Y => n7);
   U144 : INVX2 port map( A => n10, Y => n246);
   U155 : OR2X2 port map( A => n201, B => n605, Y => n8);
   U157 : AND2X2 port map( A => n504, B => n478_port, Y => n9);
   U190 : OR2X2 port map( A => n110, B => n623, Y => n10);
   U194 : AND2X2 port map( A => n162, B => n469, Y => n14);
   U198 : INVX2 port map( A => n258, Y => n259);
   U199 : INVX2 port map( A => keyi_1_port, Y => n950);
   U201 : INVX2 port map( A => n8, Y => n244);
   U202 : AND2X2 port map( A => n8, B => n601, Y => n15);
   U204 : AND2X2 port map( A => n529, B => n528, Y => n16);
   U205 : INVX2 port map( A => n249, Y => n250);
   U207 : INVX4 port map( A => RST, Y => n292);
   n17 <= '1';
   n19 <= '1';
   n20 <= '1';
   n22 <= '1';
   n24 <= '1';
   n27 <= '1';
   n29 <= '1';
   n32 <= '1';
   n34 <= '1';
   n37 <= '1';
   n39 <= '1';
   n42 <= '1';
   n44 <= '1';
   n47 <= '1';
   n49 <= '1';
   n52 <= '1';
   n54 <= '1';
   n62 <= '1';
   n64 <= '1';
   n69 <= '1';
   n117 <= '1';
   n121 <= '1';
   n122 <= '1';
   n129 <= '1';
   n131 <= '1';
   n135 <= '1';
   n136 <= '1';
   n141 <= '1';
   n151 <= '1';
   n160 <= '1';
   U281 : INVX1 port map( A => n241, Y => n507);
   U284 : BUFX4 port map( A => n644, Y => n212);
   U288 : INVX1 port map( A => n4, Y => n161);
   U291 : INVX1 port map( A => n4, Y => n610);
   U295 : NAND2X1 port map( A => n175, B => n177, Y => n172);
   U298 : INVX1 port map( A => n172, Y => n127);
   U302 : AND2X1 port map( A => n522_port, B => n612, Y => n177);
   U305 : BUFX2 port map( A => n206, Y => n180);
   U309 : INVX2 port map( A => n5, Y => n185);
   U312 : INVX2 port map( A => n196, Y => n484_port);
   U316 : INVX1 port map( A => n610, Y => n187);
   U317 : INVX2 port map( A => n187, Y => n188);
   U320 : NAND3X1 port map( A => n249, B => n197, C => n15, Y => n196);
   U321 : INVX1 port map( A => n15, Y => n252);
   U323 : NAND2X1 port map( A => n527_port, B => n16, Y => n526_port);
   U325 : NAND2X1 port map( A => n522_port, B => n612, Y => n201);
   U327 : NAND2X1 port map( A => n522_port, B => n612, Y => n203);
   U329 : INVX2 port map( A => n142, Y => n605);
   U331 : INVX2 port map( A => n326, Y => n297);
   U333 : INVX2 port map( A => n318, Y => n300);
   U335 : INVX2 port map( A => n311, Y => n305);
   U337 : INVX2 port map( A => n317, Y => n302);
   U338 : INVX2 port map( A => n327, Y => n295);
   U341 : BUFX2 port map( A => n265, Y => n275);
   U344 : BUFX2 port map( A => n264, Y => n270);
   U347 : BUFX2 port map( A => n264, Y => n268);
   U350 : BUFX2 port map( A => n264, Y => n271);
   U353 : BUFX2 port map( A => n265, Y => n277);
   U356 : BUFX2 port map( A => n265, Y => n280);
   U359 : BUFX2 port map( A => n267, Y => n282);
   U362 : BUFX2 port map( A => n267, Y => n285);
   U365 : BUFX2 port map( A => n267, Y => n287);
   U368 : BUFX2 port map( A => n333, Y => n329);
   U371 : BUFX2 port map( A => n335, Y => n327);
   U374 : BUFX2 port map( A => n307, Y => n326);
   U377 : BUFX2 port map( A => n335, Y => n318);
   U380 : BUFX2 port map( A => n307, Y => n317);
   U383 : BUFX2 port map( A => n337, Y => n311);
   U386 : BUFX2 port map( A => n337, Y => n307);
   U389 : BUFX2 port map( A => n333, Y => n331);
   U392 : INVX2 port map( A => n171, Y => n581);
   U395 : INVX4 port map( A => n6, Y => n262);
   U398 : NOR2X1 port map( A => n477_port, B => n478_port, Y => n206);
   U401 : BUFX2 port map( A => n328, Y => n265);
   U404 : BUFX2 port map( A => n328, Y => n267);
   U407 : BUFX2 port map( A => n328, Y => n264);
   U410 : INVX2 port map( A => n290, Y => n335);
   U413 : INVX2 port map( A => n290, Y => n333);
   U416 : INVX2 port map( A => n290, Y => n337);
   U419 : INVX2 port map( A => n199, Y => n594);
   U422 : INVX2 port map( A => n559, Y => n407_port);
   U425 : INVX2 port map( A => n487_port, Y => n258);
   U428 : INVX2 port map( A => n210, Y => n247);
   U431 : INVX2 port map( A => n208, Y => n253);
   U434 : INVX2 port map( A => n292, Y => n290);
   U502 : INVX2 port map( A => n197, Y => n572);
   U505 : INVX2 port map( A => n689, Y => n948);
   U508 : OR2X2 port map( A => n506, B => n593, Y => n208);
   U511 : OR2X2 port map( A => n170, B => n116, Y => n210);
   U514 : INVX2 port map( A => n239, Y => n240);
   U517 : INVX2 port map( A => n63, Y => n249);
   U520 : INVX2 port map( A => n690, Y => n949);
   U523 : INVX2 port map( A => n634, Y => n575);
   U524 : INVX2 port map( A => keyi_2_port, Y => n945);
   U525 : BUFX2 port map( A => keyi_2_port, Y => n235);
   U526 : BUFX2 port map( A => n950, Y => n228);
   U529 : BUFX2 port map( A => n532, Y => n214);
   U531 : BUFX2 port map( A => n532, Y => n216);
   U533 : BUFX2 port map( A => state_3_port, Y => n218);
   U535 : INVX2 port map( A => sj_0_port, Y => n220);
   U537 : INVX2 port map( A => keyi_0_port, Y => n951);
   U539 : BUFX2 port map( A => keyi_0_port, Y => n230);
   U541 : BUFX2 port map( A => n646, Y => n237);
   U543 : INVX2 port map( A => n531, Y => n255);
   U545 : INVX1 port map( A => n457, Y => n467);
   U547 : INVX2 port map( A => n67, Y => n239);
   U549 : OR2X2 port map( A => n407_port, B => n938, Y => n238);
   U554 : NAND2X1 port map( A => n238, B => n558, Y => n898);
   U558 : INVX1 port map( A => n110, Y => n606);
   U562 : INVX4 port map( A => n526_port, Y => n409_port);
   U565 : NAND2X1 port map( A => n357, B => n924, Y => n339);
   U568 : OAI21X1 port map( A => n924, B => n357, C => n339, Y => N442);
   U571 : NOR2X1 port map( A => n339, B => si_2_port, Y => n343);
   U574 : AOI21X1 port map( A => n339, B => si_2_port, C => n343, Y => n341);
   U577 : NAND2X1 port map( A => n343, B => n355, Y => n345);
   U580 : OAI21X1 port map( A => n343, B => n355, C => n345, Y => N444);
   U584 : NOR2X1 port map( A => n345, B => si_4_port, Y => n349);
   U585 : AOI21X1 port map( A => n345, B => si_4_port, C => n349, Y => n347);
   U586 : NAND2X1 port map( A => n349, B => n927, Y => n351);
   U588 : OAI21X1 port map( A => n349, B => n927, C => n351, Y => N446);
   U590 : XNOR2X1 port map( A => si_6_port, B => n351, Y => N447);
   U592 : NOR2X1 port map( A => si_6_port, B => n351, Y => n353);
   U594 : XOR2X1 port map( A => si_7_port, B => n353, Y => N448);
   U596 : INVX2 port map( A => si_3_port, Y => n355);
   U598 : INVX2 port map( A => si_1_port, Y => n357);
   U600 : INVX2 port map( A => n347, Y => N445);
   U602 : INVX2 port map( A => n341, Y => N443);
   U608 : INVX2 port map( A => KEY_ERROR, Y => n359);
   U611 : INVX2 port map( A => BYTE_READY, Y => n361);
   U614 : INVX2 port map( A => n130, Y => n363);
   U617 : INVX2 port map( A => OPCODE(1), Y => n365);
   U620 : INVX2 port map( A => OPCODE(0), Y => n367);
   U623 : INVX2 port map( A => nextProcessedData_7_port, Y => n369);
   U626 : INVX2 port map( A => n316, Y => n371);
   U627 : INVX2 port map( A => nextProcessedData_6_port, Y => n373);
   U629 : INVX2 port map( A => n325, Y => n375);
   U630 : INVX2 port map( A => nextProcessedData_5_port, Y => n377);
   U636 : INVX2 port map( A => n324, Y => n379);
   U640 : INVX2 port map( A => nextProcessedData_4_port, Y => n381);
   U642 : INVX2 port map( A => n323, Y => n383);
   U644 : INVX2 port map( A => nextProcessedData_3_port, Y => n385);
   U645 : INVX2 port map( A => n322, Y => n387);
   U648 : INVX2 port map( A => nextProcessedData_2_port, Y => n389);
   U651 : INVX2 port map( A => n321, Y => n391);
   U658 : INVX2 port map( A => nextProcessedData_1_port, Y => n393);
   U661 : INVX2 port map( A => n320, Y => n395);
   U670 : INVX2 port map( A => nextProcessedData_0_port, Y => n397);
   U671 : INVX2 port map( A => n319, Y => n399);
   U674 : INVX2 port map( A => prefillCounter_0_port, Y => n401);
   U675 : INVX2 port map( A => nfdata_0_port, Y => n403);
   U676 : INVX2 port map( A => nfaddr_0_port, Y => n405);
   U680 : INVX2 port map( A => n539, Y => n411_port);
   U682 : INVX2 port map( A => n538, Y => n413_port);
   U683 : INVX2 port map( A => n537, Y => n415);
   U687 : INVX2 port map( A => n536, Y => n417);
   U688 : INVX2 port map( A => n535, Y => n419);
   U689 : INVX2 port map( A => n534, Y => n421);
   U691 : INVX2 port map( A => n533, Y => n423);
   U695 : INVX2 port map( A => n530, Y => n425_port);
   U698 : INVX2 port map( A => n508, Y => n427_port);
   U701 : INVX2 port map( A => n502_port, Y => n429_port);
   U704 : INVX2 port map( A => n570, Y => n431_port);
   U707 : INVX2 port map( A => n590, Y => n433);
   U710 : INVX2 port map( A => n596, Y => n435);
   U713 : INVX2 port map( A => nfdata_7_port, Y => n437);
   U717 : INVX2 port map( A => nfdata_6_port, Y => n439);
   U718 : INVX2 port map( A => nfdata_5_port, Y => n441);
   U719 : INVX2 port map( A => nfdata_4_port, Y => n443_port);
   U720 : INVX2 port map( A => nfdata_3_port, Y => n445_port);
   U725 : INVX2 port map( A => nfdata_2_port, Y => n447_port);
   U726 : INVX2 port map( A => nfdata_1_port, Y => n449_port);
   U728 : INVX2 port map( A => n56, Y => n451_port);
   U729 : INVX2 port map( A => n486_port, Y => n453_port);
   U730 : INVX2 port map( A => n489, Y => n455_port);
   U734 : INVX2 port map( A => n490, Y => n458);
   U736 : INVX2 port map( A => n491, Y => n459);
   U740 : INVX2 port map( A => n492, Y => n461);
   U741 : INVX2 port map( A => n493, Y => n462);
   U742 : INVX2 port map( A => n494, Y => n463);
   U744 : INVX2 port map( A => n495, Y => n465);
   U747 : INVX2 port map( A => nfaddr_1_port, Y => n471);
   U749 : INVX2 port map( A => nfaddr_2_port, Y => n473_port);
   U753 : INVX2 port map( A => nfaddr_3_port, Y => n475_port);
   U756 : INVX2 port map( A => nfaddr_4_port, Y => n480_port);
   U758 : INVX2 port map( A => nfaddr_5_port, Y => n482_port);
   U763 : INVX2 port map( A => nfaddr_6_port, Y => n488);
   U768 : INVX2 port map( A => nfaddr_7_port, Y => n498_port);
   U770 : INVX2 port map( A => n310, Y => n500_port);
   U773 : INVX2 port map( A => n156, Y => n501_port);
   U776 : INVX2 port map( A => n118, Y => n503_port);
   U777 : INVX2 port map( A => n225, Y => n504);
   U778 : INVX2 port map( A => n315, Y => n505);
   U779 : INVX2 port map( A => n3, Y => n506);
   U782 : INVX2 port map( A => n485_port, Y => n509);
   U786 : INVX2 port map( A => n627, Y => n512_port);
   U789 : INVX2 port map( A => n229, Y => n514_port);
   U791 : INVX2 port map( A => n631, Y => n516_port);
   U793 : INVX2 port map( A => n157, Y => n518_port);
   U795 : INVX2 port map( A => n313, Y => n520_port);
   U796 : INVX2 port map( A => n148, Y => n522_port);
   U798 : INVX2 port map( A => n595, Y => n524_port);
   U802 : INVX2 port map( A => n205, Y => n528);
   U803 : INVX2 port map( A => n139, Y => n540);
   U805 : INVX2 port map( A => n53, Y => n541);
   U810 : INVX2 port map( A => n48, Y => n542);
   U811 : INVX2 port map( A => n43, Y => n543);
   U813 : INVX2 port map( A => n38, Y => n545);
   U814 : INVX2 port map( A => n33, Y => n547);
   U820 : INVX2 port map( A => n28, Y => n549);
   U821 : INVX2 port map( A => n23, Y => n551);
   U823 : INVX2 port map( A => n13, Y => n553);
   U824 : INVX2 port map( A => state_1_port, Y => n555);
   U830 : INVX2 port map( A => n567, Y => n557);
   U831 : INVX2 port map( A => n149, Y => n562);
   U833 : INVX2 port map( A => n625, Y => n569);
   U834 : INVX2 port map( A => n153, Y => n571);
   U840 : INVX2 port map( A => n112, Y => n577);
   U841 : INVX2 port map( A => n499_port, Y => n579);
   U843 : INVX2 port map( A => n115, Y => n592);
   U844 : INVX2 port map( A => n198, Y => n600);
   U850 : INVX2 port map( A => state_2_port, Y => n604);
   U851 : INVX2 port map( A => state_0_port, Y => n612);
   U853 : INVX2 port map( A => state_3_port, Y => n614);
   U854 : INVX2 port map( A => keyTable_7_0_port, Y => n616);
   U860 : INVX2 port map( A => keyTable_7_1_port, Y => n618);
   U861 : INVX2 port map( A => keyTable_7_2_port, Y => n624);
   U863 : INVX2 port map( A => keyTable_7_3_port, Y => n626);
   U864 : INVX2 port map( A => keyTable_7_4_port, Y => n629);
   U870 : INVX2 port map( A => keyTable_7_5_port, Y => n630);
   U871 : INVX2 port map( A => keyTable_7_6_port, Y => n632);
   U873 : INVX2 port map( A => keyTable_7_7_port, Y => n636);
   U874 : INVX2 port map( A => keyTable_6_0_port, Y => n637);
   U881 : INVX2 port map( A => keyTable_6_1_port, Y => n638);
   U883 : INVX2 port map( A => keyTable_6_2_port, Y => n648);
   U886 : INVX2 port map( A => keyTable_6_3_port, Y => n649);
   U888 : INVX2 port map( A => keyTable_6_4_port, Y => n650);
   U889 : INVX2 port map( A => keyTable_6_5_port, Y => n651);
   U891 : INVX2 port map( A => keyTable_6_6_port, Y => n692);
   U893 : INVX2 port map( A => keyTable_6_7_port, Y => n701);
   U895 : INVX2 port map( A => keyTable_5_0_port, Y => n746);
   U897 : INVX2 port map( A => keyTable_5_1_port, Y => n748);
   U899 : INVX2 port map( A => keyTable_5_2_port, Y => n750);
   U900 : INVX2 port map( A => keyTable_5_3_port, Y => n752);
   U902 : INVX2 port map( A => keyTable_5_4_port, Y => n754);
   U903 : INVX2 port map( A => keyTable_5_5_port, Y => n756);
   U904 : INVX2 port map( A => keyTable_5_6_port, Y => n758);
   U905 : INVX2 port map( A => keyTable_5_7_port, Y => n760);
   U906 : INVX2 port map( A => keyTable_4_0_port, Y => n761);
   U907 : INVX2 port map( A => keyTable_4_1_port, Y => n762);
   U908 : INVX2 port map( A => keyTable_4_2_port, Y => n763);
   U909 : INVX2 port map( A => keyTable_4_3_port, Y => n764);
   U910 : INVX2 port map( A => keyTable_4_4_port, Y => n765);
   U911 : INVX2 port map( A => keyTable_4_5_port, Y => n766);
   U912 : INVX2 port map( A => keyTable_4_6_port, Y => n767);
   U913 : INVX2 port map( A => keyTable_4_7_port, Y => n768);
   U914 : INVX2 port map( A => keyTable_3_0_port, Y => n769);
   U915 : INVX2 port map( A => keyTable_3_1_port, Y => n770);
   U916 : INVX2 port map( A => keyTable_3_2_port, Y => n771);
   U917 : INVX2 port map( A => keyTable_3_3_port, Y => n772);
   U918 : INVX2 port map( A => keyTable_3_4_port, Y => n773);
   U919 : INVX2 port map( A => keyTable_3_5_port, Y => n774);
   U920 : INVX2 port map( A => keyTable_3_6_port, Y => n775);
   U921 : INVX2 port map( A => keyTable_3_7_port, Y => n776);
   U922 : INVX2 port map( A => keyTable_2_0_port, Y => n777);
   U923 : INVX2 port map( A => keyTable_2_1_port, Y => n778);
   U924 : INVX2 port map( A => keyTable_2_2_port, Y => n779);
   U925 : INVX2 port map( A => keyTable_2_3_port, Y => n780);
   U926 : INVX2 port map( A => keyTable_2_4_port, Y => n781);
   U927 : INVX2 port map( A => keyTable_2_5_port, Y => n782);
   U928 : INVX2 port map( A => keyTable_2_6_port, Y => n783);
   U929 : INVX2 port map( A => keyTable_2_7_port, Y => n784);
   U930 : INVX2 port map( A => keyTable_1_0_port, Y => n785);
   U931 : INVX2 port map( A => keyTable_1_1_port, Y => n786);
   U932 : INVX2 port map( A => keyTable_1_2_port, Y => n787);
   U933 : INVX2 port map( A => keyTable_1_3_port, Y => n788);
   U934 : INVX2 port map( A => keyTable_1_4_port, Y => n789);
   U935 : INVX2 port map( A => keyTable_1_5_port, Y => n790);
   U936 : INVX2 port map( A => keyTable_1_6_port, Y => n791);
   U937 : INVX2 port map( A => keyTable_0_6_port, Y => n864);
   U938 : INVX2 port map( A => keyTable_0_5_port, Y => n865);
   U939 : INVX2 port map( A => keyTable_0_4_port, Y => n866);
   U940 : INVX2 port map( A => keyTable_0_3_port, Y => n867);
   U941 : INVX2 port map( A => keyTable_0_2_port, Y => n868);
   U942 : INVX2 port map( A => keyTable_0_1_port, Y => n869);
   U943 : INVX2 port map( A => keyTable_0_0_port, Y => n870);
   U944 : INVX2 port map( A => keyTable_1_7_port, Y => n871);
   U945 : INVX2 port map( A => keyTable_0_7_port, Y => n883);
   U946 : INVX2 port map( A => prefillCounter_7_port, Y => n884);
   U947 : INVX2 port map( A => prefillCounter_1_port, Y => n885);
   U948 : INVX2 port map( A => prefillCounter_2_port, Y => n886);
   U949 : INVX2 port map( A => prefillCounter_3_port, Y => n887);
   U950 : INVX2 port map( A => prefillCounter_4_port, Y => n888);
   U951 : INVX2 port map( A => prefillCounter_5_port, Y => n889);
   U952 : INVX2 port map( A => prefillCounter_6_port, Y => n890);
   U953 : INVX2 port map( A => temp_7_port, Y => n916);
   U954 : INVX2 port map( A => temp_0_port, Y => n917);
   U955 : INVX2 port map( A => temp_1_port, Y => n918);
   U956 : INVX2 port map( A => temp_2_port, Y => n919);
   U957 : INVX2 port map( A => temp_3_port, Y => n920);
   U958 : INVX2 port map( A => temp_4_port, Y => n921);
   U959 : INVX2 port map( A => temp_5_port, Y => n922);
   U960 : INVX2 port map( A => temp_6_port, Y => n923);
   U961 : INVX2 port map( A => si_0_port, Y => n924);
   U962 : INVX2 port map( A => si_2_port, Y => n925);
   U963 : INVX2 port map( A => si_4_port, Y => n926);
   U964 : INVX2 port map( A => si_5_port, Y => n927);
   U965 : INVX2 port map( A => si_6_port, Y => n928);
   U966 : INVX2 port map( A => si_7_port, Y => n929);
   U967 : INVX2 port map( A => intj_7_port, Y => n930);
   U968 : INVX2 port map( A => intj_0_port, Y => n931);
   U969 : INVX2 port map( A => intj_1_port, Y => n932);
   U970 : INVX2 port map( A => intj_2_port, Y => n933);
   U971 : INVX2 port map( A => intj_3_port, Y => n934);
   U972 : INVX2 port map( A => intj_4_port, Y => n935);
   U973 : INVX2 port map( A => intj_5_port, Y => n936);
   U974 : INVX2 port map( A => intj_6_port, Y => n937);
   U975 : INVX2 port map( A => sj_7_port, Y => n938);
   U976 : INVX2 port map( A => sj_6_port, Y => n939);
   U977 : INVX2 port map( A => sj_5_port, Y => n940);
   U978 : INVX2 port map( A => sj_4_port, Y => n941);
   U979 : INVX2 port map( A => sj_3_port, Y => n942);
   U980 : INVX2 port map( A => sj_2_port, Y => n943);
   U981 : INVX2 port map( A => sj_1_port, Y => n944);
   U982 : INVX2 port map( A => currentProcessedData_0_port, Y => n952);
   U983 : INVX2 port map( A => currentProcessedData_1_port, Y => n953);
   U984 : INVX2 port map( A => currentProcessedData_2_port, Y => n954);
   U985 : INVX2 port map( A => currentProcessedData_3_port, Y => n955);
   U986 : INVX2 port map( A => currentProcessedData_4_port, Y => n956);
   U987 : INVX2 port map( A => currentProcessedData_5_port, Y => n957);
   U988 : INVX2 port map( A => currentProcessedData_6_port, Y => n958);
   U989 : INVX2 port map( A => currentProcessedData_7_port, Y => n959);
   U990 : INVX2 port map( A => faddr_7_port, Y => n960);
   U991 : INVX2 port map( A => faddr_6_port, Y => n961);
   U992 : INVX2 port map( A => faddr_5_port, Y => n962);
   U993 : INVX2 port map( A => faddr_4_port, Y => n963);
   U994 : INVX2 port map( A => faddr_3_port, Y => n964);
   U995 : INVX2 port map( A => faddr_2_port, Y => n965);
   U996 : INVX2 port map( A => faddr_1_port, Y => n966);
   U997 : INVX2 port map( A => faddr_0_port, Y => n967);
   U998 : INVX2 port map( A => fdata_7_port, Y => n968);
   U999 : INVX2 port map( A => fdata_6_port, Y => n969);
   U1000 : INVX2 port map( A => fdata_5_port, Y => n970);
   U1001 : INVX2 port map( A => fdata_4_port, Y => n971);
   U1002 : INVX2 port map( A => fdata_3_port, Y => n972);
   U1003 : INVX2 port map( A => fdata_2_port, Y => n973);
   U1004 : INVX2 port map( A => fdata_1_port, Y => n974);
   U1005 : INVX2 port map( A => fdata_0_port, Y => n975);
   n976 <= '0';
   n977 <= '0';

end SYN_bksa;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity transmitter_block_1 is

   port( PRGA_OUT : in std_logic_vector (7 downto 0);  clk, p_ready : in 
         std_logic;  prga_opcode : in std_logic_vector (1 downto 0);  rst : in 
         std_logic;  SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE : out std_logic);

end transmitter_block_1;

architecture SYN_struct of transmitter_block_1 is

   component tx_timer_1
      port( CLK, RST, SENDING : in std_logic;  SHIFT_ENABLE_R, SHIFT_ENABLE_E :
            out std_logic);
   end component;
   
   component tx_tcu_1
      port( clk, rst, p_ready, t_bitstuff : in std_logic;  PRGA_OUT : in 
            std_logic_vector (7 downto 0);  prga_opcode : in std_logic_vector 
            (1 downto 0);  t_crc : in std_logic_vector (15 downto 0);  sending,
            EOP, next_byte : out std_logic;  send_data : out std_logic_vector 
            (7 downto 0);  t_strobe : out std_logic);
   end component;
   
   component tx_shiftreg_1
      port( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe : in std_logic;  
            send_data : in std_logic_vector (7 downto 0);  d_encode : out 
            std_logic);
   end component;
   
   component tx_encode_1
      port( clk, rst, SHIFT_ENABLE_E, d_encode, EOP : in std_logic;  t_bitstuff
            , dp_tx_out, dm_tx_out : out std_logic);
   end component;
   
   component tx_CRC_CALC_1
      port( CLK, RST, EOP, T_STROBE : in std_logic;  PRGA_OPCODE : in 
            std_logic_vector (1 downto 0);  PRGA_OUT : in std_logic_vector (7 
            downto 0);  TX_CRC : out std_logic_vector (15 downto 0));
   end component;
   
   signal SENDING_port, t_strobe, EOP, TX_CRC_15_port, TX_CRC_14_port, 
      TX_CRC_13_port, TX_CRC_12_port, TX_CRC_11_port, TX_CRC_10_port, 
      TX_CRC_9_port, TX_CRC_8_port, TX_CRC_7_port, TX_CRC_6_port, TX_CRC_5_port
      , TX_CRC_4_port, TX_CRC_3_port, TX_CRC_2_port, TX_CRC_1_port, 
      TX_CRC_0_port, SHIFT_ENABLE_E, d_encode, t_bitstuff, SHIFT_ENABLE_R, 
      send_data_7_port, send_data_6_port, send_data_5_port, send_data_4_port, 
      send_data_3_port, send_data_2_port, send_data_1_port, send_data_0_port : 
      std_logic;

begin
   SENDING <= SENDING_port;
   
   U_1 : tx_CRC_CALC_1 port map( CLK => clk, RST => rst, EOP => EOP, T_STROBE 
                           => t_strobe, PRGA_OPCODE(1) => prga_opcode(1), 
                           PRGA_OPCODE(0) => prga_opcode(0), PRGA_OUT(7) => 
                           PRGA_OUT(7), PRGA_OUT(6) => PRGA_OUT(6), PRGA_OUT(5)
                           => PRGA_OUT(5), PRGA_OUT(4) => PRGA_OUT(4), 
                           PRGA_OUT(3) => PRGA_OUT(3), PRGA_OUT(2) => 
                           PRGA_OUT(2), PRGA_OUT(1) => PRGA_OUT(1), PRGA_OUT(0)
                           => PRGA_OUT(0), TX_CRC(15) => TX_CRC_15_port, 
                           TX_CRC(14) => TX_CRC_14_port, TX_CRC(13) => 
                           TX_CRC_13_port, TX_CRC(12) => TX_CRC_12_port, 
                           TX_CRC(11) => TX_CRC_11_port, TX_CRC(10) => 
                           TX_CRC_10_port, TX_CRC(9) => TX_CRC_9_port, 
                           TX_CRC(8) => TX_CRC_8_port, TX_CRC(7) => 
                           TX_CRC_7_port, TX_CRC(6) => TX_CRC_6_port, TX_CRC(5)
                           => TX_CRC_5_port, TX_CRC(4) => TX_CRC_4_port, 
                           TX_CRC(3) => TX_CRC_3_port, TX_CRC(2) => 
                           TX_CRC_2_port, TX_CRC(1) => TX_CRC_1_port, TX_CRC(0)
                           => TX_CRC_0_port);
   U_0 : tx_encode_1 port map( clk => clk, rst => rst, SHIFT_ENABLE_E => 
                           SHIFT_ENABLE_E, d_encode => d_encode, EOP => EOP, 
                           t_bitstuff => t_bitstuff, dp_tx_out => dp_tx_out, 
                           dm_tx_out => dm_tx_out);
   U_2 : tx_shiftreg_1 port map( clk => clk, rst => rst, SHIFT_ENABLE_R => 
                           SHIFT_ENABLE_R, t_bitstuff => t_bitstuff, t_strobe 
                           => t_strobe, send_data(7) => send_data_7_port, 
                           send_data(6) => send_data_6_port, send_data(5) => 
                           send_data_5_port, send_data(4) => send_data_4_port, 
                           send_data(3) => send_data_3_port, send_data(2) => 
                           send_data_2_port, send_data(1) => send_data_1_port, 
                           send_data(0) => send_data_0_port, d_encode => 
                           d_encode);
   U_3 : tx_tcu_1 port map( clk => clk, rst => rst, p_ready => p_ready, 
                           t_bitstuff => t_bitstuff, PRGA_OUT(7) => PRGA_OUT(7)
                           , PRGA_OUT(6) => PRGA_OUT(6), PRGA_OUT(5) => 
                           PRGA_OUT(5), PRGA_OUT(4) => PRGA_OUT(4), PRGA_OUT(3)
                           => PRGA_OUT(3), PRGA_OUT(2) => PRGA_OUT(2), 
                           PRGA_OUT(1) => PRGA_OUT(1), PRGA_OUT(0) => 
                           PRGA_OUT(0), prga_opcode(1) => prga_opcode(1), 
                           prga_opcode(0) => prga_opcode(0), t_crc(15) => 
                           TX_CRC_15_port, t_crc(14) => TX_CRC_14_port, 
                           t_crc(13) => TX_CRC_13_port, t_crc(12) => 
                           TX_CRC_12_port, t_crc(11) => TX_CRC_11_port, 
                           t_crc(10) => TX_CRC_10_port, t_crc(9) => 
                           TX_CRC_9_port, t_crc(8) => TX_CRC_8_port, t_crc(7) 
                           => TX_CRC_7_port, t_crc(6) => TX_CRC_6_port, 
                           t_crc(5) => TX_CRC_5_port, t_crc(4) => TX_CRC_4_port
                           , t_crc(3) => TX_CRC_3_port, t_crc(2) => 
                           TX_CRC_2_port, t_crc(1) => TX_CRC_1_port, t_crc(0) 
                           => TX_CRC_0_port, sending => SENDING_port, EOP => 
                           EOP, next_byte => NEXT_BYTE, send_data(7) => 
                           send_data_7_port, send_data(6) => send_data_6_port, 
                           send_data(5) => send_data_5_port, send_data(4) => 
                           send_data_4_port, send_data(3) => send_data_3_port, 
                           send_data(2) => send_data_2_port, send_data(1) => 
                           send_data_1_port, send_data(0) => send_data_0_port, 
                           t_strobe => t_strobe);
   U_4 : tx_timer_1 port map( CLK => clk, RST => rst, SENDING => SENDING_port, 
                           SHIFT_ENABLE_R => SHIFT_ENABLE_R, SHIFT_ENABLE_E => 
                           SHIFT_ENABLE_E);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity receiver_block_rewire_1 is

   port( CLK, DM1_RX, DP1_RX, RST : in std_logic;  BS_ERROR, CRC_ERROR, 
         EOP_external : out std_logic;  OPCODE : out std_logic_vector (1 downto
         0);  RCV_DATA : out std_logic_vector (7 downto 0);  R_ERROR, W_ENABLE 
         : out std_logic);

end receiver_block_rewire_1;

architecture SYN_struct of receiver_block_rewire_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component rx_timer_1
      port( CLK, RST, D_EDGE, RCVING : in std_logic;  SHIFT_ENABLE : out 
            std_logic);
   end component;
   
   component rx_shift_reg_1
      port( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF : in std_logic;  RCV_DATA 
            : out std_logic_vector (7 downto 0));
   end component;
   
   component rx_rcu_1
      port( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR : in 
            std_logic;  RX_CRC, RX_CHECK_CRC : in std_logic_vector (15 downto 
            0);  RCV_DATA : in std_logic_vector (7 downto 0);  RCVING, W_ENABLE
            , R_ERROR, CRC_ERROR : out std_logic;  OPCODE : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component rx_eopdetect_1
      port( DP1_RX, DM1_RX : in std_logic;  EOP : out std_logic);
   end component;
   
   component rx_edgedetect_1
      port( CLK, RST, DP1_RX : in std_logic;  D_EDGE : out std_logic);
   end component;
   
   component rx_decode_1
      port( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP : in std_logic;  D_ORIG, 
            BITSTUFF, BS_ERROR : out std_logic);
   end component;
   
   component rx_accumulator_1
      port( CLK, RST : in std_logic;  RCV_DATA : in std_logic_vector (7 downto 
            0);  W_ENABLE : in std_logic;  rx_CHECK_CRC : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component rx_CRC_CALC_1
      port( CLK, RST, W_ENABLE : in std_logic;  OPCODE : in std_logic_vector (1
            downto 0);  RCV_DATA : in std_logic_vector (7 downto 0);  RX_CRC : 
            out std_logic_vector (15 downto 0));
   end component;
   
   signal BS_ERROR_port, EOP_external_port, OPCODE_1_port, OPCODE_0_port, 
      RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      W_ENABLE_port, RX_CRC_15_port, RX_CRC_14_port, RX_CRC_13_port, 
      RX_CRC_12_port, RX_CRC_11_port, RX_CRC_10_port, RX_CRC_9_port, 
      RX_CRC_8_port, RX_CRC_7_port, RX_CRC_6_port, RX_CRC_5_port, RX_CRC_4_port
      , RX_CRC_3_port, RX_CRC_2_port, RX_CRC_1_port, RX_CRC_0_port, 
      rx_CHECK_CRC_15_port, rx_CHECK_CRC_14_port, rx_CHECK_CRC_13_port, 
      rx_CHECK_CRC_12_port, rx_CHECK_CRC_11_port, rx_CHECK_CRC_10_port, 
      rx_CHECK_CRC_9_port, rx_CHECK_CRC_8_port, rx_CHECK_CRC_7_port, 
      rx_CHECK_CRC_6_port, rx_CHECK_CRC_5_port, rx_CHECK_CRC_4_port, 
      rx_CHECK_CRC_3_port, rx_CHECK_CRC_2_port, rx_CHECK_CRC_1_port, 
      rx_CHECK_CRC_0_port, SHIFT_ENABLE, BITSTUFF, D_ORIG, D_EDGE, RCVING, n1, 
      n2 : std_logic;

begin
   BS_ERROR <= BS_ERROR_port;
   EOP_external <= EOP_external_port;
   OPCODE <= ( OPCODE_1_port, OPCODE_0_port );
   RCV_DATA <= ( RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, 
      RCV_DATA_4_port, RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, 
      RCV_DATA_0_port );
   W_ENABLE <= W_ENABLE_port;
   
   U_2 : rx_CRC_CALC_1 port map( CLK => CLK, RST => n1, W_ENABLE => 
                           W_ENABLE_port, OPCODE(1) => OPCODE_1_port, OPCODE(0)
                           => OPCODE_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, RX_CRC(15) => 
                           RX_CRC_15_port, RX_CRC(14) => RX_CRC_14_port, 
                           RX_CRC(13) => RX_CRC_13_port, RX_CRC(12) => 
                           RX_CRC_12_port, RX_CRC(11) => RX_CRC_11_port, 
                           RX_CRC(10) => RX_CRC_10_port, RX_CRC(9) => 
                           RX_CRC_9_port, RX_CRC(8) => RX_CRC_8_port, RX_CRC(7)
                           => RX_CRC_7_port, RX_CRC(6) => RX_CRC_6_port, 
                           RX_CRC(5) => RX_CRC_5_port, RX_CRC(4) => 
                           RX_CRC_4_port, RX_CRC(3) => RX_CRC_3_port, RX_CRC(2)
                           => RX_CRC_2_port, RX_CRC(1) => RX_CRC_1_port, 
                           RX_CRC(0) => RX_CRC_0_port);
   U_3 : rx_accumulator_1 port map( CLK => CLK, RST => n1, RCV_DATA(7) => 
                           RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           W_ENABLE => W_ENABLE_port, rx_CHECK_CRC(15) => 
                           rx_CHECK_CRC_15_port, rx_CHECK_CRC(14) => 
                           rx_CHECK_CRC_14_port, rx_CHECK_CRC(13) => 
                           rx_CHECK_CRC_13_port, rx_CHECK_CRC(12) => 
                           rx_CHECK_CRC_12_port, rx_CHECK_CRC(11) => 
                           rx_CHECK_CRC_11_port, rx_CHECK_CRC(10) => 
                           rx_CHECK_CRC_10_port, rx_CHECK_CRC(9) => 
                           rx_CHECK_CRC_9_port, rx_CHECK_CRC(8) => 
                           rx_CHECK_CRC_8_port, rx_CHECK_CRC(7) => 
                           rx_CHECK_CRC_7_port, rx_CHECK_CRC(6) => 
                           rx_CHECK_CRC_6_port, rx_CHECK_CRC(5) => 
                           rx_CHECK_CRC_5_port, rx_CHECK_CRC(4) => 
                           rx_CHECK_CRC_4_port, rx_CHECK_CRC(3) => 
                           rx_CHECK_CRC_3_port, rx_CHECK_CRC(2) => 
                           rx_CHECK_CRC_2_port, rx_CHECK_CRC(1) => 
                           rx_CHECK_CRC_1_port, rx_CHECK_CRC(0) => 
                           rx_CHECK_CRC_0_port);
   U_1 : rx_decode_1 port map( CLK => CLK, RST => n1, DP1_RX => DP1_RX, 
                           SHIFT_ENABLE => SHIFT_ENABLE, EOP => 
                           EOP_external_port, D_ORIG => D_ORIG, BITSTUFF => 
                           BITSTUFF, BS_ERROR => BS_ERROR_port);
   U_0 : rx_edgedetect_1 port map( CLK => CLK, RST => n1, DP1_RX => DP1_RX, 
                           D_EDGE => D_EDGE);
   U_4 : rx_eopdetect_1 port map( DP1_RX => DP1_RX, DM1_RX => DM1_RX, EOP => 
                           EOP_external_port);
   U_5 : rx_rcu_1 port map( CLK => CLK, RST => n1, D_EDGE => D_EDGE, EOP => 
                           EOP_external_port, SHIFT_ENABLE => SHIFT_ENABLE, 
                           BITSTUFF => BITSTUFF, BS_ERROR => BS_ERROR_port, 
                           RX_CRC(15) => RX_CRC_15_port, RX_CRC(14) => 
                           RX_CRC_14_port, RX_CRC(13) => RX_CRC_13_port, 
                           RX_CRC(12) => RX_CRC_12_port, RX_CRC(11) => 
                           RX_CRC_11_port, RX_CRC(10) => RX_CRC_10_port, 
                           RX_CRC(9) => RX_CRC_9_port, RX_CRC(8) => 
                           RX_CRC_8_port, RX_CRC(7) => RX_CRC_7_port, RX_CRC(6)
                           => RX_CRC_6_port, RX_CRC(5) => RX_CRC_5_port, 
                           RX_CRC(4) => RX_CRC_4_port, RX_CRC(3) => 
                           RX_CRC_3_port, RX_CRC(2) => RX_CRC_2_port, RX_CRC(1)
                           => RX_CRC_1_port, RX_CRC(0) => RX_CRC_0_port, 
                           RX_CHECK_CRC(15) => rx_CHECK_CRC_15_port, 
                           RX_CHECK_CRC(14) => rx_CHECK_CRC_14_port, 
                           RX_CHECK_CRC(13) => rx_CHECK_CRC_13_port, 
                           RX_CHECK_CRC(12) => rx_CHECK_CRC_12_port, 
                           RX_CHECK_CRC(11) => rx_CHECK_CRC_11_port, 
                           RX_CHECK_CRC(10) => rx_CHECK_CRC_10_port, 
                           RX_CHECK_CRC(9) => rx_CHECK_CRC_9_port, 
                           RX_CHECK_CRC(8) => rx_CHECK_CRC_8_port, 
                           RX_CHECK_CRC(7) => rx_CHECK_CRC_7_port, 
                           RX_CHECK_CRC(6) => rx_CHECK_CRC_6_port, 
                           RX_CHECK_CRC(5) => rx_CHECK_CRC_5_port, 
                           RX_CHECK_CRC(4) => rx_CHECK_CRC_4_port, 
                           RX_CHECK_CRC(3) => rx_CHECK_CRC_3_port, 
                           RX_CHECK_CRC(2) => rx_CHECK_CRC_2_port, 
                           RX_CHECK_CRC(1) => rx_CHECK_CRC_1_port, 
                           RX_CHECK_CRC(0) => rx_CHECK_CRC_0_port, RCV_DATA(7) 
                           => RCV_DATA_7_port, RCV_DATA(6) => RCV_DATA_6_port, 
                           RCV_DATA(5) => RCV_DATA_5_port, RCV_DATA(4) => 
                           RCV_DATA_4_port, RCV_DATA(3) => RCV_DATA_3_port, 
                           RCV_DATA(2) => RCV_DATA_2_port, RCV_DATA(1) => 
                           RCV_DATA_1_port, RCV_DATA(0) => RCV_DATA_0_port, 
                           RCVING => RCVING, W_ENABLE => W_ENABLE_port, R_ERROR
                           => R_ERROR, CRC_ERROR => CRC_ERROR, OPCODE(1) => 
                           OPCODE_1_port, OPCODE(0) => OPCODE_0_port);
   U_6 : rx_shift_reg_1 port map( CLK => CLK, RST => n1, SHIFT_ENABLE => 
                           SHIFT_ENABLE, D_ORIG => D_ORIG, BITSTUFF => BITSTUFF
                           , RCV_DATA(7) => RCV_DATA_7_port, RCV_DATA(6) => 
                           RCV_DATA_6_port, RCV_DATA(5) => RCV_DATA_5_port, 
                           RCV_DATA(4) => RCV_DATA_4_port, RCV_DATA(3) => 
                           RCV_DATA_3_port, RCV_DATA(2) => RCV_DATA_2_port, 
                           RCV_DATA(1) => RCV_DATA_1_port, RCV_DATA(0) => 
                           RCV_DATA_0_port);
   U_7 : rx_timer_1 port map( CLK => CLK, RST => n1, D_EDGE => D_EDGE, RCVING 
                           => RCVING, SHIFT_ENABLE => SHIFT_ENABLE);
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity memoryblock_1 is

   port( CLK, NEXT_BYTE : in std_logic;  RCV_DATA : in std_logic_vector (7 
         downto 0);  RCV_OPCODE : in std_logic_vector (1 downto 0);  RST, 
         W_ENABLE, EOP : in std_logic;  EMPTY, FULL, B_READY : out std_logic;  
         PRGA_IN : out std_logic_vector (7 downto 0);  PRGA_OPCODE : out 
         std_logic_vector (1 downto 0));

end memoryblock_1;

architecture SYN_struct of memoryblock_1 is

   component RFIFO_1
      port( CLK, RST, W_ENABLE, R_ENABLE : in std_logic;  RCV_DATA : in 
            std_logic_vector (7 downto 0);  RCV_OPCODE : in std_logic_vector (1
            downto 0);  DATA : out std_logic_vector (7 downto 0);  OUT_OPCODE :
            out std_logic_vector (1 downto 0);  BYTE_COUNT : out 
            std_logic_vector (4 downto 0);  EMPTY, FULL : out std_logic);
   end component;
   
   component RBUFFER_1
      port( CLK, RST, NEXT_BYTE : in std_logic;  DATA : in std_logic_vector (7 
            downto 0);  OPCODE : in std_logic_vector (1 downto 0);  BYTE_COUNT 
            : in std_logic_vector (4 downto 0);  EOP : in std_logic;  B_READY, 
            R_ENABLE : out std_logic;  PRGA_IN : out std_logic_vector (7 downto
            0);  PRGA_OPCODE : out std_logic_vector (1 downto 0));
   end component;
   
   signal BYTE_COUNT_4_port, BYTE_COUNT_3_port, BYTE_COUNT_2_port, 
      BYTE_COUNT_1_port, BYTE_COUNT_0_port, DATA_7_port, DATA_6_port, 
      DATA_5_port, DATA_4_port, DATA_3_port, DATA_2_port, DATA_1_port, 
      DATA_0_port, OUT_OPCODE_1_port, OUT_OPCODE_0_port, R_ENABLE : std_logic;

begin
   
   U_0 : RBUFFER_1 port map( CLK => CLK, RST => RST, NEXT_BYTE => NEXT_BYTE, 
                           DATA(7) => DATA_7_port, DATA(6) => DATA_6_port, 
                           DATA(5) => DATA_5_port, DATA(4) => DATA_4_port, 
                           DATA(3) => DATA_3_port, DATA(2) => DATA_2_port, 
                           DATA(1) => DATA_1_port, DATA(0) => DATA_0_port, 
                           OPCODE(1) => OUT_OPCODE_1_port, OPCODE(0) => 
                           OUT_OPCODE_0_port, BYTE_COUNT(4) => 
                           BYTE_COUNT_4_port, BYTE_COUNT(3) => 
                           BYTE_COUNT_3_port, BYTE_COUNT(2) => 
                           BYTE_COUNT_2_port, BYTE_COUNT(1) => 
                           BYTE_COUNT_1_port, BYTE_COUNT(0) => 
                           BYTE_COUNT_0_port, EOP => EOP, B_READY => B_READY, 
                           R_ENABLE => R_ENABLE, PRGA_IN(7) => PRGA_IN(7), 
                           PRGA_IN(6) => PRGA_IN(6), PRGA_IN(5) => PRGA_IN(5), 
                           PRGA_IN(4) => PRGA_IN(4), PRGA_IN(3) => PRGA_IN(3), 
                           PRGA_IN(2) => PRGA_IN(2), PRGA_IN(1) => PRGA_IN(1), 
                           PRGA_IN(0) => PRGA_IN(0), PRGA_OPCODE(1) => 
                           PRGA_OPCODE(1), PRGA_OPCODE(0) => PRGA_OPCODE(0));
   U_1 : RFIFO_1 port map( CLK => CLK, RST => RST, W_ENABLE => W_ENABLE, 
                           R_ENABLE => R_ENABLE, RCV_DATA(7) => RCV_DATA(7), 
                           RCV_DATA(6) => RCV_DATA(6), RCV_DATA(5) => 
                           RCV_DATA(5), RCV_DATA(4) => RCV_DATA(4), RCV_DATA(3)
                           => RCV_DATA(3), RCV_DATA(2) => RCV_DATA(2), 
                           RCV_DATA(1) => RCV_DATA(1), RCV_DATA(0) => 
                           RCV_DATA(0), RCV_OPCODE(1) => RCV_OPCODE(1), 
                           RCV_OPCODE(0) => RCV_OPCODE(0), DATA(7) => 
                           DATA_7_port, DATA(6) => DATA_6_port, DATA(5) => 
                           DATA_5_port, DATA(4) => DATA_4_port, DATA(3) => 
                           DATA_3_port, DATA(2) => DATA_2_port, DATA(1) => 
                           DATA_1_port, DATA(0) => DATA_0_port, OUT_OPCODE(1) 
                           => OUT_OPCODE_1_port, OUT_OPCODE(0) => 
                           OUT_OPCODE_0_port, BYTE_COUNT(4) => 
                           BYTE_COUNT_4_port, BYTE_COUNT(3) => 
                           BYTE_COUNT_3_port, BYTE_COUNT(2) => 
                           BYTE_COUNT_2_port, BYTE_COUNT(1) => 
                           BYTE_COUNT_1_port, BYTE_COUNT(0) => 
                           BYTE_COUNT_0_port, EMPTY => EMPTY, FULL => FULL);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity EDBlock_1 is

   port( BYTE : in std_logic_vector (7 downto 0);  BYTE_READY, CLK : in 
         std_logic;  OPCODE : in std_logic_vector (1 downto 0);  RST, SERIAL_IN
         : in std_logic;  DATA_IN : in std_logic_vector (7 downto 0);  
         KEY_ERROR, PARITY_ERROR, PDATA_READY : out std_logic;  PROCESSED_DATA 
         : out std_logic_vector (7 downto 0);  PROG_ERROR, RBUF_FULL, W_ENABLE,
         R_ENABLE : out std_logic;  DATA, ADDR : out std_logic_vector (7 downto
         0));

end EDBlock_1;

architecture SYN_struct of EDBlock_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component uart_rcv_block_1
      port( CLK, RST, SERIAL_IN : in std_logic;  KEY_ERROR, PROG_ERROR : out 
            std_logic;  PLAINKEY : out std_logic_vector (63 downto 0);  
            RBUF_FULL, PARITY_ERROR : out std_logic);
   end component;
   
   component KSA_1
      port( KEY : in std_logic_vector (63 downto 0);  CLK, RST, KEY_ERROR, 
            BYTE_READY : in std_logic;  BYTE : in std_logic_vector (7 downto 0)
            ;  OPCODE : in std_logic_vector (1 downto 0);  DATA_IN : in 
            std_logic_vector (7 downto 0);  PROCESSED_DATA : out 
            std_logic_vector (7 downto 0);  PDATA_READY, W_ENABLE, R_ENABLE : 
            out std_logic;  ADDR, DATA : out std_logic_vector (7 downto 0));
   end component;
   
   signal KEY_ERROR_port, PLAINKEY_63_port, PLAINKEY_62_port, PLAINKEY_61_port,
      PLAINKEY_60_port, PLAINKEY_59_port, PLAINKEY_58_port, PLAINKEY_57_port, 
      PLAINKEY_56_port, PLAINKEY_55_port, PLAINKEY_54_port, PLAINKEY_53_port, 
      PLAINKEY_52_port, PLAINKEY_51_port, PLAINKEY_50_port, PLAINKEY_49_port, 
      PLAINKEY_48_port, PLAINKEY_47_port, PLAINKEY_46_port, PLAINKEY_45_port, 
      PLAINKEY_44_port, PLAINKEY_43_port, PLAINKEY_42_port, PLAINKEY_41_port, 
      PLAINKEY_40_port, PLAINKEY_39_port, PLAINKEY_38_port, PLAINKEY_37_port, 
      PLAINKEY_36_port, PLAINKEY_35_port, PLAINKEY_34_port, PLAINKEY_33_port, 
      PLAINKEY_32_port, PLAINKEY_31_port, PLAINKEY_30_port, PLAINKEY_29_port, 
      PLAINKEY_28_port, PLAINKEY_27_port, PLAINKEY_26_port, PLAINKEY_25_port, 
      PLAINKEY_24_port, PLAINKEY_23_port, PLAINKEY_22_port, PLAINKEY_21_port, 
      PLAINKEY_20_port, PLAINKEY_19_port, PLAINKEY_18_port, PLAINKEY_17_port, 
      PLAINKEY_16_port, PLAINKEY_15_port, PLAINKEY_14_port, PLAINKEY_13_port, 
      PLAINKEY_12_port, PLAINKEY_11_port, PLAINKEY_10_port, PLAINKEY_9_port, 
      PLAINKEY_8_port, PLAINKEY_7_port, PLAINKEY_6_port, PLAINKEY_5_port, 
      PLAINKEY_4_port, PLAINKEY_3_port, PLAINKEY_2_port, PLAINKEY_1_port, 
      PLAINKEY_0_port, n1, n2 : std_logic;

begin
   KEY_ERROR <= KEY_ERROR_port;
   
   U_0 : KSA_1 port map( KEY(63) => PLAINKEY_63_port, KEY(62) => 
                           PLAINKEY_62_port, KEY(61) => PLAINKEY_61_port, 
                           KEY(60) => PLAINKEY_60_port, KEY(59) => 
                           PLAINKEY_59_port, KEY(58) => PLAINKEY_58_port, 
                           KEY(57) => PLAINKEY_57_port, KEY(56) => 
                           PLAINKEY_56_port, KEY(55) => PLAINKEY_55_port, 
                           KEY(54) => PLAINKEY_54_port, KEY(53) => 
                           PLAINKEY_53_port, KEY(52) => PLAINKEY_52_port, 
                           KEY(51) => PLAINKEY_51_port, KEY(50) => 
                           PLAINKEY_50_port, KEY(49) => PLAINKEY_49_port, 
                           KEY(48) => PLAINKEY_48_port, KEY(47) => 
                           PLAINKEY_47_port, KEY(46) => PLAINKEY_46_port, 
                           KEY(45) => PLAINKEY_45_port, KEY(44) => 
                           PLAINKEY_44_port, KEY(43) => PLAINKEY_43_port, 
                           KEY(42) => PLAINKEY_42_port, KEY(41) => 
                           PLAINKEY_41_port, KEY(40) => PLAINKEY_40_port, 
                           KEY(39) => PLAINKEY_39_port, KEY(38) => 
                           PLAINKEY_38_port, KEY(37) => PLAINKEY_37_port, 
                           KEY(36) => PLAINKEY_36_port, KEY(35) => 
                           PLAINKEY_35_port, KEY(34) => PLAINKEY_34_port, 
                           KEY(33) => PLAINKEY_33_port, KEY(32) => 
                           PLAINKEY_32_port, KEY(31) => PLAINKEY_31_port, 
                           KEY(30) => PLAINKEY_30_port, KEY(29) => 
                           PLAINKEY_29_port, KEY(28) => PLAINKEY_28_port, 
                           KEY(27) => PLAINKEY_27_port, KEY(26) => 
                           PLAINKEY_26_port, KEY(25) => PLAINKEY_25_port, 
                           KEY(24) => PLAINKEY_24_port, KEY(23) => 
                           PLAINKEY_23_port, KEY(22) => PLAINKEY_22_port, 
                           KEY(21) => PLAINKEY_21_port, KEY(20) => 
                           PLAINKEY_20_port, KEY(19) => PLAINKEY_19_port, 
                           KEY(18) => PLAINKEY_18_port, KEY(17) => 
                           PLAINKEY_17_port, KEY(16) => PLAINKEY_16_port, 
                           KEY(15) => PLAINKEY_15_port, KEY(14) => 
                           PLAINKEY_14_port, KEY(13) => PLAINKEY_13_port, 
                           KEY(12) => PLAINKEY_12_port, KEY(11) => 
                           PLAINKEY_11_port, KEY(10) => PLAINKEY_10_port, 
                           KEY(9) => PLAINKEY_9_port, KEY(8) => PLAINKEY_8_port
                           , KEY(7) => PLAINKEY_7_port, KEY(6) => 
                           PLAINKEY_6_port, KEY(5) => PLAINKEY_5_port, KEY(4) 
                           => PLAINKEY_4_port, KEY(3) => PLAINKEY_3_port, 
                           KEY(2) => PLAINKEY_2_port, KEY(1) => PLAINKEY_1_port
                           , KEY(0) => PLAINKEY_0_port, CLK => CLK, RST => n1, 
                           KEY_ERROR => KEY_ERROR_port, BYTE_READY => 
                           BYTE_READY, BYTE(7) => BYTE(7), BYTE(6) => BYTE(6), 
                           BYTE(5) => BYTE(5), BYTE(4) => BYTE(4), BYTE(3) => 
                           BYTE(3), BYTE(2) => BYTE(2), BYTE(1) => BYTE(1), 
                           BYTE(0) => BYTE(0), OPCODE(1) => OPCODE(1), 
                           OPCODE(0) => OPCODE(0), DATA_IN(7) => DATA_IN(7), 
                           DATA_IN(6) => DATA_IN(6), DATA_IN(5) => DATA_IN(5), 
                           DATA_IN(4) => DATA_IN(4), DATA_IN(3) => DATA_IN(3), 
                           DATA_IN(2) => DATA_IN(2), DATA_IN(1) => DATA_IN(1), 
                           DATA_IN(0) => DATA_IN(0), PROCESSED_DATA(7) => 
                           PROCESSED_DATA(7), PROCESSED_DATA(6) => 
                           PROCESSED_DATA(6), PROCESSED_DATA(5) => 
                           PROCESSED_DATA(5), PROCESSED_DATA(4) => 
                           PROCESSED_DATA(4), PROCESSED_DATA(3) => 
                           PROCESSED_DATA(3), PROCESSED_DATA(2) => 
                           PROCESSED_DATA(2), PROCESSED_DATA(1) => 
                           PROCESSED_DATA(1), PROCESSED_DATA(0) => 
                           PROCESSED_DATA(0), PDATA_READY => PDATA_READY, 
                           W_ENABLE => W_ENABLE, R_ENABLE => R_ENABLE, ADDR(7) 
                           => ADDR(7), ADDR(6) => ADDR(6), ADDR(5) => ADDR(5), 
                           ADDR(4) => ADDR(4), ADDR(3) => ADDR(3), ADDR(2) => 
                           ADDR(2), ADDR(1) => ADDR(1), ADDR(0) => ADDR(0), 
                           DATA(7) => DATA(7), DATA(6) => DATA(6), DATA(5) => 
                           DATA(5), DATA(4) => DATA(4), DATA(3) => DATA(3), 
                           DATA(2) => DATA(2), DATA(1) => DATA(1), DATA(0) => 
                           DATA(0));
   U_1 : uart_rcv_block_1 port map( CLK => CLK, RST => n1, SERIAL_IN => 
                           SERIAL_IN, KEY_ERROR => KEY_ERROR_port, PROG_ERROR 
                           => PROG_ERROR, PLAINKEY(63) => PLAINKEY_63_port, 
                           PLAINKEY(62) => PLAINKEY_62_port, PLAINKEY(61) => 
                           PLAINKEY_61_port, PLAINKEY(60) => PLAINKEY_60_port, 
                           PLAINKEY(59) => PLAINKEY_59_port, PLAINKEY(58) => 
                           PLAINKEY_58_port, PLAINKEY(57) => PLAINKEY_57_port, 
                           PLAINKEY(56) => PLAINKEY_56_port, PLAINKEY(55) => 
                           PLAINKEY_55_port, PLAINKEY(54) => PLAINKEY_54_port, 
                           PLAINKEY(53) => PLAINKEY_53_port, PLAINKEY(52) => 
                           PLAINKEY_52_port, PLAINKEY(51) => PLAINKEY_51_port, 
                           PLAINKEY(50) => PLAINKEY_50_port, PLAINKEY(49) => 
                           PLAINKEY_49_port, PLAINKEY(48) => PLAINKEY_48_port, 
                           PLAINKEY(47) => PLAINKEY_47_port, PLAINKEY(46) => 
                           PLAINKEY_46_port, PLAINKEY(45) => PLAINKEY_45_port, 
                           PLAINKEY(44) => PLAINKEY_44_port, PLAINKEY(43) => 
                           PLAINKEY_43_port, PLAINKEY(42) => PLAINKEY_42_port, 
                           PLAINKEY(41) => PLAINKEY_41_port, PLAINKEY(40) => 
                           PLAINKEY_40_port, PLAINKEY(39) => PLAINKEY_39_port, 
                           PLAINKEY(38) => PLAINKEY_38_port, PLAINKEY(37) => 
                           PLAINKEY_37_port, PLAINKEY(36) => PLAINKEY_36_port, 
                           PLAINKEY(35) => PLAINKEY_35_port, PLAINKEY(34) => 
                           PLAINKEY_34_port, PLAINKEY(33) => PLAINKEY_33_port, 
                           PLAINKEY(32) => PLAINKEY_32_port, PLAINKEY(31) => 
                           PLAINKEY_31_port, PLAINKEY(30) => PLAINKEY_30_port, 
                           PLAINKEY(29) => PLAINKEY_29_port, PLAINKEY(28) => 
                           PLAINKEY_28_port, PLAINKEY(27) => PLAINKEY_27_port, 
                           PLAINKEY(26) => PLAINKEY_26_port, PLAINKEY(25) => 
                           PLAINKEY_25_port, PLAINKEY(24) => PLAINKEY_24_port, 
                           PLAINKEY(23) => PLAINKEY_23_port, PLAINKEY(22) => 
                           PLAINKEY_22_port, PLAINKEY(21) => PLAINKEY_21_port, 
                           PLAINKEY(20) => PLAINKEY_20_port, PLAINKEY(19) => 
                           PLAINKEY_19_port, PLAINKEY(18) => PLAINKEY_18_port, 
                           PLAINKEY(17) => PLAINKEY_17_port, PLAINKEY(16) => 
                           PLAINKEY_16_port, PLAINKEY(15) => PLAINKEY_15_port, 
                           PLAINKEY(14) => PLAINKEY_14_port, PLAINKEY(13) => 
                           PLAINKEY_13_port, PLAINKEY(12) => PLAINKEY_12_port, 
                           PLAINKEY(11) => PLAINKEY_11_port, PLAINKEY(10) => 
                           PLAINKEY_10_port, PLAINKEY(9) => PLAINKEY_9_port, 
                           PLAINKEY(8) => PLAINKEY_8_port, PLAINKEY(7) => 
                           PLAINKEY_7_port, PLAINKEY(6) => PLAINKEY_6_port, 
                           PLAINKEY(5) => PLAINKEY_5_port, PLAINKEY(4) => 
                           PLAINKEY_4_port, PLAINKEY(3) => PLAINKEY_3_port, 
                           PLAINKEY(2) => PLAINKEY_2_port, PLAINKEY(1) => 
                           PLAINKEY_1_port, PLAINKEY(0) => PLAINKEY_0_port, 
                           RBUF_FULL => RBUF_FULL, PARITY_ERROR => PARITY_ERROR
                           );
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity RMEDT_REWIRE_1 is

   port( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN : in std_logic;  DATA_IN : in 
         std_logic_vector (7 downto 0);  BS_ERROR, CRC_ERROR, EMPTY, FULL, 
         KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, R_ERROR, SENDING, 
         dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE : out std_logic;  DATA, 
         ADDR : out std_logic_vector (7 downto 0));

end RMEDT_REWIRE_1;

architecture SYN_struct of RMEDT_REWIRE_1 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component transmitter_block_1
      port( PRGA_OUT : in std_logic_vector (7 downto 0);  clk, p_ready : in 
            std_logic;  prga_opcode : in std_logic_vector (1 downto 0);  rst : 
            in std_logic;  SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE : out 
            std_logic);
   end component;
   
   component receiver_block_rewire_1
      port( CLK, DM1_RX, DP1_RX, RST : in std_logic;  BS_ERROR, CRC_ERROR, 
            EOP_external : out std_logic;  OPCODE : out std_logic_vector (1 
            downto 0);  RCV_DATA : out std_logic_vector (7 downto 0);  R_ERROR,
            W_ENABLE : out std_logic);
   end component;
   
   component memoryblock_1
      port( CLK, NEXT_BYTE : in std_logic;  RCV_DATA : in std_logic_vector (7 
            downto 0);  RCV_OPCODE : in std_logic_vector (1 downto 0);  RST, 
            W_ENABLE, EOP : in std_logic;  EMPTY, FULL, B_READY : out std_logic
            ;  PRGA_IN : out std_logic_vector (7 downto 0);  PRGA_OPCODE : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component EDBlock_1
      port( BYTE : in std_logic_vector (7 downto 0);  BYTE_READY, CLK : in 
            std_logic;  OPCODE : in std_logic_vector (1 downto 0);  RST, 
            SERIAL_IN : in std_logic;  DATA_IN : in std_logic_vector (7 downto 
            0);  KEY_ERROR, PARITY_ERROR, PDATA_READY : out std_logic;  
            PROCESSED_DATA : out std_logic_vector (7 downto 0);  PROG_ERROR, 
            RBUF_FULL, W_ENABLE, R_ENABLE : out std_logic;  DATA, ADDR : out 
            std_logic_vector (7 downto 0));
   end component;
   
   signal PRGA_IN_7_port, PRGA_IN_6_port, PRGA_IN_5_port, PRGA_IN_4_port, 
      PRGA_IN_3_port, PRGA_IN_2_port, PRGA_IN_1_port, PRGA_IN_0_port, B_READY, 
      PRGA_OPCODE_1_port, PRGA_OPCODE_0_port, PDATA_READY, 
      PROCESSED_DATA_7_port, PROCESSED_DATA_6_port, PROCESSED_DATA_5_port, 
      PROCESSED_DATA_4_port, PROCESSED_DATA_3_port, PROCESSED_DATA_2_port, 
      PROCESSED_DATA_1_port, PROCESSED_DATA_0_port, EOP_external, NEXT_BYTE, 
      RCV_DATA_7_port, RCV_DATA_6_port, RCV_DATA_5_port, RCV_DATA_4_port, 
      RCV_DATA_3_port, RCV_DATA_2_port, RCV_DATA_1_port, RCV_DATA_0_port, 
      OPCODE_1_port, OPCODE_0_port, W_ENABLE, n1, n2 : std_logic;

begin
   
   U_0 : EDBlock_1 port map( BYTE(7) => PRGA_IN_7_port, BYTE(6) => 
                           PRGA_IN_6_port, BYTE(5) => PRGA_IN_5_port, BYTE(4) 
                           => PRGA_IN_4_port, BYTE(3) => PRGA_IN_3_port, 
                           BYTE(2) => PRGA_IN_2_port, BYTE(1) => PRGA_IN_1_port
                           , BYTE(0) => PRGA_IN_0_port, BYTE_READY => B_READY, 
                           CLK => CLK, OPCODE(1) => PRGA_OPCODE_1_port, 
                           OPCODE(0) => PRGA_OPCODE_0_port, RST => n1, 
                           SERIAL_IN => SERIAL_IN, DATA_IN(7) => DATA_IN(7), 
                           DATA_IN(6) => DATA_IN(6), DATA_IN(5) => DATA_IN(5), 
                           DATA_IN(4) => DATA_IN(4), DATA_IN(3) => DATA_IN(3), 
                           DATA_IN(2) => DATA_IN(2), DATA_IN(1) => DATA_IN(1), 
                           DATA_IN(0) => DATA_IN(0), KEY_ERROR => KEY_ERROR, 
                           PARITY_ERROR => PARITY_ERROR, PDATA_READY => 
                           PDATA_READY, PROCESSED_DATA(7) => 
                           PROCESSED_DATA_7_port, PROCESSED_DATA(6) => 
                           PROCESSED_DATA_6_port, PROCESSED_DATA(5) => 
                           PROCESSED_DATA_5_port, PROCESSED_DATA(4) => 
                           PROCESSED_DATA_4_port, PROCESSED_DATA(3) => 
                           PROCESSED_DATA_3_port, PROCESSED_DATA(2) => 
                           PROCESSED_DATA_2_port, PROCESSED_DATA(1) => 
                           PROCESSED_DATA_1_port, PROCESSED_DATA(0) => 
                           PROCESSED_DATA_0_port, PROG_ERROR => PROG_ERROR, 
                           RBUF_FULL => RBUF_FULL, W_ENABLE => W_ENABLE_R, 
                           R_ENABLE => R_ENABLE, DATA(7) => DATA(7), DATA(6) =>
                           DATA(6), DATA(5) => DATA(5), DATA(4) => DATA(4), 
                           DATA(3) => DATA(3), DATA(2) => DATA(2), DATA(1) => 
                           DATA(1), DATA(0) => DATA(0), ADDR(7) => ADDR(7), 
                           ADDR(6) => ADDR(6), ADDR(5) => ADDR(5), ADDR(4) => 
                           ADDR(4), ADDR(3) => ADDR(3), ADDR(2) => ADDR(2), 
                           ADDR(1) => ADDR(1), ADDR(0) => ADDR(0));
   U_1 : memoryblock_1 port map( CLK => CLK, NEXT_BYTE => NEXT_BYTE, 
                           RCV_DATA(7) => RCV_DATA_7_port, RCV_DATA(6) => 
                           RCV_DATA_6_port, RCV_DATA(5) => RCV_DATA_5_port, 
                           RCV_DATA(4) => RCV_DATA_4_port, RCV_DATA(3) => 
                           RCV_DATA_3_port, RCV_DATA(2) => RCV_DATA_2_port, 
                           RCV_DATA(1) => RCV_DATA_1_port, RCV_DATA(0) => 
                           RCV_DATA_0_port, RCV_OPCODE(1) => OPCODE_1_port, 
                           RCV_OPCODE(0) => OPCODE_0_port, RST => n1, W_ENABLE 
                           => W_ENABLE, EOP => EOP_external, EMPTY => EMPTY, 
                           FULL => FULL, B_READY => B_READY, PRGA_IN(7) => 
                           PRGA_IN_7_port, PRGA_IN(6) => PRGA_IN_6_port, 
                           PRGA_IN(5) => PRGA_IN_5_port, PRGA_IN(4) => 
                           PRGA_IN_4_port, PRGA_IN(3) => PRGA_IN_3_port, 
                           PRGA_IN(2) => PRGA_IN_2_port, PRGA_IN(1) => 
                           PRGA_IN_1_port, PRGA_IN(0) => PRGA_IN_0_port, 
                           PRGA_OPCODE(1) => PRGA_OPCODE_1_port, PRGA_OPCODE(0)
                           => PRGA_OPCODE_0_port);
   U_2 : receiver_block_rewire_1 port map( CLK => CLK, DM1_RX => DM1_RX, DP1_RX
                           => DP1_RX, RST => n1, BS_ERROR => BS_ERROR, 
                           CRC_ERROR => CRC_ERROR, EOP_external => EOP_external
                           , OPCODE(1) => OPCODE_1_port, OPCODE(0) => 
                           OPCODE_0_port, RCV_DATA(7) => RCV_DATA_7_port, 
                           RCV_DATA(6) => RCV_DATA_6_port, RCV_DATA(5) => 
                           RCV_DATA_5_port, RCV_DATA(4) => RCV_DATA_4_port, 
                           RCV_DATA(3) => RCV_DATA_3_port, RCV_DATA(2) => 
                           RCV_DATA_2_port, RCV_DATA(1) => RCV_DATA_1_port, 
                           RCV_DATA(0) => RCV_DATA_0_port, R_ERROR => R_ERROR, 
                           W_ENABLE => W_ENABLE);
   U_3 : transmitter_block_1 port map( PRGA_OUT(7) => PROCESSED_DATA_7_port, 
                           PRGA_OUT(6) => PROCESSED_DATA_6_port, PRGA_OUT(5) =>
                           PROCESSED_DATA_5_port, PRGA_OUT(4) => 
                           PROCESSED_DATA_4_port, PRGA_OUT(3) => 
                           PROCESSED_DATA_3_port, PRGA_OUT(2) => 
                           PROCESSED_DATA_2_port, PRGA_OUT(1) => 
                           PROCESSED_DATA_1_port, PRGA_OUT(0) => 
                           PROCESSED_DATA_0_port, clk => CLK, p_ready => 
                           PDATA_READY, prga_opcode(1) => PRGA_OPCODE_1_port, 
                           prga_opcode(0) => PRGA_OPCODE_0_port, rst => n1, 
                           SENDING => SENDING, dm_tx_out => dm_tx_out, 
                           dp_tx_out => dp_tx_out, NEXT_BYTE => NEXT_BYTE);
   U1 : INVX2 port map( A => n2, Y => n1);
   U2 : INVX2 port map( A => RST, Y => n2);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_rmedt_square.all;

entity rmedt_square is

   port( CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN : in std_logic;  DATA_IN_H
         , DATA_IN_S : in std_logic_vector (7 downto 0);  BSE_H, BSE_S, CRCE_H,
         CRCE_S, DMTH, DMTS, DPTH, DPTS, EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H
         , RE_S, c_key_error, c_parity_error, c_prog_error, host_is_sending, 
         slave_is_sending, W_ENABLE_H, W_ENABLE_S, R_ENABLE_H, R_ENABLE_S : out
         std_logic;  DATA_H, DATA_S, ADDR_H, ADDR_S : out std_logic_vector (7 
         downto 0));

end rmedt_square;

architecture SYN_struct of rmedt_square is

   component RMEDT_REWIRE_0
      port( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN : in std_logic;  DATA_IN : in 
            std_logic_vector (7 downto 0);  BS_ERROR, CRC_ERROR, EMPTY, FULL, 
            KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, R_ERROR, SENDING, 
            dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE : out std_logic;  DATA, 
            ADDR : out std_logic_vector (7 downto 0));
   end component;
   
   component RMEDT_REWIRE_1
      port( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN : in std_logic;  DATA_IN : in 
            std_logic_vector (7 downto 0);  BS_ERROR, CRC_ERROR, EMPTY, FULL, 
            KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, R_ERROR, SENDING, 
            dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE : out std_logic;  DATA, 
            ADDR : out std_logic_vector (7 downto 0));
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal KEY_ERROR, KEY_ERROR1, PARITY_ERROR, PARITY_ERROR1, PROG_ERROR, 
      PROG_ERROR1, n_1030, n_1031 : std_logic;

begin
   
   U1 : OR2X2 port map( A => PROG_ERROR, B => PROG_ERROR1, Y => c_prog_error);
   U2 : OR2X2 port map( A => PARITY_ERROR, B => PARITY_ERROR1, Y => 
                           c_parity_error);
   U3 : OR2X2 port map( A => KEY_ERROR, B => KEY_ERROR1, Y => c_key_error);
   U_0 : RMEDT_REWIRE_1 port map( CLK => CLK, DM1_RX => DMRH, DP1_RX => DPRH, 
                           RST => RST, SERIAL_IN => SERIAL_IN, DATA_IN(7) => 
                           DATA_IN_H(7), DATA_IN(6) => DATA_IN_H(6), DATA_IN(5)
                           => DATA_IN_H(5), DATA_IN(4) => DATA_IN_H(4), 
                           DATA_IN(3) => DATA_IN_H(3), DATA_IN(2) => 
                           DATA_IN_H(2), DATA_IN(1) => DATA_IN_H(1), DATA_IN(0)
                           => DATA_IN_H(0), BS_ERROR => BSE_H, CRC_ERROR => 
                           CRCE_H, EMPTY => EMPTY_H, FULL => FULL_H, KEY_ERROR 
                           => KEY_ERROR, PROG_ERROR => PROG_ERROR, PARITY_ERROR
                           => PARITY_ERROR, RBUF_FULL => n_1030, R_ERROR => 
                           RE_H, SENDING => host_is_sending, dm_tx_out => DMTS,
                           dp_tx_out => DPTS, W_ENABLE_R => W_ENABLE_H, 
                           R_ENABLE => R_ENABLE_H, DATA(7) => DATA_H(7), 
                           DATA(6) => DATA_H(6), DATA(5) => DATA_H(5), DATA(4) 
                           => DATA_H(4), DATA(3) => DATA_H(3), DATA(2) => 
                           DATA_H(2), DATA(1) => DATA_H(1), DATA(0) => 
                           DATA_H(0), ADDR(7) => ADDR_H(7), ADDR(6) => 
                           ADDR_H(6), ADDR(5) => ADDR_H(5), ADDR(4) => 
                           ADDR_H(4), ADDR(3) => ADDR_H(3), ADDR(2) => 
                           ADDR_H(2), ADDR(1) => ADDR_H(1), ADDR(0) => 
                           ADDR_H(0));
   U_1 : RMEDT_REWIRE_0 port map( CLK => CLK, DM1_RX => DMRS, DP1_RX => DPRS, 
                           RST => RST, SERIAL_IN => SERIAL_IN, DATA_IN(7) => 
                           DATA_IN_S(7), DATA_IN(6) => DATA_IN_S(6), DATA_IN(5)
                           => DATA_IN_S(5), DATA_IN(4) => DATA_IN_S(4), 
                           DATA_IN(3) => DATA_IN_S(3), DATA_IN(2) => 
                           DATA_IN_S(2), DATA_IN(1) => DATA_IN_S(1), DATA_IN(0)
                           => DATA_IN_S(0), BS_ERROR => BSE_S, CRC_ERROR => 
                           CRCE_S, EMPTY => EMPTY_S, FULL => FULL_S, KEY_ERROR 
                           => KEY_ERROR1, PROG_ERROR => PROG_ERROR1, 
                           PARITY_ERROR => PARITY_ERROR1, RBUF_FULL => n_1031, 
                           R_ERROR => RE_S, SENDING => slave_is_sending, 
                           dm_tx_out => DMTH, dp_tx_out => DPTH, W_ENABLE_R => 
                           W_ENABLE_S, R_ENABLE => R_ENABLE_S, DATA(7) => 
                           DATA_S(7), DATA(6) => DATA_S(6), DATA(5) => 
                           DATA_S(5), DATA(4) => DATA_S(4), DATA(3) => 
                           DATA_S(3), DATA(2) => DATA_S(2), DATA(1) => 
                           DATA_S(1), DATA(0) => DATA_S(0), ADDR(7) => 
                           ADDR_S(7), ADDR(6) => ADDR_S(6), ADDR(5) => 
                           ADDR_S(5), ADDR(4) => ADDR_S(4), ADDR(3) => 
                           ADDR_S(3), ADDR(2) => ADDR_S(2), ADDR(1) => 
                           ADDR_S(1), ADDR(0) => ADDR_S(0));

end SYN_struct;
