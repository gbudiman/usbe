
module KSA_1_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_1_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_1_DW01_add_6 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;

  AND2X2 U2 ( .A(n18), .B(n14), .Y(n1) );
  NAND2X1 U3 ( .A(n33), .B(n34), .Y(n19) );
  INVX2 U4 ( .A(n38), .Y(SUM[0]) );
  XNOR2X1 U5 ( .A(n2), .B(n3), .Y(SUM[7]) );
  XOR2X1 U6 ( .A(B[7]), .B(A[7]), .Y(n3) );
  AOI21X1 U7 ( .A(n4), .B(n5), .C(n6), .Y(n2) );
  INVX2 U8 ( .A(n7), .Y(n6) );
  XNOR2X1 U9 ( .A(n4), .B(n8), .Y(SUM[6]) );
  NAND2X1 U10 ( .A(n5), .B(n7), .Y(n8) );
  NAND2X1 U11 ( .A(B[6]), .B(A[6]), .Y(n7) );
  OR2X2 U12 ( .A(A[6]), .B(B[6]), .Y(n5) );
  NAND2X1 U13 ( .A(n9), .B(n10), .Y(n4) );
  NAND2X1 U14 ( .A(n11), .B(n12), .Y(n10) );
  XNOR2X1 U15 ( .A(n11), .B(n13), .Y(SUM[5]) );
  NAND2X1 U16 ( .A(n9), .B(n12), .Y(n13) );
  OR2X2 U17 ( .A(A[5]), .B(B[5]), .Y(n12) );
  NAND2X1 U18 ( .A(B[5]), .B(A[5]), .Y(n9) );
  NAND3X1 U19 ( .A(n14), .B(n15), .C(n16), .Y(n11) );
  NAND3X1 U20 ( .A(n17), .B(n18), .C(n19), .Y(n16) );
  INVX2 U21 ( .A(n20), .Y(n17) );
  NAND3X1 U22 ( .A(n21), .B(n18), .C(n22), .Y(n15) );
  XOR2X1 U23 ( .A(n23), .B(n1), .Y(SUM[4]) );
  NAND2X1 U24 ( .A(B[4]), .B(A[4]), .Y(n14) );
  OR2X2 U25 ( .A(A[4]), .B(B[4]), .Y(n18) );
  OAI21X1 U26 ( .A(n24), .B(n20), .C(n25), .Y(n23) );
  NAND2X1 U27 ( .A(n21), .B(n22), .Y(n25) );
  NAND2X1 U28 ( .A(n26), .B(n27), .Y(n22) );
  NAND2X1 U29 ( .A(n28), .B(n21), .Y(n20) );
  INVX2 U30 ( .A(n19), .Y(n24) );
  XNOR2X1 U31 ( .A(n29), .B(n30), .Y(SUM[3]) );
  AND2X2 U32 ( .A(n21), .B(n26), .Y(n30) );
  NAND2X1 U33 ( .A(B[3]), .B(A[3]), .Y(n26) );
  OR2X2 U34 ( .A(A[3]), .B(B[3]), .Y(n21) );
  AOI21X1 U35 ( .A(n19), .B(n28), .C(n31), .Y(n29) );
  INVX2 U36 ( .A(n27), .Y(n31) );
  XNOR2X1 U37 ( .A(n32), .B(n19), .Y(SUM[2]) );
  NAND3X1 U38 ( .A(A[0]), .B(B[0]), .C(n35), .Y(n34) );
  NAND2X1 U39 ( .A(n28), .B(n27), .Y(n32) );
  NAND2X1 U40 ( .A(B[2]), .B(A[2]), .Y(n27) );
  OR2X2 U41 ( .A(A[2]), .B(B[2]), .Y(n28) );
  XOR2X1 U42 ( .A(n36), .B(n37), .Y(SUM[1]) );
  NAND2X1 U43 ( .A(n35), .B(n33), .Y(n36) );
  NAND2X1 U44 ( .A(B[1]), .B(A[1]), .Y(n33) );
  OR2X2 U45 ( .A(A[1]), .B(B[1]), .Y(n35) );
  OAI21X1 U46 ( .A(A[0]), .B(B[0]), .C(n37), .Y(n38) );
  NAND2X1 U47 ( .A(B[0]), .B(A[0]), .Y(n37) );
endmodule


module KSA_1_DW01_add_7 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  NAND2X1 U2 ( .A(n35), .B(n36), .Y(n30) );
  INVX2 U3 ( .A(n40), .Y(SUM[0]) );
  XNOR2X1 U4 ( .A(n1), .B(n2), .Y(SUM[7]) );
  XOR2X1 U5 ( .A(B[7]), .B(A[7]), .Y(n2) );
  AOI21X1 U6 ( .A(n3), .B(n4), .C(n5), .Y(n1) );
  INVX2 U7 ( .A(n6), .Y(n5) );
  XNOR2X1 U8 ( .A(n3), .B(n7), .Y(SUM[6]) );
  NAND2X1 U9 ( .A(n4), .B(n6), .Y(n7) );
  NAND2X1 U10 ( .A(B[6]), .B(A[6]), .Y(n6) );
  OR2X2 U11 ( .A(A[6]), .B(B[6]), .Y(n4) );
  NAND2X1 U12 ( .A(n8), .B(n9), .Y(n3) );
  NAND2X1 U13 ( .A(n10), .B(n11), .Y(n9) );
  XNOR2X1 U14 ( .A(n10), .B(n12), .Y(SUM[5]) );
  NAND2X1 U15 ( .A(n8), .B(n11), .Y(n12) );
  OR2X2 U16 ( .A(A[5]), .B(B[5]), .Y(n11) );
  NAND2X1 U17 ( .A(B[5]), .B(A[5]), .Y(n8) );
  OAI21X1 U18 ( .A(n13), .B(n14), .C(n15), .Y(n10) );
  AOI21X1 U19 ( .A(n16), .B(n17), .C(n18), .Y(n15) );
  INVX2 U20 ( .A(n19), .Y(n18) );
  INVX2 U21 ( .A(n20), .Y(n16) );
  NAND2X1 U22 ( .A(n21), .B(n17), .Y(n14) );
  INVX2 U23 ( .A(n22), .Y(n21) );
  XNOR2X1 U24 ( .A(n23), .B(n24), .Y(SUM[4]) );
  OAI21X1 U25 ( .A(n13), .B(n22), .C(n20), .Y(n24) );
  OAI21X1 U26 ( .A(n25), .B(n26), .C(n27), .Y(n20) );
  INVX2 U27 ( .A(n28), .Y(n26) );
  NAND2X1 U28 ( .A(n29), .B(n27), .Y(n22) );
  INVX2 U29 ( .A(n30), .Y(n13) );
  NAND2X1 U30 ( .A(n17), .B(n19), .Y(n23) );
  NAND2X1 U31 ( .A(B[4]), .B(A[4]), .Y(n19) );
  OR2X2 U32 ( .A(A[4]), .B(B[4]), .Y(n17) );
  XNOR2X1 U33 ( .A(n31), .B(n32), .Y(SUM[3]) );
  AND2X2 U34 ( .A(n27), .B(n28), .Y(n32) );
  NAND2X1 U35 ( .A(B[3]), .B(A[3]), .Y(n28) );
  OR2X2 U36 ( .A(A[3]), .B(B[3]), .Y(n27) );
  AOI21X1 U37 ( .A(n30), .B(n29), .C(n25), .Y(n31) );
  INVX2 U38 ( .A(n33), .Y(n25) );
  XNOR2X1 U39 ( .A(n34), .B(n30), .Y(SUM[2]) );
  NAND3X1 U40 ( .A(A[0]), .B(B[0]), .C(n37), .Y(n36) );
  NAND2X1 U41 ( .A(n29), .B(n33), .Y(n34) );
  NAND2X1 U42 ( .A(B[2]), .B(A[2]), .Y(n33) );
  OR2X2 U43 ( .A(A[2]), .B(B[2]), .Y(n29) );
  XOR2X1 U44 ( .A(n38), .B(n39), .Y(SUM[1]) );
  NAND2X1 U45 ( .A(n37), .B(n35), .Y(n38) );
  NAND2X1 U46 ( .A(B[1]), .B(A[1]), .Y(n35) );
  OR2X2 U47 ( .A(A[1]), .B(B[1]), .Y(n37) );
  OAI21X1 U48 ( .A(A[0]), .B(B[0]), .C(n39), .Y(n40) );
  NAND2X1 U49 ( .A(B[0]), .B(A[0]), .Y(n39) );
endmodule


module KSA_1_DW01_add_8 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49;

  BUFX2 U2 ( .A(n6), .Y(n1) );
  XNOR2X1 U3 ( .A(n6), .B(n10), .Y(SUM[6]) );
  XNOR2X1 U4 ( .A(n27), .B(n2), .Y(SUM[4]) );
  NAND2X1 U5 ( .A(n21), .B(n23), .Y(n2) );
  XOR2X1 U6 ( .A(n48), .B(n47), .Y(SUM[1]) );
  XOR2X1 U7 ( .A(n35), .B(n36), .Y(SUM[3]) );
  AND2X2 U8 ( .A(n33), .B(n31), .Y(n3) );
  INVX2 U9 ( .A(n39), .Y(n38) );
  NAND2X1 U10 ( .A(n45), .B(n42), .Y(n43) );
  INVX2 U11 ( .A(n49), .Y(SUM[0]) );
  XNOR2X1 U12 ( .A(n4), .B(n5), .Y(SUM[7]) );
  XOR2X1 U13 ( .A(B[7]), .B(A[7]), .Y(n5) );
  AOI21X1 U14 ( .A(n1), .B(n7), .C(n8), .Y(n4) );
  INVX2 U15 ( .A(n9), .Y(n8) );
  NAND2X1 U16 ( .A(n7), .B(n9), .Y(n10) );
  NAND2X1 U17 ( .A(B[6]), .B(A[6]), .Y(n9) );
  OR2X2 U18 ( .A(A[6]), .B(B[6]), .Y(n7) );
  OAI21X1 U19 ( .A(n11), .B(n12), .C(n13), .Y(n6) );
  INVX2 U20 ( .A(n14), .Y(n12) );
  INVX2 U21 ( .A(n15), .Y(n11) );
  XNOR2X1 U22 ( .A(n14), .B(n16), .Y(SUM[5]) );
  OAI21X1 U23 ( .A(n17), .B(n18), .C(n19), .Y(n14) );
  AOI21X1 U24 ( .A(n20), .B(n21), .C(n22), .Y(n19) );
  INVX2 U25 ( .A(n23), .Y(n22) );
  NAND2X1 U26 ( .A(n24), .B(n25), .Y(n20) );
  NAND3X1 U27 ( .A(n26), .B(n21), .C(n3), .Y(n18) );
  NAND2X1 U28 ( .A(n13), .B(n15), .Y(n16) );
  OR2X2 U29 ( .A(A[5]), .B(B[5]), .Y(n15) );
  NAND2X1 U30 ( .A(B[5]), .B(A[5]), .Y(n13) );
  NAND2X1 U31 ( .A(B[4]), .B(A[4]), .Y(n23) );
  OR2X2 U32 ( .A(A[4]), .B(B[4]), .Y(n21) );
  OAI21X1 U33 ( .A(n17), .B(n28), .C(n29), .Y(n27) );
  AND2X2 U34 ( .A(n24), .B(n25), .Y(n29) );
  NAND2X1 U35 ( .A(n30), .B(n31), .Y(n24) );
  INVX2 U36 ( .A(n32), .Y(n30) );
  NAND2X1 U37 ( .A(n3), .B(n26), .Y(n28) );
  AOI21X1 U38 ( .A(B[0]), .B(A[0]), .C(n34), .Y(n17) );
  NAND2X1 U39 ( .A(n25), .B(n31), .Y(n36) );
  OR2X2 U40 ( .A(A[3]), .B(B[3]), .Y(n31) );
  NAND2X1 U41 ( .A(B[3]), .B(A[3]), .Y(n25) );
  NOR2X1 U42 ( .A(n37), .B(n38), .Y(n35) );
  NAND3X1 U43 ( .A(n26), .B(n33), .C(n40), .Y(n39) );
  AND2X2 U44 ( .A(B[0]), .B(A[0]), .Y(n40) );
  NAND2X1 U45 ( .A(n41), .B(n32), .Y(n37) );
  NAND2X1 U46 ( .A(n34), .B(n33), .Y(n41) );
  INVX2 U47 ( .A(n42), .Y(n34) );
  XNOR2X1 U48 ( .A(n43), .B(n44), .Y(SUM[2]) );
  NAND2X1 U49 ( .A(n33), .B(n32), .Y(n44) );
  NAND2X1 U50 ( .A(B[2]), .B(A[2]), .Y(n32) );
  OR2X2 U51 ( .A(A[2]), .B(B[2]), .Y(n33) );
  NAND2X1 U52 ( .A(n46), .B(n26), .Y(n45) );
  AND2X2 U53 ( .A(A[0]), .B(B[0]), .Y(n46) );
  NAND2X1 U54 ( .A(n42), .B(n26), .Y(n47) );
  OR2X2 U55 ( .A(A[1]), .B(B[1]), .Y(n26) );
  NAND2X1 U56 ( .A(B[1]), .B(A[1]), .Y(n42) );
  OAI21X1 U57 ( .A(A[0]), .B(B[0]), .C(n48), .Y(n49) );
  NAND2X1 U58 ( .A(B[0]), .B(A[0]), .Y(n48) );
endmodule


module KSA_1_DW01_add_9 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;

  NAND2X1 U2 ( .A(n5), .B(n39), .Y(n1) );
  NAND2X1 U3 ( .A(n5), .B(n39), .Y(n2) );
  INVX1 U4 ( .A(n19), .Y(n3) );
  INVX1 U5 ( .A(B[6]), .Y(n19) );
  INVX1 U6 ( .A(n7), .Y(n23) );
  AND2X2 U7 ( .A(n29), .B(n13), .Y(n4) );
  NAND2X1 U8 ( .A(n5), .B(n39), .Y(n17) );
  AND2X2 U9 ( .A(n40), .B(n41), .Y(n5) );
  AND2X2 U10 ( .A(B[0]), .B(A[0]), .Y(n6) );
  OAI21X1 U11 ( .A(B[6]), .B(A[6]), .C(n13), .Y(n7) );
  OR2X2 U12 ( .A(B[6]), .B(A[6]), .Y(n14) );
  INVX2 U13 ( .A(n39), .Y(n36) );
  INVX2 U14 ( .A(n61), .Y(SUM[0]) );
  XOR2X1 U15 ( .A(n8), .B(n9), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(B[7]), .B(A[7]), .Y(n9) );
  NAND3X1 U17 ( .A(n10), .B(n11), .C(n12), .Y(n8) );
  NAND3X1 U18 ( .A(n13), .B(n14), .C(n15), .Y(n12) );
  NAND3X1 U19 ( .A(n16), .B(n13), .C(n17), .Y(n11) );
  AOI21X1 U20 ( .A(n18), .B(n19), .C(n20), .Y(n16) );
  NAND2X1 U21 ( .A(n21), .B(n22), .Y(n20) );
  INVX2 U22 ( .A(A[6]), .Y(n18) );
  AOI21X1 U23 ( .A(n23), .B(n24), .C(n25), .Y(n10) );
  NAND2X1 U24 ( .A(n26), .B(n27), .Y(n25) );
  OAI21X1 U25 ( .A(A[6]), .B(B[6]), .C(n28), .Y(n27) );
  INVX2 U26 ( .A(n29), .Y(n28) );
  XOR2X1 U27 ( .A(n30), .B(n31), .Y(SUM[6]) );
  INVX2 U28 ( .A(n32), .Y(n31) );
  OAI21X1 U29 ( .A(n3), .B(A[6]), .C(n26), .Y(n32) );
  NAND2X1 U30 ( .A(B[6]), .B(A[6]), .Y(n26) );
  NAND3X1 U31 ( .A(n29), .B(n33), .C(n34), .Y(n30) );
  OAI21X1 U32 ( .A(n35), .B(n36), .C(n37), .Y(n34) );
  AND2X2 U33 ( .A(n38), .B(n13), .Y(n37) );
  NAND2X1 U34 ( .A(n40), .B(n41), .Y(n35) );
  AOI22X1 U35 ( .A(n24), .B(n13), .C(n15), .D(n13), .Y(n33) );
  INVX2 U36 ( .A(n42), .Y(n15) );
  INVX2 U37 ( .A(n43), .Y(n24) );
  XNOR2X1 U38 ( .A(n44), .B(n4), .Y(SUM[5]) );
  OR2X2 U39 ( .A(A[5]), .B(B[5]), .Y(n13) );
  NAND2X1 U40 ( .A(B[5]), .B(A[5]), .Y(n29) );
  AOI21X1 U41 ( .A(n38), .B(n1), .C(n45), .Y(n44) );
  NAND2X1 U42 ( .A(n42), .B(n43), .Y(n45) );
  NAND3X1 U43 ( .A(A[3]), .B(B[3]), .C(n21), .Y(n42) );
  INVX2 U44 ( .A(n46), .Y(n38) );
  OAI21X1 U45 ( .A(A[4]), .B(B[4]), .C(n22), .Y(n46) );
  XNOR2X1 U46 ( .A(n47), .B(n48), .Y(SUM[4]) );
  AND2X2 U47 ( .A(n21), .B(n43), .Y(n48) );
  NAND2X1 U48 ( .A(B[4]), .B(A[4]), .Y(n43) );
  OR2X2 U49 ( .A(A[4]), .B(B[4]), .Y(n21) );
  AOI21X1 U50 ( .A(n2), .B(n22), .C(n49), .Y(n47) );
  INVX2 U51 ( .A(n50), .Y(n49) );
  XNOR2X1 U52 ( .A(n17), .B(n51), .Y(SUM[3]) );
  NAND2X1 U53 ( .A(n22), .B(n50), .Y(n51) );
  NAND2X1 U54 ( .A(B[3]), .B(A[3]), .Y(n50) );
  OR2X2 U55 ( .A(A[3]), .B(B[3]), .Y(n22) );
  NAND3X1 U56 ( .A(n52), .B(n53), .C(n54), .Y(n39) );
  AND2X2 U57 ( .A(B[0]), .B(A[0]), .Y(n54) );
  NAND3X1 U58 ( .A(A[1]), .B(B[1]), .C(n53), .Y(n40) );
  XOR2X1 U59 ( .A(n55), .B(n56), .Y(SUM[2]) );
  AOI21X1 U60 ( .A(n6), .B(n52), .C(n57), .Y(n56) );
  INVX2 U61 ( .A(n58), .Y(n57) );
  NAND2X1 U62 ( .A(n53), .B(n41), .Y(n55) );
  NAND2X1 U63 ( .A(B[2]), .B(A[2]), .Y(n41) );
  OR2X2 U64 ( .A(A[2]), .B(B[2]), .Y(n53) );
  XNOR2X1 U65 ( .A(n59), .B(n6), .Y(SUM[1]) );
  NAND2X1 U66 ( .A(n52), .B(n58), .Y(n59) );
  NAND2X1 U67 ( .A(B[1]), .B(A[1]), .Y(n58) );
  OR2X2 U68 ( .A(A[1]), .B(B[1]), .Y(n52) );
  OAI21X1 U69 ( .A(A[0]), .B(B[0]), .C(n60), .Y(n61) );
  NAND2X1 U70 ( .A(B[0]), .B(A[0]), .Y(n60) );
endmodule


module KSA_1_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  XOR2X1 U2 ( .A(n5), .B(A[4]), .Y(SUM[4]) );
  XOR2X1 U3 ( .A(n1), .B(A[2]), .Y(SUM[2]) );
  XOR2X1 U4 ( .A(n3), .B(A[6]), .Y(SUM[6]) );
  AND2X2 U5 ( .A(A[1]), .B(A[0]), .Y(n1) );
  XNOR2X1 U6 ( .A(A[7]), .B(n2), .Y(SUM[7]) );
  NAND2X1 U7 ( .A(A[6]), .B(n3), .Y(n2) );
  INVX2 U8 ( .A(n4), .Y(n3) );
  NAND3X1 U9 ( .A(A[4]), .B(A[5]), .C(n5), .Y(n4) );
  XNOR2X1 U10 ( .A(A[5]), .B(n6), .Y(SUM[5]) );
  NAND2X1 U11 ( .A(A[4]), .B(n5), .Y(n6) );
  INVX2 U12 ( .A(n7), .Y(n5) );
  NAND3X1 U13 ( .A(A[2]), .B(A[3]), .C(n1), .Y(n7) );
  XNOR2X1 U14 ( .A(A[3]), .B(n8), .Y(SUM[3]) );
  NAND2X1 U15 ( .A(A[2]), .B(n1), .Y(n8) );
  XOR2X1 U16 ( .A(A[1]), .B(A[0]), .Y(SUM[1]) );
  INVX2 U17 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module KSA_1 ( KEY, CLK, RST, KEY_ERROR, BYTE_READY, BYTE, OPCODE, DATA_IN, 
        PROCESSED_DATA, PDATA_READY, W_ENABLE, R_ENABLE, ADDR, DATA );
  input [63:0] KEY;
  input [7:0] BYTE;
  input [1:0] OPCODE;
  input [7:0] DATA_IN;
  output [7:0] PROCESSED_DATA;
  output [7:0] ADDR;
  output [7:0] DATA;
  input CLK, RST, KEY_ERROR, BYTE_READY;
  output PDATA_READY, W_ENABLE, R_ENABLE;
  wire   permuteComplete, \keyTable[0][7] , \keyTable[0][6] , \keyTable[0][5] ,
         \keyTable[0][4] , \keyTable[0][3] , \keyTable[0][2] ,
         \keyTable[0][1] , \keyTable[0][0] , \keyTable[1][7] ,
         \keyTable[1][6] , \keyTable[1][5] , \keyTable[1][4] ,
         \keyTable[1][3] , \keyTable[1][2] , \keyTable[1][1] ,
         \keyTable[1][0] , \keyTable[2][7] , \keyTable[2][6] ,
         \keyTable[2][5] , \keyTable[2][4] , \keyTable[2][3] ,
         \keyTable[2][2] , \keyTable[2][1] , \keyTable[2][0] ,
         \keyTable[3][7] , \keyTable[3][6] , \keyTable[3][5] ,
         \keyTable[3][4] , \keyTable[3][3] , \keyTable[3][2] ,
         \keyTable[3][1] , \keyTable[3][0] , \keyTable[4][7] ,
         \keyTable[4][6] , \keyTable[4][5] , \keyTable[4][4] ,
         \keyTable[4][3] , \keyTable[4][2] , \keyTable[4][1] ,
         \keyTable[4][0] , \keyTable[5][7] , \keyTable[5][6] ,
         \keyTable[5][5] , \keyTable[5][4] , \keyTable[5][3] ,
         \keyTable[5][2] , \keyTable[5][1] , \keyTable[5][0] ,
         \keyTable[6][7] , \keyTable[6][6] , \keyTable[6][5] ,
         \keyTable[6][4] , \keyTable[6][3] , \keyTable[6][2] ,
         \keyTable[6][1] , \keyTable[6][0] , \keyTable[7][7] ,
         \keyTable[7][6] , \keyTable[7][5] , \keyTable[7][4] ,
         \keyTable[7][3] , \keyTable[7][2] , \keyTable[7][1] ,
         \keyTable[7][0] , fw_enable, fr_enable, N407, N408, N409, N410, N411,
         N412, N413, N414, N424, N425, N426, N427, N428, N429, N430, N431,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N496, N497, N498, N499, N500, N501,
         N502, N503, N512, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N522, N523, N524, N525, N526, N527, n124, n126, n128, n130,
         n155, n158, n159, n163, n165, n168, n173, n174, n176, n186, n204,
         n588, n589, n691, n693, n694, n695, n696, n697, n698, n699, n700,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n747, n749, n751, n753, n755, n757, n759, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n891, n892, n893, n894, n895, n896, n897, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, N456, N455, N454, N453, N452, N451, N450,
         N449, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n125, n127,
         n129, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n156, n157, n160, n161, n162, n164, n166, n167,
         n169, n170, n171, n172, n175, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n692, n701,
         n765, n766, n769, n770, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n864, n865, n866, n867, n868, n869, n870, n871, n883,
         n884, n885, n886, n887, n888, n889, n890, n898, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136;
  wire   [4:0] state;
  wire   [7:0] si;
  wire   [7:0] sj;
  wire   [7:0] currentProcessedData;
  wire   [4:0] nextState;
  wire   [7:0] inti;
  wire   [7:0] intj;
  wire   [2:0] keyi;
  wire   [7:0] temp;
  wire   [7:0] extratemp;
  wire   [7:0] nextProcessedData;
  wire   [7:0] delaydata;
  wire   [7:0] prefillCounter;
  wire   [7:0] faddr;
  wire   [7:0] fdata;
  tri   [7:0] nfaddr;
  tri   [7:0] nfdata;

  DFFPOSX1 \prefillCounter_reg[0]  ( .D(n915), .CLK(CLK), .Q(prefillCounter[0]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n212), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n212), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[4]  ( .D(nextState[4]), .CLK(CLK), .R(n211), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n211), .S(1'b1), .Q(
        state[0]) );
  DFFPOSX1 permuteComplete_reg ( .D(n899), .CLK(CLK), .Q(permuteComplete) );
  DFFSR \state_reg[3]  ( .D(nextState[3]), .CLK(CLK), .R(n211), .S(1'b1), .Q(
        state[3]) );
  DFFSR PDATA_READY_reg ( .D(n1135), .CLK(CLK), .R(n211), .S(1'b1), .Q(
        PDATA_READY) );
  DFFPOSX1 \extratemp_reg[7]  ( .D(n1134), .CLK(CLK), .Q(extratemp[7]) );
  DFFPOSX1 \extratemp_reg[6]  ( .D(n1133), .CLK(CLK), .Q(extratemp[6]) );
  DFFPOSX1 \extratemp_reg[5]  ( .D(n1132), .CLK(CLK), .Q(extratemp[5]) );
  DFFPOSX1 \extratemp_reg[4]  ( .D(n1131), .CLK(CLK), .Q(extratemp[4]) );
  DFFPOSX1 \extratemp_reg[3]  ( .D(n1130), .CLK(CLK), .Q(extratemp[3]) );
  DFFPOSX1 \extratemp_reg[2]  ( .D(n1129), .CLK(CLK), .Q(extratemp[2]) );
  DFFPOSX1 \extratemp_reg[1]  ( .D(n1128), .CLK(CLK), .Q(extratemp[1]) );
  DFFPOSX1 \extratemp_reg[0]  ( .D(n1127), .CLK(CLK), .Q(extratemp[0]) );
  DFFPOSX1 \keyTable_reg[7][0]  ( .D(n792), .CLK(CLK), .Q(\keyTable[7][0] ) );
  DFFPOSX1 \keyTable_reg[7][1]  ( .D(n793), .CLK(CLK), .Q(\keyTable[7][1] ) );
  DFFPOSX1 \keyTable_reg[7][2]  ( .D(n794), .CLK(CLK), .Q(\keyTable[7][2] ) );
  DFFPOSX1 \keyTable_reg[7][3]  ( .D(n795), .CLK(CLK), .Q(\keyTable[7][3] ) );
  DFFPOSX1 \keyTable_reg[7][4]  ( .D(n796), .CLK(CLK), .Q(\keyTable[7][4] ) );
  DFFPOSX1 \keyTable_reg[7][5]  ( .D(n797), .CLK(CLK), .Q(\keyTable[7][5] ) );
  DFFPOSX1 \keyTable_reg[7][6]  ( .D(n798), .CLK(CLK), .Q(\keyTable[7][6] ) );
  DFFPOSX1 \keyTable_reg[7][7]  ( .D(n799), .CLK(CLK), .Q(\keyTable[7][7] ) );
  DFFPOSX1 \keyTable_reg[6][0]  ( .D(n800), .CLK(CLK), .Q(\keyTable[6][0] ) );
  DFFPOSX1 \keyTable_reg[6][1]  ( .D(n801), .CLK(CLK), .Q(\keyTable[6][1] ) );
  DFFPOSX1 \keyTable_reg[6][2]  ( .D(n802), .CLK(CLK), .Q(\keyTable[6][2] ) );
  DFFPOSX1 \keyTable_reg[6][3]  ( .D(n803), .CLK(CLK), .Q(\keyTable[6][3] ) );
  DFFPOSX1 \keyTable_reg[6][4]  ( .D(n804), .CLK(CLK), .Q(\keyTable[6][4] ) );
  DFFPOSX1 \keyTable_reg[6][5]  ( .D(n805), .CLK(CLK), .Q(\keyTable[6][5] ) );
  DFFPOSX1 \keyTable_reg[6][6]  ( .D(n806), .CLK(CLK), .Q(\keyTable[6][6] ) );
  DFFPOSX1 \keyTable_reg[6][7]  ( .D(n807), .CLK(CLK), .Q(\keyTable[6][7] ) );
  DFFPOSX1 \keyTable_reg[5][0]  ( .D(n808), .CLK(CLK), .Q(\keyTable[5][0] ) );
  DFFPOSX1 \keyTable_reg[5][1]  ( .D(n809), .CLK(CLK), .Q(\keyTable[5][1] ) );
  DFFPOSX1 \keyTable_reg[5][2]  ( .D(n810), .CLK(CLK), .Q(\keyTable[5][2] ) );
  DFFPOSX1 \keyTable_reg[5][3]  ( .D(n811), .CLK(CLK), .Q(\keyTable[5][3] ) );
  DFFPOSX1 \keyTable_reg[5][4]  ( .D(n812), .CLK(CLK), .Q(\keyTable[5][4] ) );
  DFFPOSX1 \keyTable_reg[5][5]  ( .D(n813), .CLK(CLK), .Q(\keyTable[5][5] ) );
  DFFPOSX1 \keyTable_reg[5][6]  ( .D(n814), .CLK(CLK), .Q(\keyTable[5][6] ) );
  DFFPOSX1 \keyTable_reg[5][7]  ( .D(n815), .CLK(CLK), .Q(\keyTable[5][7] ) );
  DFFPOSX1 \keyTable_reg[4][0]  ( .D(n816), .CLK(CLK), .Q(\keyTable[4][0] ) );
  DFFPOSX1 \keyTable_reg[4][1]  ( .D(n817), .CLK(CLK), .Q(\keyTable[4][1] ) );
  DFFPOSX1 \keyTable_reg[4][2]  ( .D(n818), .CLK(CLK), .Q(\keyTable[4][2] ) );
  DFFPOSX1 \keyTable_reg[4][3]  ( .D(n819), .CLK(CLK), .Q(\keyTable[4][3] ) );
  DFFPOSX1 \keyTable_reg[4][4]  ( .D(n820), .CLK(CLK), .Q(\keyTable[4][4] ) );
  DFFPOSX1 \keyTable_reg[4][5]  ( .D(n821), .CLK(CLK), .Q(\keyTable[4][5] ) );
  DFFPOSX1 \keyTable_reg[4][6]  ( .D(n822), .CLK(CLK), .Q(\keyTable[4][6] ) );
  DFFPOSX1 \keyTable_reg[4][7]  ( .D(n823), .CLK(CLK), .Q(\keyTable[4][7] ) );
  DFFPOSX1 \keyTable_reg[3][0]  ( .D(n824), .CLK(CLK), .Q(\keyTable[3][0] ) );
  DFFPOSX1 \keyTable_reg[3][1]  ( .D(n825), .CLK(CLK), .Q(\keyTable[3][1] ) );
  DFFPOSX1 \keyTable_reg[3][2]  ( .D(n826), .CLK(CLK), .Q(\keyTable[3][2] ) );
  DFFPOSX1 \keyTable_reg[3][3]  ( .D(n827), .CLK(CLK), .Q(\keyTable[3][3] ) );
  DFFPOSX1 \keyTable_reg[3][4]  ( .D(n828), .CLK(CLK), .Q(\keyTable[3][4] ) );
  DFFPOSX1 \keyTable_reg[3][5]  ( .D(n829), .CLK(CLK), .Q(\keyTable[3][5] ) );
  DFFPOSX1 \keyTable_reg[3][6]  ( .D(n830), .CLK(CLK), .Q(\keyTable[3][6] ) );
  DFFPOSX1 \keyTable_reg[3][7]  ( .D(n831), .CLK(CLK), .Q(\keyTable[3][7] ) );
  DFFPOSX1 \keyTable_reg[2][0]  ( .D(n832), .CLK(CLK), .Q(\keyTable[2][0] ) );
  DFFPOSX1 \keyTable_reg[2][1]  ( .D(n833), .CLK(CLK), .Q(\keyTable[2][1] ) );
  DFFPOSX1 \keyTable_reg[2][2]  ( .D(n834), .CLK(CLK), .Q(\keyTable[2][2] ) );
  DFFPOSX1 \keyTable_reg[2][3]  ( .D(n835), .CLK(CLK), .Q(\keyTable[2][3] ) );
  DFFPOSX1 \keyTable_reg[2][4]  ( .D(n836), .CLK(CLK), .Q(\keyTable[2][4] ) );
  DFFPOSX1 \keyTable_reg[2][5]  ( .D(n837), .CLK(CLK), .Q(\keyTable[2][5] ) );
  DFFPOSX1 \keyTable_reg[2][6]  ( .D(n838), .CLK(CLK), .Q(\keyTable[2][6] ) );
  DFFPOSX1 \keyTable_reg[2][7]  ( .D(n839), .CLK(CLK), .Q(\keyTable[2][7] ) );
  DFFPOSX1 \keyTable_reg[1][0]  ( .D(n840), .CLK(CLK), .Q(\keyTable[1][0] ) );
  DFFPOSX1 \keyTable_reg[1][1]  ( .D(n841), .CLK(CLK), .Q(\keyTable[1][1] ) );
  DFFPOSX1 \keyTable_reg[1][2]  ( .D(n842), .CLK(CLK), .Q(\keyTable[1][2] ) );
  DFFPOSX1 \keyTable_reg[1][3]  ( .D(n843), .CLK(CLK), .Q(\keyTable[1][3] ) );
  DFFPOSX1 \keyTable_reg[1][4]  ( .D(n844), .CLK(CLK), .Q(\keyTable[1][4] ) );
  DFFPOSX1 \keyTable_reg[1][5]  ( .D(n845), .CLK(CLK), .Q(\keyTable[1][5] ) );
  DFFPOSX1 \keyTable_reg[1][6]  ( .D(n846), .CLK(CLK), .Q(\keyTable[1][6] ) );
  DFFPOSX1 \keyTable_reg[0][6]  ( .D(n847), .CLK(CLK), .Q(\keyTable[0][6] ) );
  DFFPOSX1 \keyTable_reg[0][5]  ( .D(n848), .CLK(CLK), .Q(\keyTable[0][5] ) );
  DFFPOSX1 \keyTable_reg[0][4]  ( .D(n849), .CLK(CLK), .Q(\keyTable[0][4] ) );
  DFFPOSX1 \keyTable_reg[0][3]  ( .D(n850), .CLK(CLK), .Q(\keyTable[0][3] ) );
  DFFPOSX1 \keyTable_reg[0][2]  ( .D(n851), .CLK(CLK), .Q(\keyTable[0][2] ) );
  DFFPOSX1 \keyTable_reg[0][1]  ( .D(n852), .CLK(CLK), .Q(\keyTable[0][1] ) );
  DFFPOSX1 \keyTable_reg[0][0]  ( .D(n853), .CLK(CLK), .Q(\keyTable[0][0] ) );
  DFFPOSX1 \keyTable_reg[1][7]  ( .D(n854), .CLK(CLK), .Q(\keyTable[1][7] ) );
  DFFPOSX1 \keyTable_reg[0][7]  ( .D(n855), .CLK(CLK), .Q(\keyTable[0][7] ) );
  DFFPOSX1 \prefillCounter_reg[7]  ( .D(n914), .CLK(CLK), .Q(prefillCounter[7]) );
  DFFPOSX1 \prefillCounter_reg[1]  ( .D(n913), .CLK(CLK), .Q(prefillCounter[1]) );
  DFFPOSX1 \prefillCounter_reg[2]  ( .D(n912), .CLK(CLK), .Q(prefillCounter[2]) );
  DFFPOSX1 \prefillCounter_reg[3]  ( .D(n911), .CLK(CLK), .Q(prefillCounter[3]) );
  DFFPOSX1 \prefillCounter_reg[4]  ( .D(n910), .CLK(CLK), .Q(prefillCounter[4]) );
  DFFPOSX1 \prefillCounter_reg[5]  ( .D(n909), .CLK(CLK), .Q(prefillCounter[5]) );
  DFFPOSX1 \prefillCounter_reg[6]  ( .D(n908), .CLK(CLK), .Q(prefillCounter[6]) );
  DFFPOSX1 \temp_reg[7]  ( .D(n856), .CLK(CLK), .Q(temp[7]) );
  DFFPOSX1 \temp_reg[0]  ( .D(n863), .CLK(CLK), .Q(temp[0]) );
  DFFPOSX1 \temp_reg[1]  ( .D(n862), .CLK(CLK), .Q(temp[1]) );
  DFFPOSX1 \temp_reg[2]  ( .D(n861), .CLK(CLK), .Q(temp[2]) );
  DFFPOSX1 \temp_reg[3]  ( .D(n860), .CLK(CLK), .Q(temp[3]) );
  DFFPOSX1 \temp_reg[4]  ( .D(n859), .CLK(CLK), .Q(temp[4]) );
  DFFPOSX1 \temp_reg[5]  ( .D(n858), .CLK(CLK), .Q(temp[5]) );
  DFFPOSX1 \temp_reg[6]  ( .D(n857), .CLK(CLK), .Q(temp[6]) );
  DFFSR \si_reg[0]  ( .D(n907), .CLK(CLK), .R(n211), .S(1'b1), .Q(si[0]) );
  DFFSR \si_reg[1]  ( .D(n906), .CLK(CLK), .R(n210), .S(1'b1), .Q(si[1]) );
  DFFSR \si_reg[2]  ( .D(n905), .CLK(CLK), .R(n210), .S(1'b1), .Q(si[2]) );
  DFFSR \si_reg[3]  ( .D(n904), .CLK(CLK), .R(n210), .S(1'b1), .Q(si[3]) );
  DFFSR \si_reg[4]  ( .D(n903), .CLK(CLK), .R(n209), .S(1'b1), .Q(si[4]) );
  DFFSR \si_reg[5]  ( .D(n902), .CLK(CLK), .R(n210), .S(1'b1), .Q(si[5]) );
  DFFPOSX1 \delaydata_reg[7]  ( .D(n1111), .CLK(CLK), .Q(delaydata[7]) );
  DFFPOSX1 \delaydata_reg[0]  ( .D(n1118), .CLK(CLK), .Q(delaydata[0]) );
  DFFPOSX1 \delaydata_reg[1]  ( .D(n1117), .CLK(CLK), .Q(delaydata[1]) );
  DFFPOSX1 \delaydata_reg[2]  ( .D(n1116), .CLK(CLK), .Q(delaydata[2]) );
  DFFPOSX1 \delaydata_reg[3]  ( .D(n1115), .CLK(CLK), .Q(delaydata[3]) );
  DFFPOSX1 \delaydata_reg[4]  ( .D(n1114), .CLK(CLK), .Q(delaydata[4]) );
  DFFPOSX1 \delaydata_reg[5]  ( .D(n1113), .CLK(CLK), .Q(delaydata[5]) );
  DFFPOSX1 \delaydata_reg[6]  ( .D(n1112), .CLK(CLK), .Q(delaydata[6]) );
  DFFPOSX1 \intj_reg[7]  ( .D(n875), .CLK(CLK), .Q(intj[7]) );
  DFFPOSX1 \intj_reg[0]  ( .D(n882), .CLK(CLK), .Q(intj[0]) );
  DFFPOSX1 \intj_reg[1]  ( .D(n881), .CLK(CLK), .Q(intj[1]) );
  DFFPOSX1 \intj_reg[2]  ( .D(n880), .CLK(CLK), .Q(intj[2]) );
  DFFPOSX1 \intj_reg[3]  ( .D(n879), .CLK(CLK), .Q(intj[3]) );
  DFFPOSX1 \intj_reg[4]  ( .D(n878), .CLK(CLK), .Q(intj[4]) );
  DFFPOSX1 \intj_reg[5]  ( .D(n877), .CLK(CLK), .Q(intj[5]) );
  DFFPOSX1 \intj_reg[6]  ( .D(n876), .CLK(CLK), .Q(intj[6]) );
  DFFSR \sj_reg[7]  ( .D(n1099), .CLK(CLK), .R(n209), .S(1'b1), .Q(sj[7]) );
  DFFSR \sj_reg[6]  ( .D(n897), .CLK(CLK), .R(n209), .S(1'b1), .Q(sj[6]) );
  DFFSR \sj_reg[3]  ( .D(n894), .CLK(CLK), .R(n208), .S(1'b1), .Q(sj[3]) );
  DFFSR \sj_reg[2]  ( .D(n893), .CLK(CLK), .R(n208), .S(1'b1), .Q(sj[2]) );
  DFFSR \sj_reg[1]  ( .D(n892), .CLK(CLK), .R(n208), .S(1'b1), .Q(sj[1]) );
  DFFSR \sj_reg[0]  ( .D(n891), .CLK(CLK), .R(n207), .S(1'b1), .Q(sj[0]) );
  DFFPOSX1 \keyi_reg[2]  ( .D(n874), .CLK(CLK), .Q(keyi[2]) );
  DFFPOSX1 \keyi_reg[1]  ( .D(n873), .CLK(CLK), .Q(keyi[1]) );
  DFFPOSX1 \keyi_reg[0]  ( .D(n872), .CLK(CLK), .Q(keyi[0]) );
  DFFPOSX1 \inti_reg[7]  ( .D(n1126), .CLK(CLK), .Q(inti[7]) );
  DFFPOSX1 \inti_reg[0]  ( .D(n1119), .CLK(CLK), .Q(inti[0]) );
  DFFPOSX1 \inti_reg[1]  ( .D(n1120), .CLK(CLK), .Q(inti[1]) );
  DFFPOSX1 \inti_reg[2]  ( .D(n1121), .CLK(CLK), .Q(inti[2]) );
  DFFPOSX1 \inti_reg[3]  ( .D(n1122), .CLK(CLK), .Q(inti[3]) );
  DFFPOSX1 \inti_reg[4]  ( .D(n1123), .CLK(CLK), .Q(inti[4]) );
  DFFPOSX1 \inti_reg[5]  ( .D(n1124), .CLK(CLK), .Q(inti[5]) );
  DFFPOSX1 \inti_reg[6]  ( .D(n1125), .CLK(CLK), .Q(inti[6]) );
  DFFSR \currentProcessedData_reg[0]  ( .D(nextProcessedData[0]), .CLK(CLK), 
        .R(n207), .S(1'b1), .Q(currentProcessedData[0]) );
  DFFPOSX1 \PROCESSED_DATA_reg[0]  ( .D(n759), .CLK(CLK), .Q(PROCESSED_DATA[0]) );
  DFFSR \currentProcessedData_reg[1]  ( .D(nextProcessedData[1]), .CLK(CLK), 
        .R(n206), .S(1'b1), .Q(currentProcessedData[1]) );
  DFFPOSX1 \PROCESSED_DATA_reg[1]  ( .D(n757), .CLK(CLK), .Q(PROCESSED_DATA[1]) );
  DFFSR \currentProcessedData_reg[2]  ( .D(n37), .CLK(CLK), .R(n206), .S(1'b1), 
        .Q(currentProcessedData[2]) );
  DFFPOSX1 \PROCESSED_DATA_reg[2]  ( .D(n755), .CLK(CLK), .Q(PROCESSED_DATA[2]) );
  DFFSR \currentProcessedData_reg[3]  ( .D(n38), .CLK(CLK), .R(n205), .S(1'b1), 
        .Q(currentProcessedData[3]) );
  DFFPOSX1 \PROCESSED_DATA_reg[3]  ( .D(n753), .CLK(CLK), .Q(PROCESSED_DATA[3]) );
  DFFSR \currentProcessedData_reg[4]  ( .D(n39), .CLK(CLK), .R(n205), .S(1'b1), 
        .Q(currentProcessedData[4]) );
  DFFPOSX1 \PROCESSED_DATA_reg[4]  ( .D(n751), .CLK(CLK), .Q(PROCESSED_DATA[4]) );
  DFFSR \currentProcessedData_reg[5]  ( .D(n40), .CLK(CLK), .R(n203), .S(1'b1), 
        .Q(currentProcessedData[5]) );
  DFFPOSX1 \PROCESSED_DATA_reg[5]  ( .D(n749), .CLK(CLK), .Q(PROCESSED_DATA[5]) );
  DFFSR \currentProcessedData_reg[6]  ( .D(n95), .CLK(CLK), .R(n203), .S(1'b1), 
        .Q(currentProcessedData[6]) );
  DFFPOSX1 \PROCESSED_DATA_reg[6]  ( .D(n747), .CLK(CLK), .Q(PROCESSED_DATA[6]) );
  DFFSR \currentProcessedData_reg[7]  ( .D(nextProcessedData[7]), .CLK(CLK), 
        .R(n210), .S(1'b1), .Q(currentProcessedData[7]) );
  DFFPOSX1 \PROCESSED_DATA_reg[7]  ( .D(n745), .CLK(CLK), .Q(PROCESSED_DATA[7]) );
  DFFPOSX1 \faddr_reg[7]  ( .D(n744), .CLK(CLK), .Q(faddr[7]) );
  DFFPOSX1 \ADDR_reg[7]  ( .D(n743), .CLK(CLK), .Q(ADDR[7]) );
  DFFPOSX1 \faddr_reg[6]  ( .D(n742), .CLK(CLK), .Q(faddr[6]) );
  DFFPOSX1 \ADDR_reg[6]  ( .D(n741), .CLK(CLK), .Q(ADDR[6]) );
  DFFPOSX1 \faddr_reg[5]  ( .D(n740), .CLK(CLK), .Q(faddr[5]) );
  DFFPOSX1 \ADDR_reg[5]  ( .D(n739), .CLK(CLK), .Q(ADDR[5]) );
  DFFPOSX1 \faddr_reg[4]  ( .D(n738), .CLK(CLK), .Q(faddr[4]) );
  DFFPOSX1 \ADDR_reg[4]  ( .D(n737), .CLK(CLK), .Q(ADDR[4]) );
  DFFPOSX1 \faddr_reg[3]  ( .D(n736), .CLK(CLK), .Q(faddr[3]) );
  DFFPOSX1 \ADDR_reg[3]  ( .D(n735), .CLK(CLK), .Q(ADDR[3]) );
  DFFPOSX1 \faddr_reg[2]  ( .D(n734), .CLK(CLK), .Q(faddr[2]) );
  DFFPOSX1 \ADDR_reg[2]  ( .D(n733), .CLK(CLK), .Q(ADDR[2]) );
  DFFPOSX1 \faddr_reg[1]  ( .D(n732), .CLK(CLK), .Q(faddr[1]) );
  DFFPOSX1 \ADDR_reg[1]  ( .D(n731), .CLK(CLK), .Q(ADDR[1]) );
  DFFPOSX1 \faddr_reg[0]  ( .D(n730), .CLK(CLK), .Q(faddr[0]) );
  DFFPOSX1 \ADDR_reg[0]  ( .D(n729), .CLK(CLK), .Q(ADDR[0]) );
  DFFPOSX1 \fdata_reg[7]  ( .D(n728), .CLK(CLK), .Q(fdata[7]) );
  DFFPOSX1 \fdata_reg[6]  ( .D(n727), .CLK(CLK), .Q(fdata[6]) );
  DFFPOSX1 \fdata_reg[5]  ( .D(n726), .CLK(CLK), .Q(fdata[5]) );
  DFFPOSX1 \fdata_reg[4]  ( .D(n725), .CLK(CLK), .Q(fdata[4]) );
  DFFPOSX1 \fdata_reg[3]  ( .D(n724), .CLK(CLK), .Q(fdata[3]) );
  DFFPOSX1 \fdata_reg[2]  ( .D(n723), .CLK(CLK), .Q(fdata[2]) );
  DFFPOSX1 \fdata_reg[1]  ( .D(n722), .CLK(CLK), .Q(fdata[1]) );
  DFFPOSX1 \fdata_reg[0]  ( .D(n721), .CLK(CLK), .Q(fdata[0]) );
  DFFPOSX1 fw_enable_reg ( .D(n720), .CLK(CLK), .Q(fw_enable) );
  DFFPOSX1 fr_enable_reg ( .D(n719), .CLK(CLK), .Q(fr_enable) );
  DFFPOSX1 W_ENABLE_reg ( .D(n718), .CLK(CLK), .Q(W_ENABLE) );
  DFFPOSX1 R_ENABLE_reg ( .D(n717), .CLK(CLK), .Q(R_ENABLE) );
  DFFPOSX1 \DATA_reg[7]  ( .D(n716), .CLK(CLK), .Q(DATA[7]) );
  DFFPOSX1 \DATA_reg[6]  ( .D(n715), .CLK(CLK), .Q(DATA[6]) );
  DFFPOSX1 \DATA_reg[5]  ( .D(n714), .CLK(CLK), .Q(DATA[5]) );
  DFFPOSX1 \DATA_reg[4]  ( .D(n713), .CLK(CLK), .Q(DATA[4]) );
  DFFPOSX1 \DATA_reg[3]  ( .D(n712), .CLK(CLK), .Q(DATA[3]) );
  DFFPOSX1 \DATA_reg[2]  ( .D(n711), .CLK(CLK), .Q(DATA[2]) );
  DFFPOSX1 \DATA_reg[1]  ( .D(n710), .CLK(CLK), .Q(DATA[1]) );
  DFFPOSX1 \DATA_reg[0]  ( .D(n709), .CLK(CLK), .Q(DATA[0]) );
  NOR2X1 U110 ( .A(KEY_ERROR), .B(n128), .Y(n126) );
  OAI21X1 U111 ( .A(n1107), .B(n130), .C(n1106), .Y(n124) );
  NOR2X1 U123 ( .A(n159), .B(n1107), .Y(n155) );
  NAND3X1 U126 ( .A(n163), .B(n1101), .C(n165), .Y(nextState[1]) );
  NOR2X1 U130 ( .A(prefillCounter[2]), .B(prefillCounter[1]), .Y(n173) );
  NAND3X1 U131 ( .A(n174), .B(n1136), .C(n176), .Y(n168) );
  NOR2X1 U132 ( .A(prefillCounter[4]), .B(prefillCounter[3]), .Y(n176) );
  NOR2X1 U133 ( .A(prefillCounter[7]), .B(prefillCounter[6]), .Y(n174) );
  NAND3X1 U143 ( .A(n1110), .B(n1109), .C(BYTE_READY), .Y(n158) );
  NAND2X1 U156 ( .A(OPCODE[0]), .B(n1109), .Y(n130) );
  NAND2X1 U158 ( .A(BYTE_READY), .B(n204), .Y(n128) );
  OAI21X1 U159 ( .A(OPCODE[0]), .B(OPCODE[1]), .C(n186), .Y(n204) );
  NAND2X1 U160 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n186) );
  NOR2X1 U669 ( .A(n1104), .B(n1105), .Y(n588) );
  NOR2X1 U673 ( .A(n1102), .B(n1103), .Y(n589) );
  AND2X2 U142 ( .A(n130), .B(n186), .Y(n159) );
  KSA_1_DW01_inc_0 add_289 ( .A({si[7:1], n24}), .SUM({N431, N430, N429, N428, 
        N427, N426, N425, N424}) );
  KSA_1_DW01_inc_1 add_263 ( .A(prefillCounter), .SUM({N414, N413, N412, N411, 
        N410, N409, N408, N407}) );
  KSA_1_DW01_add_6 add_377 ( .A(temp), .B(extratemp), .CI(1'b0), .SUM({N527, 
        N526, N525, N524, N523, N522, N521, N520}) );
  KSA_1_DW01_add_7 add_337 ( .A(intj), .B(DATA_IN), .CI(1'b0), .SUM({N519, 
        N518, N517, N516, N515, N514, N513, N512}) );
  KSA_1_DW01_add_8 add_1_root_add_0_root_add_302_2 ( .A(DATA_IN), .B({sj[7:1], 
        n48}), .CI(1'b0), .SUM({N456, N455, N454, N453, N452, N451, N450, N449}) );
  KSA_1_DW01_add_9 add_0_root_add_0_root_add_302_2 ( .A({N472, N473, N474, 
        N475, N476, N477, N478, N479}), .B({N456, N455, N454, N453, N452, N451, 
        N450, N449}), .CI(1'b0), .SUM({N487, N486, N485, N484, N483, N482, 
        N481, N480}) );
  KSA_1_DW01_inc_3 r126 ( .A(inti), .SUM({N503, N502, N501, N500, N499, N498, 
        N497, N496}) );
  TBUFX1 \nfaddr_tri[0]  ( .A(n708), .EN(n1100), .Y(nfaddr[0]) );
  TBUFX1 \nfaddr_tri[1]  ( .A(n707), .EN(n1100), .Y(nfaddr[1]) );
  TBUFX1 \nfaddr_tri[2]  ( .A(n706), .EN(n1100), .Y(nfaddr[2]) );
  TBUFX1 \nfaddr_tri[3]  ( .A(n705), .EN(n1100), .Y(nfaddr[3]) );
  TBUFX1 \nfaddr_tri[4]  ( .A(n704), .EN(n1100), .Y(nfaddr[4]) );
  TBUFX1 \nfaddr_tri[5]  ( .A(n703), .EN(n1100), .Y(nfaddr[5]) );
  TBUFX1 \nfdata_tri[1]  ( .A(n698), .EN(n29), .Y(nfdata[1]) );
  TBUFX1 \nfdata_tri[2]  ( .A(n697), .EN(n29), .Y(nfdata[2]) );
  TBUFX1 \nfdata_tri[3]  ( .A(n696), .EN(n29), .Y(nfdata[3]) );
  TBUFX1 \nfdata_tri[4]  ( .A(n695), .EN(n29), .Y(nfdata[4]) );
  TBUFX1 \nfdata_tri[5]  ( .A(n694), .EN(n29), .Y(nfdata[5]) );
  TBUFX1 \nfdata_tri[6]  ( .A(n693), .EN(n29), .Y(nfdata[6]) );
  TBUFX1 \nfdata_tri[7]  ( .A(n691), .EN(n29), .Y(nfdata[7]) );
  TBUFX2 \nfaddr_tri[7]  ( .A(n700), .EN(n1100), .Y(nfaddr[7]) );
  TBUFX1 \nfaddr_tri[6]  ( .A(n702), .EN(n1100), .Y(nfaddr[6]) );
  TBUFX1 \nfdata_tri[0]  ( .A(n699), .EN(n29), .Y(nfdata[0]) );
  DFFSR \si_reg[6]  ( .D(n901), .CLK(CLK), .R(n199), .S(1'b1), .Q(si[6]) );
  DFFSR \si_reg[7]  ( .D(n900), .CLK(CLK), .R(n199), .S(1'b1), .Q(si[7]) );
  DFFSR \sj_reg[5]  ( .D(n896), .CLK(CLK), .R(n199), .S(1'b1), .Q(sj[5]) );
  DFFSR \sj_reg[4]  ( .D(n895), .CLK(CLK), .R(n199), .S(1'b1), .Q(sj[4]) );
  INVX8 U3 ( .A(n63), .Y(n136) );
  NAND2X1 U4 ( .A(n54), .B(n1090), .Y(n3) );
  AND2X1 U7 ( .A(n70), .B(n58), .Y(n4) );
  AND2X2 U8 ( .A(n591), .B(n590), .Y(n5) );
  BUFX4 U9 ( .A(n154), .Y(n143) );
  INVX2 U10 ( .A(n31), .Y(n552) );
  INVX2 U11 ( .A(n47), .Y(n563) );
  INVX2 U12 ( .A(n183), .Y(n1081) );
  INVX2 U13 ( .A(n269), .Y(n30) );
  INVX2 U14 ( .A(n188), .Y(n189) );
  INVX2 U15 ( .A(n89), .Y(n67) );
  INVX2 U16 ( .A(n89), .Y(n70) );
  OR2X2 U17 ( .A(n1025), .B(n1024), .Y(n6) );
  INVX2 U18 ( .A(n682), .Y(n429) );
  NAND2X1 U19 ( .A(n135), .B(n1082), .Y(n7) );
  OR2X1 U20 ( .A(n119), .B(n120), .Y(n8) );
  AND2X2 U21 ( .A(n481), .B(n482), .Y(n9) );
  AND2X2 U22 ( .A(n473), .B(n474), .Y(n10) );
  AND2X2 U23 ( .A(n437), .B(n438), .Y(n11) );
  AND2X2 U24 ( .A(n107), .B(n76), .Y(n12) );
  NAND3X1 U29 ( .A(n162), .B(n70), .C(n238), .Y(n17) );
  INVX2 U30 ( .A(n244), .Y(n18) );
  BUFX2 U31 ( .A(n242), .Y(n142) );
  BUFX2 U32 ( .A(n72), .Y(n19) );
  AOI21X1 U33 ( .A(n177), .B(n18), .C(n88), .Y(n20) );
  BUFX4 U34 ( .A(n1026), .Y(n21) );
  NOR2X1 U35 ( .A(n75), .B(n74), .Y(n22) );
  AND2X2 U36 ( .A(n433), .B(n432), .Y(n23) );
  BUFX2 U37 ( .A(si[0]), .Y(n24) );
  AND2X2 U38 ( .A(n49), .B(n32), .Y(n25) );
  INVX2 U39 ( .A(n25), .Y(n240) );
  INVX2 U40 ( .A(n240), .Y(n1046) );
  AND2X2 U41 ( .A(n64), .B(n237), .Y(n26) );
  INVX1 U42 ( .A(n1060), .Y(n1084) );
  INVX1 U43 ( .A(n66), .Y(n27) );
  INVX2 U44 ( .A(n49), .Y(n243) );
  INVX1 U45 ( .A(n119), .Y(n28) );
  INVX2 U46 ( .A(n135), .Y(n119) );
  INVX4 U47 ( .A(n76), .Y(n223) );
  INVX1 U48 ( .A(n645), .Y(n29) );
  NOR3X1 U49 ( .A(n510), .B(n512), .C(keyi[2]), .Y(n31) );
  INVX4 U50 ( .A(keyi[1]), .Y(n510) );
  INVX4 U51 ( .A(keyi[0]), .Y(n512) );
  INVX4 U52 ( .A(keyi[2]), .Y(n511) );
  BUFX2 U53 ( .A(n161), .Y(n32) );
  NAND2X1 U54 ( .A(n644), .B(n115), .Y(n33) );
  INVX2 U55 ( .A(n114), .Y(n115) );
  INVX1 U56 ( .A(n18), .Y(n34) );
  INVX1 U57 ( .A(n7), .Y(n645) );
  MUX2X1 U58 ( .B(n640), .A(n511), .S(n35), .Y(n874) );
  NAND2X1 U59 ( .A(n92), .B(n563), .Y(n35) );
  INVX1 U60 ( .A(n429), .Y(n36) );
  INVX1 U61 ( .A(n471), .Y(n37) );
  INVX1 U62 ( .A(n465), .Y(n38) );
  INVX1 U63 ( .A(n459), .Y(n39) );
  INVX1 U64 ( .A(n453), .Y(n40) );
  NAND2X1 U65 ( .A(n41), .B(n432), .Y(n297) );
  NOR2X1 U66 ( .A(n47), .B(n1135), .Y(n41) );
  INVX2 U67 ( .A(n101), .Y(n432) );
  AND2X2 U68 ( .A(n183), .B(n161), .Y(n62) );
  AND2X1 U69 ( .A(n680), .B(n681), .Y(n42) );
  NAND2X1 U70 ( .A(n644), .B(n115), .Y(n43) );
  NAND2X1 U71 ( .A(n644), .B(n115), .Y(n44) );
  INVX1 U72 ( .A(n487), .Y(n45) );
  INVX1 U73 ( .A(n45), .Y(n46) );
  NAND2X1 U74 ( .A(n188), .B(n273), .Y(n242) );
  BUFX2 U75 ( .A(state[2]), .Y(n179) );
  AND2X2 U76 ( .A(n178), .B(n1082), .Y(n47) );
  BUFX4 U77 ( .A(sj[0]), .Y(n48) );
  AND2X2 U78 ( .A(n189), .B(n273), .Y(n49) );
  NAND3X1 U79 ( .A(n96), .B(n110), .C(n223), .Y(n50) );
  NOR2X1 U80 ( .A(n562), .B(n47), .Y(n51) );
  INVX2 U81 ( .A(n57), .Y(n562) );
  BUFX2 U82 ( .A(n562), .Y(n52) );
  BUFX4 U83 ( .A(n185), .Y(n53) );
  AND2X2 U84 ( .A(n585), .B(n1048), .Y(n54) );
  INVX4 U85 ( .A(n5), .Y(n55) );
  MUX2X1 U86 ( .B(n1102), .A(n512), .S(n56), .Y(n872) );
  NAND2X1 U87 ( .A(n563), .B(n92), .Y(n56) );
  AND2X2 U88 ( .A(n670), .B(n646), .Y(n57) );
  INVX2 U89 ( .A(n1077), .Y(n58) );
  AND2X2 U90 ( .A(n90), .B(n638), .Y(n59) );
  INVX1 U91 ( .A(n59), .Y(n328) );
  INVX1 U92 ( .A(n434), .Y(n479) );
  AND2X2 U93 ( .A(n7), .B(n42), .Y(n60) );
  INVX1 U94 ( .A(n60), .Y(n1025) );
  MUX2X1 U95 ( .B(fdata[7]), .A(nfdata[7]), .S(n206), .Y(n412) );
  MUX2X1 U96 ( .B(fdata[6]), .A(nfdata[6]), .S(n205), .Y(n411) );
  MUX2X1 U97 ( .B(fdata[5]), .A(nfdata[5]), .S(n205), .Y(n410) );
  MUX2X1 U98 ( .B(fdata[4]), .A(nfdata[4]), .S(n205), .Y(n409) );
  MUX2X1 U99 ( .B(fdata[3]), .A(nfdata[3]), .S(n205), .Y(n408) );
  MUX2X1 U100 ( .B(fdata[2]), .A(nfdata[2]), .S(n205), .Y(n407) );
  MUX2X1 U101 ( .B(fdata[1]), .A(nfdata[1]), .S(n205), .Y(n406) );
  MUX2X1 U102 ( .B(fdata[0]), .A(nfdata[0]), .S(n205), .Y(n405) );
  MUX2X1 U103 ( .B(DATA[7]), .A(nfdata[7]), .S(n205), .Y(n386) );
  MUX2X1 U104 ( .B(DATA[6]), .A(nfdata[6]), .S(n205), .Y(n385) );
  MUX2X1 U105 ( .B(DATA[5]), .A(nfdata[5]), .S(n205), .Y(n384) );
  MUX2X1 U106 ( .B(DATA[4]), .A(nfdata[4]), .S(n203), .Y(n383) );
  MUX2X1 U107 ( .B(DATA[3]), .A(nfdata[3]), .S(n203), .Y(n382) );
  MUX2X1 U108 ( .B(DATA[2]), .A(nfdata[2]), .S(n203), .Y(n381) );
  MUX2X1 U109 ( .B(DATA[1]), .A(nfdata[1]), .S(n205), .Y(n380) );
  AND2X2 U112 ( .A(n682), .B(n153), .Y(n430) );
  MUX2X1 U113 ( .B(DATA[0]), .A(nfdata[0]), .S(n199), .Y(n379) );
  MUX2X1 U114 ( .B(n1103), .A(n510), .S(n61), .Y(n873) );
  NAND2X1 U115 ( .A(n563), .B(n92), .Y(n61) );
  INVX1 U116 ( .A(n62), .Y(n274) );
  INVX2 U117 ( .A(n108), .Y(n63) );
  INVX2 U118 ( .A(n108), .Y(n154) );
  BUFX4 U119 ( .A(state[4]), .Y(n197) );
  AND2X2 U120 ( .A(n182), .B(n139), .Y(n64) );
  INVX1 U121 ( .A(n64), .Y(n220) );
  INVX1 U122 ( .A(n66), .Y(n111) );
  NAND2X1 U124 ( .A(n246), .B(n1082), .Y(n65) );
  BUFX2 U125 ( .A(state[1]), .Y(n66) );
  NAND2X1 U127 ( .A(n684), .B(n141), .Y(n68) );
  INVX4 U128 ( .A(n237), .Y(n105) );
  NAND2X1 U129 ( .A(n237), .B(n169), .Y(n69) );
  INVX2 U134 ( .A(n69), .Y(n135) );
  INVX1 U135 ( .A(n194), .Y(n131) );
  BUFX2 U136 ( .A(state[0]), .Y(n182) );
  INVX1 U137 ( .A(sj[2]), .Y(n572) );
  INVX2 U138 ( .A(n297), .Y(n71) );
  AND2X2 U139 ( .A(n96), .B(n64), .Y(n72) );
  NOR2X1 U140 ( .A(n47), .B(n156), .Y(n73) );
  NOR2X1 U141 ( .A(n75), .B(n74), .Y(n565) );
  INVX1 U144 ( .A(n73), .Y(n74) );
  BUFX4 U145 ( .A(n564), .Y(n75) );
  NOR2X1 U146 ( .A(n94), .B(n486), .Y(n629) );
  INVX1 U147 ( .A(n486), .Y(n1100) );
  INVX4 U148 ( .A(n133), .Y(n1135) );
  BUFX4 U149 ( .A(state[0]), .Y(n76) );
  NAND2X1 U150 ( .A(n190), .B(n51), .Y(n1026) );
  AND2X2 U151 ( .A(n18), .B(n1071), .Y(n156) );
  INVX4 U152 ( .A(n195), .Y(n196) );
  INVX8 U153 ( .A(n136), .Y(n77) );
  INVX8 U154 ( .A(n136), .Y(n78) );
  INVX4 U155 ( .A(n148), .Y(n79) );
  INVX8 U157 ( .A(n79), .Y(n80) );
  INVX4 U161 ( .A(n198), .Y(n81) );
  INVX8 U162 ( .A(n81), .Y(n82) );
  NOR2X1 U163 ( .A(n245), .B(n25), .Y(n83) );
  AND2X2 U164 ( .A(n83), .B(n84), .Y(n289) );
  AND2X1 U165 ( .A(n8), .B(n670), .Y(n84) );
  INVX1 U166 ( .A(n50), .Y(n85) );
  INVX1 U167 ( .A(n50), .Y(n246) );
  AND2X2 U168 ( .A(n566), .B(n86), .Y(n152) );
  AND2X1 U169 ( .A(n565), .B(n591), .Y(n86) );
  BUFX2 U170 ( .A(n169), .Y(n87) );
  INVX1 U171 ( .A(n436), .Y(n480) );
  INVX4 U172 ( .A(n297), .Y(n650) );
  INVX2 U173 ( .A(n139), .Y(n184) );
  AND2X2 U174 ( .A(n32), .B(n1082), .Y(n88) );
  INVX2 U175 ( .A(n88), .Y(n560) );
  AND2X1 U176 ( .A(n193), .B(n123), .Y(n649) );
  INVX2 U177 ( .A(n131), .Y(n132) );
  AND2X2 U178 ( .A(n167), .B(n26), .Y(n89) );
  NOR2X1 U179 ( .A(n354), .B(si[2]), .Y(n90) );
  INVX1 U180 ( .A(n90), .Y(n341) );
  INVX1 U181 ( .A(si[2]), .Y(n640) );
  NOR2X1 U182 ( .A(n1046), .B(n245), .Y(n91) );
  AND2X2 U183 ( .A(n507), .B(n4), .Y(n92) );
  INVX1 U184 ( .A(n92), .Y(n1057) );
  BUFX2 U185 ( .A(n1089), .Y(n93) );
  INVX1 U186 ( .A(si[1]), .Y(n1103) );
  NAND2X1 U187 ( .A(n70), .B(n563), .Y(n94) );
  NAND2X1 U188 ( .A(n483), .B(n9), .Y(nextProcessedData[0]) );
  INVX1 U189 ( .A(nextProcessedData[0]), .Y(n485) );
  NAND2X1 U190 ( .A(n475), .B(n10), .Y(nextProcessedData[1]) );
  INVX1 U191 ( .A(nextProcessedData[1]), .Y(n477) );
  INVX1 U192 ( .A(n447), .Y(n95) );
  BUFX4 U193 ( .A(state[4]), .Y(n96) );
  OR2X1 U194 ( .A(n562), .B(n561), .Y(n97) );
  NAND2X1 U195 ( .A(n1090), .B(n157), .Y(n98) );
  INVX4 U196 ( .A(n195), .Y(n99) );
  INVX1 U197 ( .A(n223), .Y(n100) );
  NAND2X1 U198 ( .A(n121), .B(n20), .Y(n101) );
  NAND2X1 U199 ( .A(n23), .B(n629), .Y(n102) );
  NAND2X1 U200 ( .A(n23), .B(n629), .Y(n103) );
  NAND2X1 U201 ( .A(n289), .B(n54), .Y(n104) );
  INVX2 U202 ( .A(n195), .Y(n122) );
  INVX1 U203 ( .A(n785), .Y(n683) );
  BUFX2 U204 ( .A(n585), .Y(n106) );
  AND2X1 U205 ( .A(n328), .B(si[4]), .Y(n316) );
  INVX1 U206 ( .A(n24), .Y(n1102) );
  OR2X2 U207 ( .A(n213), .B(n181), .Y(n1065) );
  INVX1 U208 ( .A(n144), .Y(n107) );
  INVX4 U209 ( .A(n674), .Y(n195) );
  INVX1 U210 ( .A(n412), .Y(n728) );
  INVX1 U211 ( .A(n411), .Y(n727) );
  INVX1 U212 ( .A(n410), .Y(n726) );
  INVX1 U213 ( .A(n409), .Y(n725) );
  INVX1 U214 ( .A(n408), .Y(n724) );
  INVX1 U215 ( .A(n407), .Y(n723) );
  INVX1 U216 ( .A(n406), .Y(n722) );
  INVX1 U217 ( .A(n386), .Y(n716) );
  INVX1 U218 ( .A(n385), .Y(n715) );
  INVX1 U219 ( .A(n384), .Y(n714) );
  INVX1 U220 ( .A(n383), .Y(n713) );
  INVX1 U221 ( .A(n382), .Y(n712) );
  INVX1 U222 ( .A(n381), .Y(n711) );
  INVX1 U223 ( .A(n380), .Y(n710) );
  NAND2X1 U224 ( .A(n786), .B(n190), .Y(n108) );
  INVX2 U225 ( .A(n122), .Y(n151) );
  BUFX2 U226 ( .A(n160), .Y(n109) );
  INVX1 U227 ( .A(n66), .Y(n110) );
  INVX1 U228 ( .A(n66), .Y(n144) );
  BUFX2 U229 ( .A(n190), .Y(n112) );
  BUFX2 U230 ( .A(n305), .Y(n113) );
  INVX1 U231 ( .A(n507), .Y(n114) );
  AND2X2 U232 ( .A(n305), .B(n275), .Y(n116) );
  AND2X1 U233 ( .A(n113), .B(n275), .Y(n171) );
  NAND2X1 U234 ( .A(n23), .B(n629), .Y(n117) );
  NAND2X1 U235 ( .A(n23), .B(n629), .Y(n118) );
  INVX8 U236 ( .A(n99), .Y(n675) );
  INVX1 U237 ( .A(n428), .Y(n744) );
  AND2X1 U238 ( .A(n303), .B(si[5]), .Y(n304) );
  INVX1 U239 ( .A(n427), .Y(n743) );
  INVX2 U240 ( .A(n1071), .Y(n120) );
  NOR2X1 U241 ( .A(n194), .B(n97), .Y(n566) );
  AND2X2 U242 ( .A(n146), .B(n1060), .Y(n121) );
  INVX1 U243 ( .A(n121), .Y(n1050) );
  INVX4 U244 ( .A(n125), .Y(n608) );
  NOR2X1 U245 ( .A(n648), .B(n684), .Y(n123) );
  AND2X2 U246 ( .A(n224), .B(n152), .Y(n125) );
  INVX1 U247 ( .A(n187), .Y(n127) );
  INVX1 U248 ( .A(n187), .Y(n129) );
  NOR2X1 U249 ( .A(n197), .B(n1045), .Y(n161) );
  AND2X2 U250 ( .A(n434), .B(n436), .Y(n133) );
  BUFX2 U251 ( .A(n49), .Y(n134) );
  NAND2X1 U252 ( .A(n439), .B(n11), .Y(nextProcessedData[7]) );
  INVX1 U253 ( .A(nextProcessedData[7]), .Y(n441) );
  INVX1 U254 ( .A(state[2]), .Y(n273) );
  INVX8 U255 ( .A(n136), .Y(n137) );
  INVX2 U256 ( .A(state[1]), .Y(n139) );
  NOR3X1 U257 ( .A(n75), .B(n156), .C(n194), .Y(n138) );
  INVX4 U258 ( .A(n193), .Y(n194) );
  NOR2X1 U259 ( .A(n144), .B(n76), .Y(n140) );
  AND2X2 U260 ( .A(n683), .B(n112), .Y(n141) );
  INVX4 U261 ( .A(n141), .Y(n149) );
  BUFX2 U262 ( .A(n154), .Y(n148) );
  NOR2X1 U263 ( .A(n1135), .B(n431), .Y(n145) );
  INVX1 U264 ( .A(n145), .Y(n387) );
  AND2X2 U265 ( .A(n487), .B(n1074), .Y(n146) );
  INVX1 U266 ( .A(n146), .Y(n1085) );
  INVX2 U267 ( .A(n67), .Y(n644) );
  NAND2X1 U268 ( .A(n167), .B(n28), .Y(n147) );
  NOR2X1 U269 ( .A(n27), .B(n76), .Y(n169) );
  AND2X1 U270 ( .A(n88), .B(n1055), .Y(n166) );
  AND2X1 U271 ( .A(keyi[2]), .B(keyi[1]), .Y(n172) );
  INVX1 U272 ( .A(n19), .Y(n150) );
  INVX2 U273 ( .A(n205), .Y(n202) );
  INVX2 U274 ( .A(n206), .Y(n201) );
  INVX2 U275 ( .A(n207), .Y(n200) );
  BUFX2 U276 ( .A(n154), .Y(n198) );
  INVX4 U277 ( .A(n1027), .Y(n1042) );
  BUFX2 U278 ( .A(n199), .Y(n203) );
  BUFX2 U279 ( .A(n212), .Y(n205) );
  BUFX2 U280 ( .A(n199), .Y(n206) );
  BUFX2 U281 ( .A(n212), .Y(n207) );
  BUFX2 U282 ( .A(n199), .Y(n208) );
  BUFX2 U283 ( .A(n199), .Y(n209) );
  BUFX2 U284 ( .A(n199), .Y(n210) );
  BUFX2 U285 ( .A(n199), .Y(n211) );
  BUFX2 U286 ( .A(n199), .Y(n212) );
  AND2X2 U287 ( .A(n278), .B(n1065), .Y(n153) );
  AND2X2 U288 ( .A(n585), .B(n1048), .Y(n157) );
  INVX2 U289 ( .A(n1081), .Y(n177) );
  AND2X2 U290 ( .A(n183), .B(n140), .Y(n160) );
  AND2X2 U291 ( .A(n1089), .B(n236), .Y(n162) );
  INVX2 U292 ( .A(RST), .Y(n199) );
  AND2X2 U293 ( .A(n172), .B(n512), .Y(n164) );
  AND2X2 U294 ( .A(n189), .B(n179), .Y(n167) );
  AND2X2 U295 ( .A(n172), .B(keyi[0]), .Y(n170) );
  INVX1 U296 ( .A(n405), .Y(n721) );
  INVX1 U297 ( .A(n379), .Y(n709) );
  INVX4 U298 ( .A(n242), .Y(n1082) );
  INVX1 U299 ( .A(n189), .Y(n1071) );
  INVX4 U300 ( .A(n197), .Y(n237) );
  NOR2X1 U301 ( .A(n182), .B(n184), .Y(n175) );
  AND2X2 U302 ( .A(n175), .B(n237), .Y(n178) );
  AND2X1 U303 ( .A(n175), .B(n237), .Y(n180) );
  INVX2 U304 ( .A(n181), .Y(n183) );
  NAND2X1 U305 ( .A(n188), .B(n179), .Y(n181) );
  INVX1 U306 ( .A(n147), .Y(n224) );
  INVX1 U307 ( .A(n1074), .Y(n1077) );
  OR2X2 U308 ( .A(n6), .B(n1026), .Y(n1027) );
  INVX1 U309 ( .A(n153), .Y(n185) );
  INVX1 U310 ( .A(n681), .Y(n268) );
  INVX1 U311 ( .A(n53), .Y(n1075) );
  INVX1 U312 ( .A(n670), .Y(n676) );
  AND2X2 U313 ( .A(n276), .B(n681), .Y(n187) );
  INVX2 U314 ( .A(state[3]), .Y(n188) );
  AND2X2 U315 ( .A(n239), .B(n145), .Y(n190) );
  INVX1 U316 ( .A(n112), .Y(n401) );
  AND2X2 U317 ( .A(n152), .B(n58), .Y(n191) );
  AND2X2 U318 ( .A(n152), .B(n58), .Y(n192) );
  INVX1 U319 ( .A(n1065), .Y(n269) );
  AND2X1 U320 ( .A(n1065), .B(n208), .Y(n680) );
  INVX2 U321 ( .A(n647), .Y(n193) );
  INVX4 U322 ( .A(n1022), .Y(n684) );
  INVX2 U323 ( .A(si[4]), .Y(n1104) );
  INVX2 U324 ( .A(si[5]), .Y(n1105) );
  INVX2 U325 ( .A(prefillCounter[5]), .Y(n1136) );
  NAND3X1 U326 ( .A(n167), .B(n175), .C(n237), .Y(n1074) );
  NAND3X1 U327 ( .A(n111), .B(n96), .C(n223), .Y(n213) );
  NAND2X1 U328 ( .A(n85), .B(n167), .Y(n487) );
  INVX2 U329 ( .A(n158), .Y(n214) );
  NAND2X1 U330 ( .A(n1085), .B(n214), .Y(n219) );
  NAND2X1 U331 ( .A(n105), .B(n64), .Y(n232) );
  NAND3X1 U332 ( .A(n96), .B(n184), .C(n76), .Y(n241) );
  INVX2 U333 ( .A(n241), .Y(n215) );
  OAI21X1 U334 ( .A(n159), .B(n1107), .C(n215), .Y(n216) );
  OAI21X1 U335 ( .A(n158), .B(n150), .C(n216), .Y(n217) );
  NAND2X1 U336 ( .A(n134), .B(n217), .Y(n218) );
  NAND2X1 U337 ( .A(n219), .B(n218), .Y(n222) );
  NOR2X1 U338 ( .A(n220), .B(n142), .Y(n221) );
  AOI21X1 U339 ( .A(n1106), .B(n222), .C(n221), .Y(n163) );
  NAND2X1 U340 ( .A(n160), .B(n237), .Y(n1090) );
  NAND2X1 U341 ( .A(n184), .B(n182), .Y(n1045) );
  INVX2 U342 ( .A(permuteComplete), .Y(n1054) );
  NAND2X1 U343 ( .A(n167), .B(n135), .Y(n1048) );
  AOI21X1 U344 ( .A(n1046), .B(n1054), .C(n224), .Y(n227) );
  NAND2X1 U345 ( .A(n160), .B(n105), .Y(n1089) );
  XOR2X1 U346 ( .A(n189), .B(n96), .Y(n225) );
  NAND3X1 U347 ( .A(n87), .B(n225), .C(n273), .Y(n682) );
  AND2X2 U348 ( .A(n93), .B(n36), .Y(n226) );
  NAND3X1 U349 ( .A(n1090), .B(n227), .C(n226), .Y(n1067) );
  INVX2 U350 ( .A(n1067), .Y(n1101) );
  NOR2X1 U351 ( .A(prefillCounter[0]), .B(n168), .Y(n228) );
  NAND3X1 U352 ( .A(n173), .B(n645), .C(n228), .Y(n229) );
  NAND3X1 U353 ( .A(n49), .B(n140), .C(n105), .Y(n436) );
  NAND2X1 U354 ( .A(n229), .B(n436), .Y(n231) );
  NAND2X1 U355 ( .A(n177), .B(n72), .Y(n670) );
  NAND2X1 U356 ( .A(n64), .B(n237), .Y(n244) );
  NAND2X1 U357 ( .A(n670), .B(n34), .Y(n230) );
  NOR2X1 U358 ( .A(n231), .B(n230), .Y(n165) );
  NAND2X1 U359 ( .A(n246), .B(n49), .Y(n434) );
  AOI21X1 U360 ( .A(n177), .B(n26), .C(n88), .Y(n234) );
  NAND2X1 U361 ( .A(n241), .B(n232), .Y(n233) );
  NAND2X1 U362 ( .A(n49), .B(n233), .Y(n1060) );
  NAND2X1 U363 ( .A(n234), .B(n121), .Y(n431) );
  NAND2X1 U364 ( .A(n246), .B(n1082), .Y(n1070) );
  OAI21X1 U365 ( .A(n1081), .B(n241), .C(n1070), .Y(n235) );
  INVX2 U366 ( .A(n235), .Y(n585) );
  AOI21X1 U367 ( .A(n72), .B(n1082), .C(n62), .Y(n236) );
  NAND2X1 U368 ( .A(n178), .B(n183), .Y(n276) );
  NAND2X1 U369 ( .A(n167), .B(n32), .Y(n278) );
  AND2X2 U370 ( .A(n276), .B(n278), .Y(n238) );
  NAND3X1 U371 ( .A(n162), .B(n67), .C(n238), .Y(n398) );
  NOR2X1 U372 ( .A(n398), .B(n98), .Y(n239) );
  OAI22X1 U373 ( .A(n244), .B(n243), .C(n142), .D(n241), .Y(n245) );
  NOR2X1 U374 ( .A(n25), .B(n245), .Y(n646) );
  NAND2X1 U375 ( .A(n180), .B(n49), .Y(n681) );
  NAND2X1 U376 ( .A(n268), .B(DATA_IN[7]), .Y(n248) );
  NAND2X1 U377 ( .A(n1082), .B(n26), .Y(n1022) );
  NAND2X1 U378 ( .A(prefillCounter[7]), .B(n684), .Y(n282) );
  AOI22X1 U379 ( .A(extratemp[7]), .B(n269), .C(n429), .D(temp[7]), .Y(n247)
         );
  NAND3X1 U380 ( .A(n248), .B(n282), .C(n247), .Y(n249) );
  AOI21X1 U381 ( .A(n21), .B(fdata[7]), .C(n249), .Y(n691) );
  NAND2X1 U382 ( .A(n268), .B(DATA_IN[6]), .Y(n251) );
  NAND2X1 U383 ( .A(prefillCounter[6]), .B(n684), .Y(n295) );
  AOI22X1 U384 ( .A(extratemp[6]), .B(n269), .C(n429), .D(temp[6]), .Y(n250)
         );
  NAND3X1 U385 ( .A(n251), .B(n295), .C(n250), .Y(n252) );
  AOI21X1 U386 ( .A(n21), .B(fdata[6]), .C(n252), .Y(n693) );
  NAND2X1 U387 ( .A(n268), .B(DATA_IN[5]), .Y(n254) );
  NAND2X1 U388 ( .A(n684), .B(prefillCounter[5]), .Y(n309) );
  AOI22X1 U389 ( .A(extratemp[5]), .B(n269), .C(n429), .D(temp[5]), .Y(n253)
         );
  NAND3X1 U390 ( .A(n254), .B(n309), .C(n253), .Y(n255) );
  AOI21X1 U391 ( .A(n21), .B(fdata[5]), .C(n255), .Y(n694) );
  NAND2X1 U392 ( .A(n268), .B(DATA_IN[4]), .Y(n257) );
  NAND2X1 U393 ( .A(prefillCounter[4]), .B(n684), .Y(n321) );
  AOI22X1 U394 ( .A(extratemp[4]), .B(n269), .C(n429), .D(temp[4]), .Y(n256)
         );
  NAND3X1 U395 ( .A(n257), .B(n321), .C(n256), .Y(n258) );
  AOI21X1 U396 ( .A(n21), .B(fdata[4]), .C(n258), .Y(n695) );
  NAND2X1 U397 ( .A(n268), .B(DATA_IN[3]), .Y(n260) );
  NAND2X1 U398 ( .A(prefillCounter[3]), .B(n684), .Y(n334) );
  AOI22X1 U399 ( .A(extratemp[3]), .B(n269), .C(n429), .D(temp[3]), .Y(n259)
         );
  NAND3X1 U400 ( .A(n260), .B(n334), .C(n259), .Y(n261) );
  AOI21X1 U401 ( .A(n21), .B(fdata[3]), .C(n261), .Y(n696) );
  NAND2X1 U402 ( .A(n268), .B(DATA_IN[2]), .Y(n263) );
  NAND2X1 U403 ( .A(prefillCounter[2]), .B(n684), .Y(n347) );
  AOI22X1 U404 ( .A(extratemp[2]), .B(n269), .C(n429), .D(temp[2]), .Y(n262)
         );
  NAND3X1 U405 ( .A(n263), .B(n347), .C(n262), .Y(n264) );
  AOI21X1 U406 ( .A(n21), .B(fdata[2]), .C(n264), .Y(n697) );
  NAND2X1 U407 ( .A(n268), .B(DATA_IN[1]), .Y(n266) );
  NAND2X1 U408 ( .A(prefillCounter[1]), .B(n684), .Y(n360) );
  AOI22X1 U409 ( .A(extratemp[1]), .B(n269), .C(n429), .D(temp[1]), .Y(n265)
         );
  NAND3X1 U410 ( .A(n266), .B(n360), .C(n265), .Y(n267) );
  AOI21X1 U411 ( .A(n21), .B(fdata[1]), .C(n267), .Y(n698) );
  NAND2X1 U412 ( .A(n268), .B(DATA_IN[0]), .Y(n271) );
  NAND2X1 U413 ( .A(prefillCounter[0]), .B(n684), .Y(n371) );
  AOI22X1 U414 ( .A(extratemp[0]), .B(n269), .C(n429), .D(temp[0]), .Y(n270)
         );
  NAND3X1 U415 ( .A(n271), .B(n371), .C(n270), .Y(n272) );
  AOI21X1 U416 ( .A(n21), .B(fdata[0]), .C(n272), .Y(n699) );
  NAND2X1 U417 ( .A(n135), .B(n273), .Y(n388) );
  NAND2X1 U418 ( .A(n388), .B(n274), .Y(n367) );
  OR2X2 U419 ( .A(si[1]), .B(si[0]), .Y(n354) );
  INVX2 U420 ( .A(si[3]), .Y(n638) );
  NAND2X1 U421 ( .A(n59), .B(n1104), .Y(n303) );
  INVX2 U422 ( .A(n303), .Y(n317) );
  NAND2X1 U423 ( .A(n317), .B(n1105), .Y(n290) );
  INVX2 U424 ( .A(n290), .Y(n305) );
  INVX2 U425 ( .A(si[6]), .Y(n275) );
  XOR2X1 U426 ( .A(n116), .B(si[7]), .Y(n277) );
  AOI22X1 U427 ( .A(sj[7]), .B(n367), .C(n277), .D(n127), .Y(n287) );
  AOI22X1 U428 ( .A(N503), .B(n644), .C(intj[7]), .D(n53), .Y(n286) );
  AND2X2 U429 ( .A(faddr[7]), .B(n297), .Y(n284) );
  NAND2X1 U430 ( .A(temp[7]), .B(n109), .Y(n281) );
  OAI21X1 U431 ( .A(n87), .B(n19), .C(n1082), .Y(n279) );
  INVX2 U432 ( .A(n279), .Y(n373) );
  NAND2X1 U433 ( .A(n373), .B(inti[7]), .Y(n280) );
  NAND3X1 U434 ( .A(n282), .B(n281), .C(n280), .Y(n283) );
  NOR2X1 U435 ( .A(n284), .B(n283), .Y(n285) );
  NAND3X1 U436 ( .A(n287), .B(n286), .C(n285), .Y(n288) );
  INVX2 U437 ( .A(n288), .Y(n700) );
  NAND2X1 U438 ( .A(n54), .B(n289), .Y(n486) );
  NAND2X1 U439 ( .A(sj[6]), .B(n367), .Y(n294) );
  AND2X2 U440 ( .A(si[6]), .B(n290), .Y(n291) );
  OAI21X1 U441 ( .A(n171), .B(n291), .C(n127), .Y(n293) );
  AOI22X1 U442 ( .A(intj[6]), .B(n53), .C(N502), .D(n644), .Y(n292) );
  NAND3X1 U443 ( .A(n294), .B(n293), .C(n292), .Y(n302) );
  NAND2X1 U444 ( .A(temp[6]), .B(n109), .Y(n296) );
  NAND2X1 U445 ( .A(n296), .B(n295), .Y(n301) );
  INVX2 U446 ( .A(faddr[6]), .Y(n299) );
  NAND2X1 U447 ( .A(n373), .B(inti[6]), .Y(n298) );
  OAI21X1 U448 ( .A(n650), .B(n299), .C(n298), .Y(n300) );
  NOR3X1 U449 ( .A(n302), .B(n301), .C(n300), .Y(n702) );
  NAND2X1 U450 ( .A(sj[5]), .B(n367), .Y(n308) );
  OAI21X1 U451 ( .A(n113), .B(n304), .C(n129), .Y(n307) );
  AOI22X1 U452 ( .A(intj[5]), .B(n53), .C(N501), .D(n644), .Y(n306) );
  NAND3X1 U453 ( .A(n308), .B(n307), .C(n306), .Y(n315) );
  NAND2X1 U454 ( .A(temp[5]), .B(n109), .Y(n310) );
  NAND2X1 U455 ( .A(n310), .B(n309), .Y(n314) );
  INVX2 U456 ( .A(faddr[5]), .Y(n312) );
  NAND2X1 U457 ( .A(n373), .B(inti[5]), .Y(n311) );
  OAI21X1 U458 ( .A(n650), .B(n312), .C(n311), .Y(n313) );
  NOR3X1 U459 ( .A(n315), .B(n314), .C(n313), .Y(n703) );
  NAND2X1 U460 ( .A(sj[4]), .B(n367), .Y(n320) );
  OAI21X1 U461 ( .A(n317), .B(n316), .C(n127), .Y(n319) );
  AOI22X1 U462 ( .A(intj[4]), .B(n53), .C(N500), .D(n644), .Y(n318) );
  NAND3X1 U463 ( .A(n320), .B(n319), .C(n318), .Y(n327) );
  NAND2X1 U464 ( .A(temp[4]), .B(n109), .Y(n322) );
  NAND2X1 U465 ( .A(n322), .B(n321), .Y(n326) );
  INVX2 U466 ( .A(faddr[4]), .Y(n324) );
  NAND2X1 U467 ( .A(n373), .B(inti[4]), .Y(n323) );
  OAI21X1 U468 ( .A(n650), .B(n324), .C(n323), .Y(n325) );
  NOR3X1 U469 ( .A(n327), .B(n326), .C(n325), .Y(n704) );
  NAND2X1 U470 ( .A(sj[3]), .B(n367), .Y(n333) );
  NAND2X1 U471 ( .A(si[3]), .B(n341), .Y(n329) );
  NAND2X1 U472 ( .A(n329), .B(n328), .Y(n330) );
  NAND2X1 U473 ( .A(n330), .B(n129), .Y(n332) );
  AOI22X1 U474 ( .A(intj[3]), .B(n53), .C(N499), .D(n644), .Y(n331) );
  NAND3X1 U475 ( .A(n333), .B(n332), .C(n331), .Y(n340) );
  NAND2X1 U476 ( .A(temp[3]), .B(n109), .Y(n335) );
  NAND2X1 U477 ( .A(n335), .B(n334), .Y(n339) );
  INVX2 U478 ( .A(faddr[3]), .Y(n337) );
  NAND2X1 U479 ( .A(n373), .B(inti[3]), .Y(n336) );
  OAI21X1 U480 ( .A(n650), .B(n337), .C(n336), .Y(n338) );
  NOR3X1 U481 ( .A(n340), .B(n339), .C(n338), .Y(n705) );
  NAND2X1 U482 ( .A(sj[2]), .B(n367), .Y(n346) );
  NAND2X1 U483 ( .A(si[2]), .B(n354), .Y(n342) );
  NAND2X1 U484 ( .A(n342), .B(n341), .Y(n343) );
  NAND2X1 U485 ( .A(n343), .B(n127), .Y(n345) );
  AOI22X1 U486 ( .A(intj[2]), .B(n53), .C(N498), .D(n644), .Y(n344) );
  NAND3X1 U487 ( .A(n346), .B(n345), .C(n344), .Y(n353) );
  NAND2X1 U488 ( .A(temp[2]), .B(n109), .Y(n348) );
  NAND2X1 U489 ( .A(n348), .B(n347), .Y(n352) );
  INVX2 U490 ( .A(faddr[2]), .Y(n350) );
  NAND2X1 U491 ( .A(n373), .B(inti[2]), .Y(n349) );
  OAI21X1 U492 ( .A(n650), .B(n350), .C(n349), .Y(n351) );
  NOR3X1 U493 ( .A(n353), .B(n352), .C(n351), .Y(n706) );
  NAND2X1 U494 ( .A(sj[1]), .B(n367), .Y(n359) );
  NAND2X1 U495 ( .A(n24), .B(si[1]), .Y(n355) );
  NAND2X1 U496 ( .A(n355), .B(n354), .Y(n356) );
  NAND2X1 U497 ( .A(n356), .B(n129), .Y(n358) );
  AOI22X1 U498 ( .A(intj[1]), .B(n53), .C(N497), .D(n644), .Y(n357) );
  NAND3X1 U499 ( .A(n359), .B(n358), .C(n357), .Y(n366) );
  NAND2X1 U500 ( .A(temp[1]), .B(n109), .Y(n361) );
  NAND2X1 U501 ( .A(n361), .B(n360), .Y(n365) );
  INVX2 U502 ( .A(faddr[1]), .Y(n363) );
  NAND2X1 U503 ( .A(n373), .B(inti[1]), .Y(n362) );
  OAI21X1 U504 ( .A(n650), .B(n363), .C(n362), .Y(n364) );
  NOR3X1 U505 ( .A(n366), .B(n365), .C(n364), .Y(n707) );
  NAND2X1 U506 ( .A(n48), .B(n367), .Y(n370) );
  NAND2X1 U507 ( .A(n129), .B(n1102), .Y(n369) );
  AOI22X1 U508 ( .A(intj[0]), .B(n53), .C(N496), .D(n644), .Y(n368) );
  NAND3X1 U509 ( .A(n370), .B(n369), .C(n368), .Y(n378) );
  NAND2X1 U510 ( .A(temp[0]), .B(n109), .Y(n372) );
  NAND2X1 U511 ( .A(n372), .B(n371), .Y(n377) );
  INVX2 U512 ( .A(faddr[0]), .Y(n375) );
  NAND2X1 U513 ( .A(n373), .B(inti[0]), .Y(n374) );
  OAI21X1 U514 ( .A(n650), .B(n375), .C(n374), .Y(n376) );
  NOR3X1 U515 ( .A(n378), .B(n377), .C(n376), .Y(n708) );
  NOR2X1 U516 ( .A(n684), .B(n52), .Y(n391) );
  INVX2 U517 ( .A(n387), .Y(n390) );
  AND2X2 U518 ( .A(n388), .B(n30), .Y(n389) );
  NAND3X1 U519 ( .A(n391), .B(n390), .C(n389), .Y(n397) );
  AOI21X1 U520 ( .A(fr_enable), .B(n397), .C(n17), .Y(n393) );
  INVX2 U521 ( .A(R_ENABLE), .Y(n392) );
  MUX2X1 U522 ( .B(n393), .A(n392), .S(n202), .Y(n717) );
  AND2X2 U523 ( .A(n681), .B(n30), .Y(n394) );
  NAND3X1 U524 ( .A(n36), .B(n1022), .C(n394), .Y(n402) );
  AOI21X1 U525 ( .A(fw_enable), .B(n401), .C(n402), .Y(n396) );
  INVX2 U526 ( .A(W_ENABLE), .Y(n395) );
  MUX2X1 U527 ( .B(n396), .A(n395), .S(n202), .Y(n718) );
  OAI21X1 U528 ( .A(n202), .B(n397), .C(fr_enable), .Y(n400) );
  NAND2X1 U529 ( .A(n17), .B(n207), .Y(n399) );
  NAND2X1 U530 ( .A(n400), .B(n399), .Y(n719) );
  OAI21X1 U531 ( .A(n202), .B(n401), .C(fw_enable), .Y(n404) );
  NAND2X1 U532 ( .A(n402), .B(n206), .Y(n403) );
  NAND2X1 U533 ( .A(n404), .B(n403), .Y(n720) );
  MUX2X1 U534 ( .B(nfaddr[0]), .A(ADDR[0]), .S(n201), .Y(n413) );
  INVX2 U535 ( .A(n413), .Y(n729) );
  MUX2X1 U536 ( .B(nfaddr[0]), .A(faddr[0]), .S(n201), .Y(n414) );
  INVX2 U537 ( .A(n414), .Y(n730) );
  MUX2X1 U538 ( .B(nfaddr[1]), .A(ADDR[1]), .S(n201), .Y(n415) );
  INVX2 U539 ( .A(n415), .Y(n731) );
  MUX2X1 U540 ( .B(nfaddr[1]), .A(faddr[1]), .S(n201), .Y(n416) );
  INVX2 U541 ( .A(n416), .Y(n732) );
  MUX2X1 U542 ( .B(nfaddr[2]), .A(ADDR[2]), .S(n201), .Y(n417) );
  INVX2 U543 ( .A(n417), .Y(n733) );
  MUX2X1 U544 ( .B(nfaddr[2]), .A(faddr[2]), .S(n201), .Y(n418) );
  INVX2 U545 ( .A(n418), .Y(n734) );
  MUX2X1 U546 ( .B(nfaddr[3]), .A(ADDR[3]), .S(n201), .Y(n419) );
  INVX2 U547 ( .A(n419), .Y(n735) );
  MUX2X1 U548 ( .B(nfaddr[3]), .A(faddr[3]), .S(n201), .Y(n420) );
  INVX2 U549 ( .A(n420), .Y(n736) );
  MUX2X1 U550 ( .B(nfaddr[4]), .A(ADDR[4]), .S(n201), .Y(n421) );
  INVX2 U551 ( .A(n421), .Y(n737) );
  MUX2X1 U552 ( .B(nfaddr[4]), .A(faddr[4]), .S(n201), .Y(n422) );
  INVX2 U553 ( .A(n422), .Y(n738) );
  MUX2X1 U554 ( .B(nfaddr[5]), .A(ADDR[5]), .S(n201), .Y(n423) );
  INVX2 U555 ( .A(n423), .Y(n739) );
  MUX2X1 U556 ( .B(nfaddr[5]), .A(faddr[5]), .S(n200), .Y(n424) );
  INVX2 U557 ( .A(n424), .Y(n740) );
  MUX2X1 U558 ( .B(nfaddr[6]), .A(ADDR[6]), .S(n200), .Y(n425) );
  INVX2 U559 ( .A(n425), .Y(n741) );
  MUX2X1 U560 ( .B(nfaddr[6]), .A(faddr[6]), .S(n200), .Y(n426) );
  INVX2 U561 ( .A(n426), .Y(n742) );
  MUX2X1 U562 ( .B(nfaddr[7]), .A(ADDR[7]), .S(n201), .Y(n427) );
  MUX2X1 U563 ( .B(nfaddr[7]), .A(faddr[7]), .S(n200), .Y(n428) );
  NAND3X1 U564 ( .A(n187), .B(n162), .C(n430), .Y(n647) );
  NOR2X1 U565 ( .A(n194), .B(n684), .Y(n433) );
  NAND2X1 U566 ( .A(n103), .B(currentProcessedData[7]), .Y(n439) );
  XOR2X1 U567 ( .A(delaydata[7]), .B(temp[7]), .Y(n435) );
  NAND2X1 U568 ( .A(n479), .B(n435), .Y(n438) );
  NAND2X1 U569 ( .A(BYTE[7]), .B(n480), .Y(n437) );
  INVX2 U570 ( .A(PROCESSED_DATA[7]), .Y(n440) );
  MUX2X1 U571 ( .B(n441), .A(n440), .S(n200), .Y(n745) );
  NAND2X1 U572 ( .A(n118), .B(currentProcessedData[6]), .Y(n445) );
  XOR2X1 U573 ( .A(delaydata[6]), .B(temp[6]), .Y(n442) );
  NAND2X1 U574 ( .A(n479), .B(n442), .Y(n444) );
  NAND2X1 U575 ( .A(BYTE[6]), .B(n480), .Y(n443) );
  NAND3X1 U576 ( .A(n445), .B(n444), .C(n443), .Y(nextProcessedData[6]) );
  INVX2 U577 ( .A(nextProcessedData[6]), .Y(n447) );
  INVX2 U578 ( .A(PROCESSED_DATA[6]), .Y(n446) );
  MUX2X1 U579 ( .B(n447), .A(n446), .S(n200), .Y(n747) );
  NAND2X1 U580 ( .A(n117), .B(currentProcessedData[5]), .Y(n451) );
  XOR2X1 U581 ( .A(delaydata[5]), .B(temp[5]), .Y(n448) );
  NAND2X1 U582 ( .A(n479), .B(n448), .Y(n450) );
  NAND2X1 U583 ( .A(BYTE[5]), .B(n480), .Y(n449) );
  NAND3X1 U584 ( .A(n451), .B(n450), .C(n449), .Y(nextProcessedData[5]) );
  INVX2 U585 ( .A(nextProcessedData[5]), .Y(n453) );
  INVX2 U586 ( .A(PROCESSED_DATA[5]), .Y(n452) );
  MUX2X1 U587 ( .B(n453), .A(n452), .S(n200), .Y(n749) );
  NAND2X1 U588 ( .A(n103), .B(currentProcessedData[4]), .Y(n457) );
  XOR2X1 U589 ( .A(delaydata[4]), .B(temp[4]), .Y(n454) );
  NAND2X1 U590 ( .A(n479), .B(n454), .Y(n456) );
  NAND2X1 U591 ( .A(BYTE[4]), .B(n480), .Y(n455) );
  NAND3X1 U592 ( .A(n457), .B(n456), .C(n455), .Y(nextProcessedData[4]) );
  INVX2 U593 ( .A(nextProcessedData[4]), .Y(n459) );
  INVX2 U594 ( .A(PROCESSED_DATA[4]), .Y(n458) );
  MUX2X1 U595 ( .B(n459), .A(n458), .S(n200), .Y(n751) );
  NAND2X1 U596 ( .A(n102), .B(currentProcessedData[3]), .Y(n463) );
  XOR2X1 U597 ( .A(delaydata[3]), .B(temp[3]), .Y(n460) );
  NAND2X1 U598 ( .A(n479), .B(n460), .Y(n462) );
  NAND2X1 U599 ( .A(BYTE[3]), .B(n480), .Y(n461) );
  NAND3X1 U600 ( .A(n463), .B(n462), .C(n461), .Y(nextProcessedData[3]) );
  INVX2 U601 ( .A(nextProcessedData[3]), .Y(n465) );
  INVX2 U602 ( .A(PROCESSED_DATA[3]), .Y(n464) );
  MUX2X1 U603 ( .B(n465), .A(n464), .S(n200), .Y(n753) );
  NAND2X1 U604 ( .A(n118), .B(currentProcessedData[2]), .Y(n469) );
  XOR2X1 U605 ( .A(delaydata[2]), .B(temp[2]), .Y(n466) );
  NAND2X1 U606 ( .A(n479), .B(n466), .Y(n468) );
  NAND2X1 U607 ( .A(BYTE[2]), .B(n480), .Y(n467) );
  NAND3X1 U608 ( .A(n469), .B(n468), .C(n467), .Y(nextProcessedData[2]) );
  INVX2 U609 ( .A(nextProcessedData[2]), .Y(n471) );
  INVX2 U610 ( .A(PROCESSED_DATA[2]), .Y(n470) );
  MUX2X1 U611 ( .B(n471), .A(n470), .S(n200), .Y(n755) );
  NAND2X1 U612 ( .A(n102), .B(currentProcessedData[1]), .Y(n475) );
  XOR2X1 U613 ( .A(delaydata[1]), .B(temp[1]), .Y(n472) );
  NAND2X1 U614 ( .A(n479), .B(n472), .Y(n474) );
  NAND2X1 U615 ( .A(BYTE[1]), .B(n480), .Y(n473) );
  INVX2 U616 ( .A(PROCESSED_DATA[1]), .Y(n476) );
  MUX2X1 U617 ( .B(n477), .A(n476), .S(n200), .Y(n757) );
  NAND2X1 U618 ( .A(n117), .B(currentProcessedData[0]), .Y(n483) );
  XOR2X1 U619 ( .A(delaydata[0]), .B(temp[0]), .Y(n478) );
  NAND2X1 U620 ( .A(n479), .B(n478), .Y(n482) );
  NAND2X1 U621 ( .A(BYTE[0]), .B(n480), .Y(n481) );
  INVX2 U622 ( .A(PROCESSED_DATA[0]), .Y(n484) );
  MUX2X1 U623 ( .B(n485), .A(n484), .S(n200), .Y(n759) );
  NOR2X1 U624 ( .A(n202), .B(n104), .Y(n489) );
  NAND2X1 U625 ( .A(n46), .B(n1060), .Y(n1073) );
  INVX2 U626 ( .A(n1073), .Y(n488) );
  NAND2X1 U627 ( .A(n488), .B(n133), .Y(n564) );
  NOR3X1 U628 ( .A(n75), .B(n156), .C(n132), .Y(n628) );
  AND2X2 U629 ( .A(n138), .B(n489), .Y(n507) );
  INVX2 U630 ( .A(N502), .Y(n491) );
  NAND3X1 U631 ( .A(n560), .B(n507), .C(n563), .Y(n504) );
  NAND2X1 U632 ( .A(inti[6]), .B(n504), .Y(n490) );
  OAI21X1 U633 ( .A(n44), .B(n491), .C(n490), .Y(n1125) );
  INVX2 U634 ( .A(N501), .Y(n493) );
  NAND2X1 U635 ( .A(inti[5]), .B(n504), .Y(n492) );
  OAI21X1 U636 ( .A(n44), .B(n493), .C(n492), .Y(n1124) );
  INVX2 U637 ( .A(N500), .Y(n495) );
  NAND2X1 U638 ( .A(inti[4]), .B(n504), .Y(n494) );
  OAI21X1 U639 ( .A(n43), .B(n495), .C(n494), .Y(n1123) );
  INVX2 U640 ( .A(N499), .Y(n497) );
  NAND2X1 U641 ( .A(inti[3]), .B(n504), .Y(n496) );
  OAI21X1 U642 ( .A(n33), .B(n497), .C(n496), .Y(n1122) );
  INVX2 U643 ( .A(N498), .Y(n499) );
  NAND2X1 U644 ( .A(inti[2]), .B(n504), .Y(n498) );
  OAI21X1 U645 ( .A(n43), .B(n499), .C(n498), .Y(n1121) );
  INVX2 U646 ( .A(N497), .Y(n501) );
  NAND2X1 U647 ( .A(inti[1]), .B(n504), .Y(n500) );
  OAI21X1 U648 ( .A(n44), .B(n501), .C(n500), .Y(n1120) );
  INVX2 U649 ( .A(N496), .Y(n503) );
  NAND2X1 U650 ( .A(inti[0]), .B(n504), .Y(n502) );
  OAI21X1 U651 ( .A(n43), .B(n503), .C(n502), .Y(n1119) );
  INVX2 U652 ( .A(N503), .Y(n506) );
  NAND2X1 U653 ( .A(inti[7]), .B(n504), .Y(n505) );
  OAI21X1 U654 ( .A(n33), .B(n506), .C(n505), .Y(n1126) );
  NAND3X1 U655 ( .A(keyi[2]), .B(n510), .C(n512), .Y(n508) );
  INVX2 U656 ( .A(n508), .Y(n550) );
  NAND3X1 U657 ( .A(keyi[2]), .B(keyi[0]), .C(n510), .Y(n509) );
  INVX2 U658 ( .A(n509), .Y(n549) );
  AOI22X1 U659 ( .A(\keyTable[4][7] ), .B(n550), .C(\keyTable[5][7] ), .D(n549), .Y(n518) );
  AOI22X1 U660 ( .A(\keyTable[6][7] ), .B(n164), .C(\keyTable[7][7] ), .D(n170), .Y(n517) );
  INVX2 U661 ( .A(\keyTable[3][7] ), .Y(n943) );
  NAND3X1 U662 ( .A(keyi[1]), .B(n511), .C(n512), .Y(n551) );
  INVX2 U663 ( .A(\keyTable[2][7] ), .Y(n927) );
  OAI22X1 U664 ( .A(n552), .B(n943), .C(n551), .D(n927), .Y(n515) );
  NAND3X1 U665 ( .A(keyi[0]), .B(n511), .C(n510), .Y(n554) );
  INVX2 U666 ( .A(\keyTable[1][7] ), .Y(n790) );
  NOR2X1 U667 ( .A(keyi[2]), .B(keyi[1]), .Y(n513) );
  NAND2X1 U668 ( .A(n513), .B(n512), .Y(n553) );
  INVX2 U670 ( .A(\keyTable[0][7] ), .Y(n788) );
  OAI22X1 U671 ( .A(n554), .B(n790), .C(n553), .D(n788), .Y(n514) );
  NOR2X1 U672 ( .A(n515), .B(n514), .Y(n516) );
  NAND3X1 U674 ( .A(n518), .B(n517), .C(n516), .Y(N472) );
  AOI22X1 U675 ( .A(\keyTable[4][6] ), .B(n550), .C(\keyTable[5][6] ), .D(n549), .Y(n523) );
  AOI22X1 U676 ( .A(\keyTable[6][6] ), .B(n164), .C(\keyTable[7][6] ), .D(n170), .Y(n522) );
  INVX2 U677 ( .A(\keyTable[3][6] ), .Y(n945) );
  INVX2 U678 ( .A(\keyTable[2][6] ), .Y(n929) );
  OAI22X1 U679 ( .A(n552), .B(n945), .C(n551), .D(n929), .Y(n520) );
  INVX2 U680 ( .A(\keyTable[1][6] ), .Y(n889) );
  INVX2 U681 ( .A(\keyTable[0][6] ), .Y(n887) );
  OAI22X1 U682 ( .A(n554), .B(n889), .C(n553), .D(n887), .Y(n519) );
  NOR2X1 U683 ( .A(n520), .B(n519), .Y(n521) );
  NAND3X1 U684 ( .A(n523), .B(n522), .C(n521), .Y(N473) );
  AOI22X1 U685 ( .A(\keyTable[4][5] ), .B(n550), .C(\keyTable[5][5] ), .D(n549), .Y(n528) );
  AOI22X1 U686 ( .A(\keyTable[6][5] ), .B(n164), .C(\keyTable[7][5] ), .D(n170), .Y(n527) );
  INVX2 U687 ( .A(\keyTable[3][5] ), .Y(n947) );
  INVX2 U688 ( .A(\keyTable[2][5] ), .Y(n931) );
  OAI22X1 U689 ( .A(n552), .B(n947), .C(n551), .D(n931), .Y(n525) );
  INVX2 U690 ( .A(\keyTable[1][5] ), .Y(n898) );
  INVX2 U691 ( .A(\keyTable[0][5] ), .Y(n885) );
  OAI22X1 U692 ( .A(n554), .B(n898), .C(n553), .D(n885), .Y(n524) );
  NOR2X1 U693 ( .A(n525), .B(n524), .Y(n526) );
  NAND3X1 U694 ( .A(n528), .B(n527), .C(n526), .Y(N474) );
  AOI22X1 U695 ( .A(\keyTable[4][4] ), .B(n550), .C(\keyTable[5][4] ), .D(n549), .Y(n533) );
  AOI22X1 U696 ( .A(\keyTable[6][4] ), .B(n164), .C(\keyTable[7][4] ), .D(n170), .Y(n532) );
  INVX2 U697 ( .A(\keyTable[3][4] ), .Y(n949) );
  INVX2 U698 ( .A(\keyTable[2][4] ), .Y(n933) );
  OAI22X1 U699 ( .A(n552), .B(n949), .C(n551), .D(n933), .Y(n530) );
  INVX2 U700 ( .A(\keyTable[1][4] ), .Y(n917) );
  INVX2 U701 ( .A(\keyTable[0][4] ), .Y(n883) );
  OAI22X1 U702 ( .A(n554), .B(n917), .C(n553), .D(n883), .Y(n529) );
  NOR2X1 U703 ( .A(n530), .B(n529), .Y(n531) );
  NAND3X1 U704 ( .A(n533), .B(n532), .C(n531), .Y(N475) );
  AOI22X1 U705 ( .A(\keyTable[4][3] ), .B(n550), .C(\keyTable[5][3] ), .D(n549), .Y(n538) );
  AOI22X1 U706 ( .A(\keyTable[6][3] ), .B(n164), .C(\keyTable[7][3] ), .D(n170), .Y(n537) );
  INVX2 U707 ( .A(\keyTable[3][3] ), .Y(n951) );
  INVX2 U708 ( .A(\keyTable[2][3] ), .Y(n935) );
  OAI22X1 U709 ( .A(n552), .B(n951), .C(n551), .D(n935), .Y(n535) );
  INVX2 U710 ( .A(\keyTable[1][3] ), .Y(n919) );
  INVX2 U711 ( .A(\keyTable[0][3] ), .Y(n870) );
  OAI22X1 U712 ( .A(n554), .B(n919), .C(n553), .D(n870), .Y(n534) );
  NOR2X1 U713 ( .A(n535), .B(n534), .Y(n536) );
  NAND3X1 U714 ( .A(n538), .B(n537), .C(n536), .Y(N476) );
  AOI22X1 U715 ( .A(\keyTable[4][2] ), .B(n550), .C(\keyTable[5][2] ), .D(n549), .Y(n543) );
  AOI22X1 U716 ( .A(\keyTable[6][2] ), .B(n164), .C(\keyTable[7][2] ), .D(n170), .Y(n542) );
  INVX2 U717 ( .A(\keyTable[3][2] ), .Y(n953) );
  INVX2 U718 ( .A(\keyTable[2][2] ), .Y(n937) );
  OAI22X1 U719 ( .A(n552), .B(n953), .C(n551), .D(n937), .Y(n540) );
  INVX2 U720 ( .A(\keyTable[1][2] ), .Y(n921) );
  INVX2 U721 ( .A(\keyTable[0][2] ), .Y(n868) );
  OAI22X1 U722 ( .A(n554), .B(n921), .C(n553), .D(n868), .Y(n539) );
  NOR2X1 U723 ( .A(n540), .B(n539), .Y(n541) );
  NAND3X1 U724 ( .A(n543), .B(n542), .C(n541), .Y(N477) );
  AOI22X1 U725 ( .A(\keyTable[4][1] ), .B(n550), .C(\keyTable[5][1] ), .D(n549), .Y(n548) );
  AOI22X1 U726 ( .A(\keyTable[6][1] ), .B(n164), .C(\keyTable[7][1] ), .D(n170), .Y(n547) );
  INVX2 U727 ( .A(\keyTable[3][1] ), .Y(n955) );
  INVX2 U728 ( .A(\keyTable[2][1] ), .Y(n939) );
  OAI22X1 U729 ( .A(n552), .B(n955), .C(n551), .D(n939), .Y(n545) );
  INVX2 U730 ( .A(\keyTable[1][1] ), .Y(n923) );
  INVX2 U731 ( .A(\keyTable[0][1] ), .Y(n866) );
  OAI22X1 U732 ( .A(n554), .B(n923), .C(n553), .D(n866), .Y(n544) );
  NOR2X1 U733 ( .A(n545), .B(n544), .Y(n546) );
  NAND3X1 U734 ( .A(n548), .B(n547), .C(n546), .Y(N478) );
  AOI22X1 U735 ( .A(\keyTable[4][0] ), .B(n550), .C(\keyTable[5][0] ), .D(n549), .Y(n559) );
  AOI22X1 U736 ( .A(\keyTable[6][0] ), .B(n164), .C(\keyTable[7][0] ), .D(n170), .Y(n558) );
  INVX2 U737 ( .A(\keyTable[3][0] ), .Y(n957) );
  INVX2 U738 ( .A(\keyTable[2][0] ), .Y(n941) );
  OAI22X1 U739 ( .A(n552), .B(n957), .C(n551), .D(n941), .Y(n556) );
  INVX2 U740 ( .A(\keyTable[1][0] ), .Y(n925) );
  INVX2 U741 ( .A(\keyTable[0][0] ), .Y(n864) );
  OAI22X1 U742 ( .A(n554), .B(n925), .C(n553), .D(n864), .Y(n555) );
  NOR2X1 U743 ( .A(n556), .B(n555), .Y(n557) );
  NAND3X1 U744 ( .A(n559), .B(n558), .C(n557), .Y(N479) );
  NAND3X1 U745 ( .A(n560), .B(n7), .C(n70), .Y(n561) );
  AND2X2 U746 ( .A(n566), .B(n22), .Y(n590) );
  NAND2X1 U747 ( .A(n590), .B(n54), .Y(n582) );
  INVX2 U748 ( .A(n582), .Y(n573) );
  INVX2 U749 ( .A(n48), .Y(n568) );
  INVX2 U750 ( .A(n1090), .Y(n587) );
  NAND2X1 U751 ( .A(N480), .B(n587), .Y(n567) );
  OAI21X1 U752 ( .A(n573), .B(n568), .C(n567), .Y(n891) );
  INVX2 U753 ( .A(sj[1]), .Y(n570) );
  NAND2X1 U754 ( .A(N481), .B(n587), .Y(n569) );
  OAI21X1 U755 ( .A(n573), .B(n570), .C(n569), .Y(n892) );
  NAND2X1 U756 ( .A(N482), .B(n587), .Y(n571) );
  OAI21X1 U757 ( .A(n573), .B(n572), .C(n571), .Y(n893) );
  NAND2X1 U758 ( .A(sj[3]), .B(n582), .Y(n575) );
  NAND2X1 U759 ( .A(N483), .B(n587), .Y(n574) );
  NAND2X1 U760 ( .A(n575), .B(n574), .Y(n894) );
  NAND2X1 U761 ( .A(sj[4]), .B(n582), .Y(n577) );
  NAND2X1 U762 ( .A(N484), .B(n587), .Y(n576) );
  NAND2X1 U763 ( .A(n577), .B(n576), .Y(n895) );
  NAND2X1 U764 ( .A(sj[5]), .B(n582), .Y(n579) );
  NAND2X1 U765 ( .A(N485), .B(n587), .Y(n578) );
  NAND2X1 U766 ( .A(n579), .B(n578), .Y(n896) );
  NAND2X1 U767 ( .A(sj[6]), .B(n582), .Y(n581) );
  NAND2X1 U768 ( .A(N486), .B(n587), .Y(n580) );
  NAND2X1 U769 ( .A(n581), .B(n580), .Y(n897) );
  NAND2X1 U770 ( .A(sj[7]), .B(n582), .Y(n584) );
  INVX2 U771 ( .A(N487), .Y(n583) );
  AOI22X1 U772 ( .A(n584), .B(n1090), .C(n584), .D(n583), .Y(n1099) );
  NAND2X1 U773 ( .A(n106), .B(n205), .Y(n586) );
  NOR2X1 U774 ( .A(n587), .B(n586), .Y(n591) );
  INVX2 U775 ( .A(N518), .Y(n593) );
  NAND2X1 U776 ( .A(intj[6]), .B(n55), .Y(n592) );
  OAI21X1 U777 ( .A(n608), .B(n593), .C(n592), .Y(n876) );
  INVX2 U778 ( .A(N517), .Y(n595) );
  NAND2X1 U779 ( .A(intj[5]), .B(n55), .Y(n594) );
  OAI21X1 U780 ( .A(n608), .B(n595), .C(n594), .Y(n877) );
  INVX2 U781 ( .A(N516), .Y(n597) );
  NAND2X1 U782 ( .A(intj[4]), .B(n55), .Y(n596) );
  OAI21X1 U783 ( .A(n608), .B(n597), .C(n596), .Y(n878) );
  INVX2 U784 ( .A(N515), .Y(n599) );
  NAND2X1 U785 ( .A(intj[3]), .B(n55), .Y(n598) );
  OAI21X1 U786 ( .A(n608), .B(n599), .C(n598), .Y(n879) );
  INVX2 U787 ( .A(N514), .Y(n601) );
  NAND2X1 U788 ( .A(intj[2]), .B(n55), .Y(n600) );
  OAI21X1 U789 ( .A(n608), .B(n601), .C(n600), .Y(n880) );
  INVX2 U790 ( .A(N513), .Y(n603) );
  NAND2X1 U791 ( .A(intj[1]), .B(n55), .Y(n602) );
  OAI21X1 U792 ( .A(n608), .B(n603), .C(n602), .Y(n881) );
  INVX2 U793 ( .A(N512), .Y(n605) );
  NAND2X1 U794 ( .A(intj[0]), .B(n55), .Y(n604) );
  OAI21X1 U795 ( .A(n608), .B(n605), .C(n604), .Y(n882) );
  INVX2 U796 ( .A(N519), .Y(n607) );
  NAND2X1 U797 ( .A(intj[7]), .B(n55), .Y(n606) );
  OAI21X1 U798 ( .A(n608), .B(n607), .C(n606), .Y(n875) );
  INVX2 U799 ( .A(delaydata[6]), .Y(n610) );
  INVX2 U800 ( .A(BYTE[6]), .Y(n609) );
  MUX2X1 U801 ( .B(n610), .A(n609), .S(n191), .Y(n1112) );
  INVX2 U802 ( .A(delaydata[5]), .Y(n612) );
  INVX2 U803 ( .A(BYTE[5]), .Y(n611) );
  MUX2X1 U804 ( .B(n612), .A(n611), .S(n192), .Y(n1113) );
  INVX2 U805 ( .A(delaydata[4]), .Y(n614) );
  INVX2 U806 ( .A(BYTE[4]), .Y(n613) );
  MUX2X1 U807 ( .B(n614), .A(n613), .S(n191), .Y(n1114) );
  INVX2 U808 ( .A(delaydata[3]), .Y(n616) );
  INVX2 U809 ( .A(BYTE[3]), .Y(n615) );
  MUX2X1 U810 ( .B(n616), .A(n615), .S(n192), .Y(n1115) );
  INVX2 U811 ( .A(delaydata[2]), .Y(n618) );
  INVX2 U812 ( .A(BYTE[2]), .Y(n617) );
  MUX2X1 U813 ( .B(n618), .A(n617), .S(n191), .Y(n1116) );
  INVX2 U814 ( .A(delaydata[1]), .Y(n620) );
  INVX2 U815 ( .A(BYTE[1]), .Y(n619) );
  MUX2X1 U816 ( .B(n620), .A(n619), .S(n192), .Y(n1117) );
  INVX2 U817 ( .A(delaydata[0]), .Y(n622) );
  INVX2 U818 ( .A(BYTE[0]), .Y(n621) );
  MUX2X1 U819 ( .B(n622), .A(n621), .S(n191), .Y(n1118) );
  INVX2 U820 ( .A(delaydata[7]), .Y(n624) );
  INVX2 U821 ( .A(BYTE[7]), .Y(n623) );
  MUX2X1 U822 ( .B(n624), .A(n623), .S(n192), .Y(n1111) );
  NAND3X1 U823 ( .A(si[3]), .B(si[2]), .C(si[6]), .Y(n626) );
  NAND2X1 U824 ( .A(n588), .B(si[7]), .Y(n625) );
  NOR2X1 U825 ( .A(n626), .B(n625), .Y(n627) );
  NAND2X1 U826 ( .A(n627), .B(n589), .Y(n1055) );
  NAND2X1 U827 ( .A(N431), .B(n166), .Y(n631) );
  NAND2X1 U828 ( .A(n629), .B(n628), .Y(n634) );
  NAND2X1 U829 ( .A(si[7]), .B(n634), .Y(n630) );
  NAND2X1 U830 ( .A(n631), .B(n630), .Y(n900) );
  NAND2X1 U831 ( .A(N430), .B(n166), .Y(n633) );
  NAND2X1 U832 ( .A(si[6]), .B(n634), .Y(n632) );
  NAND2X1 U833 ( .A(n633), .B(n632), .Y(n901) );
  INVX2 U834 ( .A(n634), .Y(n643) );
  NAND2X1 U835 ( .A(N429), .B(n166), .Y(n635) );
  OAI21X1 U836 ( .A(n1105), .B(n643), .C(n635), .Y(n902) );
  NAND2X1 U837 ( .A(N428), .B(n166), .Y(n636) );
  OAI21X1 U838 ( .A(n1104), .B(n643), .C(n636), .Y(n903) );
  NAND2X1 U839 ( .A(N427), .B(n166), .Y(n637) );
  OAI21X1 U840 ( .A(n643), .B(n638), .C(n637), .Y(n904) );
  NAND2X1 U841 ( .A(N426), .B(n166), .Y(n639) );
  OAI21X1 U842 ( .A(n643), .B(n640), .C(n639), .Y(n905) );
  NAND2X1 U843 ( .A(N425), .B(n166), .Y(n641) );
  OAI21X1 U844 ( .A(n1103), .B(n643), .C(n641), .Y(n906) );
  NAND2X1 U845 ( .A(N424), .B(n166), .Y(n642) );
  OAI21X1 U846 ( .A(n1102), .B(n643), .C(n642), .Y(n907) );
  NOR2X1 U847 ( .A(n645), .B(n644), .Y(n651) );
  NAND2X1 U848 ( .A(n91), .B(n203), .Y(n648) );
  NAND3X1 U849 ( .A(n651), .B(n71), .C(n649), .Y(n674) );
  NAND2X1 U850 ( .A(temp[6]), .B(n196), .Y(n654) );
  NAND3X1 U851 ( .A(DATA_IN[6]), .B(n3), .C(n675), .Y(n653) );
  NAND3X1 U852 ( .A(N526), .B(n676), .C(n675), .Y(n652) );
  NAND3X1 U853 ( .A(n654), .B(n652), .C(n653), .Y(n857) );
  NAND2X1 U854 ( .A(temp[5]), .B(n196), .Y(n657) );
  NAND3X1 U855 ( .A(DATA_IN[5]), .B(n3), .C(n675), .Y(n656) );
  NAND3X1 U856 ( .A(N525), .B(n676), .C(n675), .Y(n655) );
  NAND3X1 U857 ( .A(n657), .B(n655), .C(n656), .Y(n858) );
  NAND2X1 U858 ( .A(temp[4]), .B(n196), .Y(n660) );
  NAND3X1 U859 ( .A(DATA_IN[4]), .B(n3), .C(n675), .Y(n659) );
  NAND3X1 U860 ( .A(N524), .B(n676), .C(n675), .Y(n658) );
  NAND3X1 U861 ( .A(n660), .B(n658), .C(n659), .Y(n859) );
  NAND2X1 U862 ( .A(temp[3]), .B(n196), .Y(n663) );
  NAND3X1 U863 ( .A(DATA_IN[3]), .B(n3), .C(n675), .Y(n662) );
  NAND3X1 U864 ( .A(N523), .B(n676), .C(n151), .Y(n661) );
  NAND3X1 U865 ( .A(n663), .B(n661), .C(n662), .Y(n860) );
  NAND2X1 U866 ( .A(temp[2]), .B(n196), .Y(n666) );
  NAND3X1 U867 ( .A(DATA_IN[2]), .B(n3), .C(n675), .Y(n665) );
  NAND3X1 U868 ( .A(N522), .B(n676), .C(n151), .Y(n664) );
  NAND3X1 U869 ( .A(n666), .B(n664), .C(n665), .Y(n861) );
  NAND2X1 U870 ( .A(temp[1]), .B(n196), .Y(n669) );
  NAND3X1 U871 ( .A(DATA_IN[1]), .B(n3), .C(n675), .Y(n668) );
  NAND3X1 U872 ( .A(N521), .B(n676), .C(n675), .Y(n667) );
  NAND3X1 U873 ( .A(n669), .B(n667), .C(n668), .Y(n862) );
  NAND2X1 U874 ( .A(temp[0]), .B(n196), .Y(n673) );
  NAND3X1 U875 ( .A(DATA_IN[0]), .B(n3), .C(n151), .Y(n672) );
  NAND3X1 U876 ( .A(N520), .B(n676), .C(n675), .Y(n671) );
  NAND3X1 U877 ( .A(n673), .B(n672), .C(n671), .Y(n863) );
  NAND2X1 U878 ( .A(temp[7]), .B(n196), .Y(n679) );
  NAND3X1 U879 ( .A(DATA_IN[7]), .B(n3), .C(n675), .Y(n678) );
  NAND3X1 U880 ( .A(N527), .B(n676), .C(n151), .Y(n677) );
  NAND3X1 U881 ( .A(n679), .B(n677), .C(n678), .Y(n856) );
  NAND3X1 U882 ( .A(n682), .B(n60), .C(n57), .Y(n785) );
  NAND2X1 U883 ( .A(n684), .B(n141), .Y(n1098) );
  INVX2 U884 ( .A(N413), .Y(n686) );
  NAND2X1 U885 ( .A(prefillCounter[6]), .B(n149), .Y(n685) );
  OAI21X1 U886 ( .A(n68), .B(n686), .C(n685), .Y(n908) );
  INVX2 U887 ( .A(N412), .Y(n688) );
  NAND2X1 U888 ( .A(n149), .B(prefillCounter[5]), .Y(n687) );
  OAI21X1 U889 ( .A(n68), .B(n688), .C(n687), .Y(n909) );
  INVX2 U890 ( .A(N411), .Y(n690) );
  NAND2X1 U891 ( .A(prefillCounter[4]), .B(n149), .Y(n689) );
  OAI21X1 U892 ( .A(n68), .B(n690), .C(n689), .Y(n910) );
  INVX2 U893 ( .A(N410), .Y(n701) );
  NAND2X1 U894 ( .A(prefillCounter[3]), .B(n149), .Y(n692) );
  OAI21X1 U895 ( .A(n68), .B(n701), .C(n692), .Y(n911) );
  INVX2 U896 ( .A(N409), .Y(n766) );
  NAND2X1 U897 ( .A(prefillCounter[2]), .B(n149), .Y(n765) );
  OAI21X1 U898 ( .A(n1098), .B(n766), .C(n765), .Y(n912) );
  INVX2 U899 ( .A(N408), .Y(n770) );
  NAND2X1 U900 ( .A(prefillCounter[1]), .B(n149), .Y(n769) );
  OAI21X1 U901 ( .A(n1098), .B(n770), .C(n769), .Y(n913) );
  INVX2 U914 ( .A(N414), .Y(n784) );
  NAND2X1 U915 ( .A(prefillCounter[7]), .B(n149), .Y(n783) );
  OAI21X1 U918 ( .A(n1098), .B(n784), .C(n783), .Y(n914) );
  INVX2 U919 ( .A(KEY[7]), .Y(n787) );
  NOR2X1 U932 ( .A(n47), .B(n785), .Y(n786) );
  MUX2X1 U933 ( .B(n788), .A(n787), .S(n137), .Y(n855) );
  INVX2 U934 ( .A(KEY[15]), .Y(n789) );
  MUX2X1 U935 ( .B(n790), .A(n789), .S(n78), .Y(n854) );
  INVX2 U936 ( .A(KEY[0]), .Y(n791) );
  MUX2X1 U937 ( .B(n864), .A(n791), .S(n137), .Y(n853) );
  INVX2 U938 ( .A(KEY[1]), .Y(n865) );
  MUX2X1 U939 ( .B(n866), .A(n865), .S(n82), .Y(n852) );
  INVX2 U940 ( .A(KEY[2]), .Y(n867) );
  MUX2X1 U941 ( .B(n868), .A(n867), .S(n80), .Y(n851) );
  INVX2 U942 ( .A(KEY[3]), .Y(n869) );
  MUX2X1 U943 ( .B(n870), .A(n869), .S(n137), .Y(n850) );
  INVX2 U944 ( .A(KEY[4]), .Y(n871) );
  MUX2X1 U945 ( .B(n883), .A(n871), .S(n137), .Y(n849) );
  INVX2 U946 ( .A(KEY[5]), .Y(n884) );
  MUX2X1 U947 ( .B(n885), .A(n884), .S(n137), .Y(n848) );
  INVX2 U948 ( .A(KEY[6]), .Y(n886) );
  MUX2X1 U949 ( .B(n887), .A(n886), .S(n137), .Y(n847) );
  INVX2 U950 ( .A(KEY[14]), .Y(n888) );
  MUX2X1 U951 ( .B(n889), .A(n888), .S(n78), .Y(n846) );
  INVX2 U952 ( .A(KEY[13]), .Y(n890) );
  MUX2X1 U953 ( .B(n898), .A(n890), .S(n137), .Y(n845) );
  INVX2 U954 ( .A(KEY[12]), .Y(n916) );
  MUX2X1 U955 ( .B(n917), .A(n916), .S(n77), .Y(n844) );
  INVX2 U956 ( .A(KEY[11]), .Y(n918) );
  MUX2X1 U957 ( .B(n919), .A(n918), .S(n77), .Y(n843) );
  INVX2 U958 ( .A(KEY[10]), .Y(n920) );
  MUX2X1 U959 ( .B(n921), .A(n920), .S(n77), .Y(n842) );
  INVX2 U960 ( .A(KEY[9]), .Y(n922) );
  MUX2X1 U961 ( .B(n923), .A(n922), .S(n78), .Y(n841) );
  INVX2 U962 ( .A(KEY[8]), .Y(n924) );
  MUX2X1 U963 ( .B(n925), .A(n924), .S(n78), .Y(n840) );
  INVX2 U964 ( .A(KEY[23]), .Y(n926) );
  MUX2X1 U965 ( .B(n927), .A(n926), .S(n80), .Y(n839) );
  INVX2 U966 ( .A(KEY[22]), .Y(n928) );
  MUX2X1 U967 ( .B(n929), .A(n928), .S(n143), .Y(n838) );
  INVX2 U968 ( .A(KEY[21]), .Y(n930) );
  MUX2X1 U969 ( .B(n931), .A(n930), .S(n137), .Y(n837) );
  INVX2 U970 ( .A(KEY[20]), .Y(n932) );
  MUX2X1 U971 ( .B(n933), .A(n932), .S(n137), .Y(n836) );
  INVX2 U972 ( .A(KEY[19]), .Y(n934) );
  MUX2X1 U973 ( .B(n935), .A(n934), .S(n137), .Y(n835) );
  INVX2 U974 ( .A(KEY[18]), .Y(n936) );
  MUX2X1 U975 ( .B(n937), .A(n936), .S(n143), .Y(n834) );
  INVX2 U976 ( .A(KEY[17]), .Y(n938) );
  MUX2X1 U977 ( .B(n939), .A(n938), .S(n82), .Y(n833) );
  INVX2 U978 ( .A(KEY[16]), .Y(n940) );
  MUX2X1 U979 ( .B(n941), .A(n940), .S(n137), .Y(n832) );
  INVX2 U980 ( .A(KEY[31]), .Y(n942) );
  MUX2X1 U981 ( .B(n943), .A(n942), .S(n80), .Y(n831) );
  INVX2 U982 ( .A(KEY[30]), .Y(n944) );
  MUX2X1 U983 ( .B(n945), .A(n944), .S(n82), .Y(n830) );
  INVX2 U984 ( .A(KEY[29]), .Y(n946) );
  MUX2X1 U985 ( .B(n947), .A(n946), .S(n82), .Y(n829) );
  INVX2 U986 ( .A(KEY[28]), .Y(n948) );
  MUX2X1 U987 ( .B(n949), .A(n948), .S(n80), .Y(n828) );
  INVX2 U988 ( .A(KEY[27]), .Y(n950) );
  MUX2X1 U989 ( .B(n951), .A(n950), .S(n137), .Y(n827) );
  INVX2 U990 ( .A(KEY[26]), .Y(n952) );
  MUX2X1 U991 ( .B(n953), .A(n952), .S(n143), .Y(n826) );
  INVX2 U992 ( .A(KEY[25]), .Y(n954) );
  MUX2X1 U993 ( .B(n955), .A(n954), .S(n137), .Y(n825) );
  INVX2 U994 ( .A(KEY[24]), .Y(n956) );
  MUX2X1 U995 ( .B(n957), .A(n956), .S(n143), .Y(n824) );
  INVX2 U996 ( .A(\keyTable[4][7] ), .Y(n959) );
  INVX2 U997 ( .A(KEY[39]), .Y(n958) );
  MUX2X1 U998 ( .B(n959), .A(n958), .S(n137), .Y(n823) );
  INVX2 U999 ( .A(\keyTable[4][6] ), .Y(n961) );
  INVX2 U1000 ( .A(KEY[38]), .Y(n960) );
  MUX2X1 U1001 ( .B(n961), .A(n960), .S(n77), .Y(n822) );
  INVX2 U1002 ( .A(\keyTable[4][5] ), .Y(n963) );
  INVX2 U1003 ( .A(KEY[37]), .Y(n962) );
  MUX2X1 U1004 ( .B(n963), .A(n962), .S(n78), .Y(n821) );
  INVX2 U1005 ( .A(\keyTable[4][4] ), .Y(n965) );
  INVX2 U1006 ( .A(KEY[36]), .Y(n964) );
  MUX2X1 U1007 ( .B(n965), .A(n964), .S(n78), .Y(n820) );
  INVX2 U1008 ( .A(\keyTable[4][3] ), .Y(n967) );
  INVX2 U1009 ( .A(KEY[35]), .Y(n966) );
  MUX2X1 U1010 ( .B(n967), .A(n966), .S(n78), .Y(n819) );
  INVX2 U1011 ( .A(\keyTable[4][2] ), .Y(n969) );
  INVX2 U1012 ( .A(KEY[34]), .Y(n968) );
  MUX2X1 U1013 ( .B(n969), .A(n968), .S(n80), .Y(n818) );
  INVX2 U1014 ( .A(\keyTable[4][1] ), .Y(n971) );
  INVX2 U1015 ( .A(KEY[33]), .Y(n970) );
  MUX2X1 U1016 ( .B(n971), .A(n970), .S(n78), .Y(n817) );
  INVX2 U1017 ( .A(\keyTable[4][0] ), .Y(n973) );
  INVX2 U1018 ( .A(KEY[32]), .Y(n972) );
  MUX2X1 U1019 ( .B(n973), .A(n972), .S(n77), .Y(n816) );
  INVX2 U1020 ( .A(\keyTable[5][7] ), .Y(n975) );
  INVX2 U1021 ( .A(KEY[47]), .Y(n974) );
  MUX2X1 U1022 ( .B(n975), .A(n974), .S(n143), .Y(n815) );
  INVX2 U1023 ( .A(\keyTable[5][6] ), .Y(n977) );
  INVX2 U1024 ( .A(KEY[46]), .Y(n976) );
  MUX2X1 U1025 ( .B(n977), .A(n976), .S(n143), .Y(n814) );
  INVX2 U1026 ( .A(\keyTable[5][5] ), .Y(n979) );
  INVX2 U1027 ( .A(KEY[45]), .Y(n978) );
  MUX2X1 U1028 ( .B(n979), .A(n978), .S(n77), .Y(n813) );
  INVX2 U1029 ( .A(\keyTable[5][4] ), .Y(n981) );
  INVX2 U1030 ( .A(KEY[44]), .Y(n980) );
  MUX2X1 U1031 ( .B(n981), .A(n980), .S(n80), .Y(n812) );
  INVX2 U1032 ( .A(\keyTable[5][3] ), .Y(n983) );
  INVX2 U1033 ( .A(KEY[43]), .Y(n982) );
  MUX2X1 U1034 ( .B(n983), .A(n982), .S(n78), .Y(n811) );
  INVX2 U1035 ( .A(\keyTable[5][2] ), .Y(n985) );
  INVX2 U1036 ( .A(KEY[42]), .Y(n984) );
  MUX2X1 U1037 ( .B(n985), .A(n984), .S(n143), .Y(n810) );
  INVX2 U1038 ( .A(\keyTable[5][1] ), .Y(n987) );
  INVX2 U1039 ( .A(KEY[41]), .Y(n986) );
  MUX2X1 U1040 ( .B(n987), .A(n986), .S(n78), .Y(n809) );
  INVX2 U1041 ( .A(\keyTable[5][0] ), .Y(n989) );
  INVX2 U1042 ( .A(KEY[40]), .Y(n988) );
  MUX2X1 U1043 ( .B(n989), .A(n988), .S(n77), .Y(n808) );
  INVX2 U1044 ( .A(\keyTable[6][7] ), .Y(n991) );
  INVX2 U1045 ( .A(KEY[55]), .Y(n990) );
  MUX2X1 U1046 ( .B(n991), .A(n990), .S(n77), .Y(n807) );
  INVX2 U1047 ( .A(\keyTable[6][6] ), .Y(n993) );
  INVX2 U1048 ( .A(KEY[54]), .Y(n992) );
  MUX2X1 U1049 ( .B(n993), .A(n992), .S(n78), .Y(n806) );
  INVX2 U1050 ( .A(\keyTable[6][5] ), .Y(n995) );
  INVX2 U1051 ( .A(KEY[53]), .Y(n994) );
  MUX2X1 U1052 ( .B(n995), .A(n994), .S(n80), .Y(n805) );
  INVX2 U1053 ( .A(\keyTable[6][4] ), .Y(n997) );
  INVX2 U1054 ( .A(KEY[52]), .Y(n996) );
  MUX2X1 U1055 ( .B(n997), .A(n996), .S(n82), .Y(n804) );
  INVX2 U1056 ( .A(\keyTable[6][3] ), .Y(n999) );
  INVX2 U1057 ( .A(KEY[51]), .Y(n998) );
  MUX2X1 U1058 ( .B(n999), .A(n998), .S(n77), .Y(n803) );
  INVX2 U1059 ( .A(\keyTable[6][2] ), .Y(n1001) );
  INVX2 U1060 ( .A(KEY[50]), .Y(n1000) );
  MUX2X1 U1061 ( .B(n1001), .A(n1000), .S(n82), .Y(n802) );
  INVX2 U1062 ( .A(\keyTable[6][1] ), .Y(n1003) );
  INVX2 U1063 ( .A(KEY[49]), .Y(n1002) );
  MUX2X1 U1064 ( .B(n1003), .A(n1002), .S(n77), .Y(n801) );
  INVX2 U1065 ( .A(\keyTable[6][0] ), .Y(n1005) );
  INVX2 U1066 ( .A(KEY[48]), .Y(n1004) );
  MUX2X1 U1067 ( .B(n1005), .A(n1004), .S(n82), .Y(n800) );
  INVX2 U1068 ( .A(\keyTable[7][7] ), .Y(n1007) );
  INVX2 U1069 ( .A(KEY[63]), .Y(n1006) );
  MUX2X1 U1070 ( .B(n1007), .A(n1006), .S(n82), .Y(n799) );
  INVX2 U1071 ( .A(\keyTable[7][6] ), .Y(n1009) );
  INVX2 U1072 ( .A(KEY[62]), .Y(n1008) );
  MUX2X1 U1073 ( .B(n1009), .A(n1008), .S(n80), .Y(n798) );
  INVX2 U1074 ( .A(\keyTable[7][5] ), .Y(n1011) );
  INVX2 U1075 ( .A(KEY[61]), .Y(n1010) );
  MUX2X1 U1076 ( .B(n1011), .A(n1010), .S(n77), .Y(n797) );
  INVX2 U1077 ( .A(\keyTable[7][4] ), .Y(n1013) );
  INVX2 U1078 ( .A(KEY[60]), .Y(n1012) );
  MUX2X1 U1079 ( .B(n1013), .A(n1012), .S(n143), .Y(n796) );
  INVX2 U1080 ( .A(\keyTable[7][3] ), .Y(n1015) );
  INVX2 U1081 ( .A(KEY[59]), .Y(n1014) );
  MUX2X1 U1082 ( .B(n1015), .A(n1014), .S(n78), .Y(n795) );
  INVX2 U1083 ( .A(\keyTable[7][2] ), .Y(n1017) );
  INVX2 U1084 ( .A(KEY[58]), .Y(n1016) );
  MUX2X1 U1085 ( .B(n1017), .A(n1016), .S(n77), .Y(n794) );
  INVX2 U1086 ( .A(\keyTable[7][1] ), .Y(n1019) );
  INVX2 U1087 ( .A(KEY[57]), .Y(n1018) );
  MUX2X1 U1088 ( .B(n1019), .A(n1018), .S(n77), .Y(n793) );
  INVX2 U1089 ( .A(\keyTable[7][0] ), .Y(n1021) );
  INVX2 U1090 ( .A(KEY[56]), .Y(n1020) );
  MUX2X1 U1091 ( .B(n1021), .A(n1020), .S(n78), .Y(n792) );
  INVX2 U1092 ( .A(extratemp[0]), .Y(n1029) );
  INVX2 U1093 ( .A(DATA_IN[0]), .Y(n1028) );
  NAND2X1 U1094 ( .A(n28), .B(n134), .Y(n1023) );
  NAND2X1 U1095 ( .A(n1023), .B(n1022), .Y(n1024) );
  MUX2X1 U1096 ( .B(n1029), .A(n1028), .S(n1042), .Y(n1127) );
  INVX2 U1097 ( .A(extratemp[1]), .Y(n1031) );
  INVX2 U1098 ( .A(DATA_IN[1]), .Y(n1030) );
  MUX2X1 U1099 ( .B(n1031), .A(n1030), .S(n1042), .Y(n1128) );
  INVX2 U1100 ( .A(extratemp[2]), .Y(n1033) );
  INVX2 U1101 ( .A(DATA_IN[2]), .Y(n1032) );
  MUX2X1 U1102 ( .B(n1033), .A(n1032), .S(n1042), .Y(n1129) );
  INVX2 U1103 ( .A(extratemp[3]), .Y(n1035) );
  INVX2 U1104 ( .A(DATA_IN[3]), .Y(n1034) );
  MUX2X1 U1105 ( .B(n1035), .A(n1034), .S(n1042), .Y(n1130) );
  INVX2 U1106 ( .A(extratemp[4]), .Y(n1037) );
  INVX2 U1107 ( .A(DATA_IN[4]), .Y(n1036) );
  MUX2X1 U1108 ( .B(n1037), .A(n1036), .S(n1042), .Y(n1131) );
  INVX2 U1109 ( .A(extratemp[5]), .Y(n1039) );
  INVX2 U1110 ( .A(DATA_IN[5]), .Y(n1038) );
  MUX2X1 U1111 ( .B(n1039), .A(n1038), .S(n1042), .Y(n1132) );
  INVX2 U1112 ( .A(extratemp[6]), .Y(n1041) );
  INVX2 U1113 ( .A(DATA_IN[6]), .Y(n1040) );
  MUX2X1 U1114 ( .B(n1041), .A(n1040), .S(n1042), .Y(n1133) );
  INVX2 U1115 ( .A(extratemp[7]), .Y(n1044) );
  INVX2 U1116 ( .A(DATA_IN[7]), .Y(n1043) );
  MUX2X1 U1117 ( .B(n1044), .A(n1043), .S(n1042), .Y(n1134) );
  AOI21X1 U1118 ( .A(n12), .B(n177), .C(n1135), .Y(n1053) );
  NAND2X1 U1119 ( .A(permuteComplete), .B(n1046), .Y(n1047) );
  NAND3X1 U1120 ( .A(n147), .B(n70), .C(n1047), .Y(n1091) );
  INVX2 U1121 ( .A(n1091), .Y(n1052) );
  OAI21X1 U1122 ( .A(n105), .B(n107), .C(n119), .Y(n1049) );
  AOI22X1 U1123 ( .A(n1106), .B(n1050), .C(n134), .D(n1049), .Y(n1051) );
  NAND3X1 U1124 ( .A(n1053), .B(n1052), .C(n1051), .Y(nextState[3]) );
  OAI21X1 U1125 ( .A(n1055), .B(n1057), .C(n1054), .Y(n1056) );
  NAND2X1 U1126 ( .A(n88), .B(n1056), .Y(n1059) );
  NAND2X1 U1127 ( .A(n1057), .B(permuteComplete), .Y(n1058) );
  NAND2X1 U1128 ( .A(n1059), .B(n1058), .Y(n899) );
  NAND3X1 U1129 ( .A(n1108), .B(BYTE_READY), .C(n1085), .Y(n1063) );
  NAND2X1 U1130 ( .A(n128), .B(n1084), .Y(n1062) );
  NAND2X1 U1131 ( .A(n178), .B(n1071), .Y(n1061) );
  NAND3X1 U1132 ( .A(n1063), .B(n1062), .C(n1061), .Y(n1064) );
  AOI21X1 U1133 ( .A(n1064), .B(n1106), .C(n645), .Y(n1069) );
  NAND2X1 U1134 ( .A(n187), .B(n30), .Y(n1066) );
  NOR3X1 U1135 ( .A(n1067), .B(n1066), .C(n1135), .Y(n1068) );
  NAND3X1 U1136 ( .A(n65), .B(n1069), .C(n1068), .Y(nextState[0]) );
  NAND2X1 U1137 ( .A(n105), .B(n1071), .Y(n1080) );
  INVX2 U1138 ( .A(n124), .Y(n1072) );
  NAND2X1 U1139 ( .A(n1073), .B(n1072), .Y(n1079) );
  NAND2X1 U1140 ( .A(n1075), .B(n133), .Y(n1076) );
  AOI21X1 U1141 ( .A(n126), .B(n1077), .C(n1076), .Y(n1078) );
  NAND3X1 U1142 ( .A(n1080), .B(n1079), .C(n1078), .Y(nextState[4]) );
  AND2X2 U1143 ( .A(n1082), .B(n100), .Y(n1083) );
  MUX2X1 U1144 ( .B(n177), .A(n1083), .S(n107), .Y(n1095) );
  NAND2X1 U1145 ( .A(n155), .B(n1084), .Y(n1087) );
  NAND2X1 U1146 ( .A(n158), .B(n1085), .Y(n1086) );
  NAND2X1 U1147 ( .A(n1087), .B(n1086), .Y(n1088) );
  NAND2X1 U1148 ( .A(n1088), .B(n1106), .Y(n1094) );
  NAND2X1 U1149 ( .A(n1090), .B(n93), .Y(n1092) );
  NOR2X1 U1150 ( .A(n1092), .B(n1091), .Y(n1093) );
  NAND3X1 U1151 ( .A(n1095), .B(n1094), .C(n1093), .Y(nextState[2]) );
  INVX2 U1152 ( .A(N407), .Y(n1097) );
  NAND2X1 U1153 ( .A(prefillCounter[0]), .B(n149), .Y(n1096) );
  OAI21X1 U1154 ( .A(n1098), .B(n1097), .C(n1096), .Y(n915) );
  INVX2 U1155 ( .A(KEY_ERROR), .Y(n1106) );
  INVX2 U1156 ( .A(BYTE_READY), .Y(n1107) );
  INVX2 U1157 ( .A(n130), .Y(n1108) );
  INVX2 U1158 ( .A(OPCODE[1]), .Y(n1109) );
  INVX2 U1159 ( .A(OPCODE[0]), .Y(n1110) );
endmodule


module uart_edge_detector_1 ( CLK, RST, SERIAL_IN, START_BIT );
  input CLK, RST, SERIAL_IN;
  output START_BIT;
  wire   Q_int, Q_int2, n2, n4;

  DFFSR Q_int_reg ( .D(SERIAL_IN), .CLK(CLK), .R(n2), .S(1'b1), .Q(Q_int) );
  DFFSR Q_int2_reg ( .D(Q_int), .CLK(CLK), .R(n2), .S(1'b1), .Q(Q_int2) );
  NOR2X1 U7 ( .A(Q_int), .B(n4), .Y(START_BIT) );
  INVX2 U4 ( .A(RST), .Y(n2) );
  INVX2 U6 ( .A(Q_int2), .Y(n4) );
endmodule


module uart_error_1 ( RST, CLK, RBUF_FULL, CHK_ERROR, OE );
  input RST, CLK, RBUF_FULL, CHK_ERROR;
  output OE;
  wire   OE_prime, n1;

  DFFSR OE_reg ( .D(OE_prime), .CLK(CLK), .R(n1), .S(1'b1), .Q(OE) );
  AND2X2 U5 ( .A(RBUF_FULL), .B(CHK_ERROR), .Y(OE_prime) );
  INVX2 U3 ( .A(RST), .Y(n1) );
endmodule


module uart_rcu_1 ( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT, RBUF_LOAD, 
        TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR );
  input CLK, RST, START_BIT, STOP_RCVING, SB_DETECT;
  output RBUF_LOAD, TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR;
  wire   timerRunning, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N99, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, \add_46/carry[6] ,
         \add_46/carry[5] , \add_46/carry[4] , \add_46/carry[3] , n3, n4, n5,
         n6, n7, n25, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n81, n82;
  wire   [2:0] state;
  wire   [7:0] count;
  wire   [7:0] nextCount;
  wire   [2:0] nextState;

  DFFSR \count_reg[0]  ( .D(nextCount[0]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[0]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(n43), .CLK(CLK), .R(n4), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[0]) );
  DFFSR SBC_CLR_reg ( .D(n78), .CLK(CLK), .R(n4), .S(1'b1), .Q(SBC_CLR) );
  DFFSR TIMER_TRIG_reg ( .D(n79), .CLK(CLK), .R(n4), .S(1'b1), .Q(TIMER_TRIG)
         );
  DFFSR RBUF_LOAD_reg ( .D(n80), .CLK(CLK), .R(n4), .S(1'b1), .Q(RBUF_LOAD) );
  DFFSR timerRunning_reg ( .D(n74), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        timerRunning) );
  DFFSR \nextCount_reg[1]  ( .D(N32), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        nextCount[1]) );
  DFFSR \count_reg[1]  ( .D(nextCount[1]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        count[1]) );
  DFFSR \nextCount_reg[0]  ( .D(N31), .CLK(CLK), .R(1'b1), .S(n5), .Q(
        nextCount[0]) );
  DFFSR \nextCount_reg[2]  ( .D(N33), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        nextCount[2]) );
  DFFSR \count_reg[2]  ( .D(nextCount[2]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[2]) );
  DFFSR \nextCount_reg[3]  ( .D(N34), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[3]) );
  DFFSR \count_reg[3]  ( .D(nextCount[3]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[3]) );
  DFFSR \nextCount_reg[4]  ( .D(N35), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[4]) );
  DFFSR \count_reg[4]  ( .D(nextCount[4]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[4]) );
  DFFSR \nextCount_reg[5]  ( .D(N36), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[5]) );
  DFFSR \count_reg[5]  ( .D(nextCount[5]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[5]) );
  DFFSR \nextCount_reg[6]  ( .D(N37), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[6]) );
  DFFSR \count_reg[6]  ( .D(nextCount[6]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[6]) );
  DFFSR \nextCount_reg[7]  ( .D(N38), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[7]) );
  DFFSR \count_reg[7]  ( .D(nextCount[7]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[7]) );
  DFFSR SBC_EN_reg ( .D(n76), .CLK(CLK), .R(n4), .S(1'b1), .Q(SBC_EN) );
  AND2X2 U33 ( .A(N30), .B(timerRunning), .Y(N38) );
  AND2X2 U34 ( .A(N29), .B(timerRunning), .Y(N37) );
  AND2X2 U35 ( .A(N28), .B(timerRunning), .Y(N36) );
  AND2X2 U36 ( .A(N27), .B(timerRunning), .Y(N35) );
  AND2X2 U37 ( .A(N26), .B(timerRunning), .Y(N34) );
  AND2X2 U38 ( .A(N25), .B(timerRunning), .Y(N33) );
  AND2X2 U39 ( .A(N24), .B(timerRunning), .Y(N32) );
  OAI21X1 U54 ( .A(n49), .B(n45), .C(n50), .Y(n48) );
  OAI21X1 U55 ( .A(n46), .B(n44), .C(n45), .Y(n50) );
  NAND2X1 U56 ( .A(n51), .B(n52), .Y(n74) );
  OAI21X1 U57 ( .A(n53), .B(n54), .C(timerRunning), .Y(n52) );
  NAND2X1 U58 ( .A(n55), .B(n56), .Y(n54) );
  NAND2X1 U59 ( .A(n57), .B(n56), .Y(n75) );
  NAND3X1 U60 ( .A(n37), .B(n51), .C(CHK_ERROR), .Y(n57) );
  OAI21X1 U61 ( .A(n58), .B(n82), .C(n59), .Y(n76) );
  NAND2X1 U62 ( .A(n56), .B(n60), .Y(n58) );
  NAND2X1 U63 ( .A(n61), .B(n40), .Y(n56) );
  NAND3X1 U64 ( .A(n62), .B(n63), .C(n64), .Y(n77) );
  NAND3X1 U65 ( .A(n36), .B(n51), .C(SET_RBUF_FULL), .Y(n64) );
  NAND2X1 U66 ( .A(n60), .B(n63), .Y(n53) );
  NAND3X1 U67 ( .A(nextState[0]), .B(nextState[1]), .C(n61), .Y(n63) );
  NAND3X1 U68 ( .A(n38), .B(n40), .C(n61), .Y(n62) );
  OAI21X1 U69 ( .A(n65), .B(n47), .C(n51), .Y(n78) );
  OAI21X1 U70 ( .A(n65), .B(n81), .C(n51), .Y(n79) );
  NAND2X1 U71 ( .A(n60), .B(n59), .Y(n65) );
  NAND3X1 U72 ( .A(nextState[1]), .B(n38), .C(n41), .Y(n59) );
  NAND2X1 U73 ( .A(n66), .B(n55), .Y(n80) );
  NAND3X1 U74 ( .A(nextState[1]), .B(n38), .C(n61), .Y(n55) );
  NAND3X1 U75 ( .A(n60), .B(n51), .C(RBUF_LOAD), .Y(n66) );
  NAND3X1 U76 ( .A(nextState[0]), .B(n40), .C(n41), .Y(n51) );
  NAND3X1 U77 ( .A(n38), .B(n40), .C(n41), .Y(n60) );
  OAI21X1 U78 ( .A(n42), .B(n45), .C(n67), .Y(n61) );
  NAND3X1 U79 ( .A(state[0]), .B(n45), .C(state[1]), .Y(n67) );
  NAND2X1 U80 ( .A(n68), .B(n69), .Y(n49) );
  OAI21X1 U81 ( .A(n70), .B(n69), .C(n68), .Y(nextState[1]) );
  NOR2X1 U82 ( .A(N99), .B(state[2]), .Y(n70) );
  OAI21X1 U83 ( .A(state[2]), .B(n71), .C(n68), .Y(nextState[0]) );
  NAND2X1 U84 ( .A(state[1]), .B(n46), .Y(n68) );
  AOI21X1 U85 ( .A(START_BIT), .B(n46), .C(n72), .Y(n71) );
  OAI21X1 U86 ( .A(N99), .B(n69), .C(n73), .Y(n72) );
  NAND2X1 U87 ( .A(SB_DETECT), .B(state[1]), .Y(n73) );
  NAND2X1 U88 ( .A(state[0]), .B(n44), .Y(n69) );
  NAND2X1 U89 ( .A(n39), .B(timerRunning), .Y(N31) );
  DFFSR SET_RBUF_FULL_reg ( .D(n77), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        SET_RBUF_FULL) );
  DFFSR CHK_ERROR_reg ( .D(n75), .CLK(CLK), .R(n4), .S(1'b1), .Q(CHK_ERROR) );
  INVX2 U7 ( .A(RST), .Y(n4) );
  INVX2 U8 ( .A(RST), .Y(n5) );
  XNOR2X1 U24 ( .A(count[7]), .B(n3), .Y(N30) );
  NAND2X1 U31 ( .A(count[6]), .B(\add_46/carry[6] ), .Y(n3) );
  XOR2X1 U40 ( .A(\add_46/carry[6] ), .B(count[6]), .Y(N29) );
  AND2X1 U41 ( .A(count[5]), .B(\add_46/carry[5] ), .Y(\add_46/carry[6] ) );
  XOR2X1 U42 ( .A(\add_46/carry[5] ), .B(count[5]), .Y(N28) );
  AND2X1 U43 ( .A(count[4]), .B(\add_46/carry[4] ), .Y(\add_46/carry[5] ) );
  XOR2X1 U44 ( .A(\add_46/carry[4] ), .B(count[4]), .Y(N27) );
  AND2X1 U45 ( .A(count[3]), .B(\add_46/carry[3] ), .Y(\add_46/carry[4] ) );
  XOR2X1 U46 ( .A(\add_46/carry[3] ), .B(count[3]), .Y(N26) );
  AND2X1 U47 ( .A(count[2]), .B(count[1]), .Y(\add_46/carry[3] ) );
  XOR2X1 U48 ( .A(count[1]), .B(count[2]), .Y(N25) );
  INVX2 U49 ( .A(count[1]), .Y(N24) );
  OAI21X1 U50 ( .A(count[0]), .B(count[1]), .C(count[2]), .Y(n6) );
  NOR2X1 U51 ( .A(n35), .B(n6), .Y(n7) );
  OAI21X1 U52 ( .A(n7), .B(count[4]), .C(count[6]), .Y(n25) );
  OAI21X1 U53 ( .A(n34), .B(n25), .C(n32), .Y(N99) );
  INVX2 U90 ( .A(count[7]), .Y(n32) );
  INVX2 U91 ( .A(count[5]), .Y(n34) );
  INVX2 U92 ( .A(count[3]), .Y(n35) );
  INVX2 U93 ( .A(n53), .Y(n36) );
  INVX2 U94 ( .A(n58), .Y(n37) );
  INVX2 U95 ( .A(nextState[0]), .Y(n38) );
  INVX2 U96 ( .A(count[0]), .Y(n39) );
  INVX2 U97 ( .A(nextState[1]), .Y(n40) );
  INVX2 U98 ( .A(n61), .Y(n41) );
  INVX2 U99 ( .A(n49), .Y(n42) );
  INVX2 U100 ( .A(n48), .Y(n43) );
  INVX2 U101 ( .A(state[1]), .Y(n44) );
  INVX2 U102 ( .A(state[2]), .Y(n45) );
  INVX2 U103 ( .A(state[0]), .Y(n46) );
  INVX2 U104 ( .A(SBC_CLR), .Y(n47) );
  INVX2 U105 ( .A(TIMER_TRIG), .Y(n81) );
  INVX2 U106 ( .A(SBC_EN), .Y(n82) );
endmodule


module uart_rcv_buf_1 ( CLK, RST, LOAD_RBUF, LOAD_DATA, RCV_DATA );
  input [7:0] LOAD_DATA;
  output [7:0] RCV_DATA;
  input CLK, RST, LOAD_RBUF;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n2, n11, n13, n15, n17, n19, n21, n23,
         n24, n26;

  DFFSR \Q_int_reg[7]  ( .D(n11), .CLK(CLK), .R(n2), .S(1'b1), .Q(RCV_DATA[7])
         );
  DFFSR \Q_int_reg[6]  ( .D(n13), .CLK(CLK), .R(n2), .S(1'b1), .Q(RCV_DATA[6])
         );
  DFFSR \Q_int_reg[5]  ( .D(n15), .CLK(CLK), .R(n2), .S(1'b1), .Q(RCV_DATA[5])
         );
  DFFSR \Q_int_reg[4]  ( .D(n17), .CLK(CLK), .R(n2), .S(1'b1), .Q(RCV_DATA[4])
         );
  DFFSR \Q_int_reg[3]  ( .D(n19), .CLK(CLK), .R(n2), .S(1'b1), .Q(RCV_DATA[3])
         );
  DFFSR \Q_int_reg[2]  ( .D(n21), .CLK(CLK), .R(n2), .S(1'b1), .Q(RCV_DATA[2])
         );
  DFFSR \Q_int_reg[1]  ( .D(n23), .CLK(CLK), .R(n2), .S(1'b1), .Q(RCV_DATA[1])
         );
  DFFSR \Q_int_reg[0]  ( .D(n24), .CLK(CLK), .R(n2), .S(1'b1), .Q(RCV_DATA[0])
         );
  AOI22X1 U3 ( .A(LOAD_RBUF), .B(LOAD_DATA[0]), .C(RCV_DATA[0]), .D(n26), .Y(
        n1) );
  AOI22X1 U5 ( .A(LOAD_DATA[1]), .B(LOAD_RBUF), .C(RCV_DATA[1]), .D(n26), .Y(
        n3) );
  AOI22X1 U7 ( .A(LOAD_DATA[2]), .B(LOAD_RBUF), .C(RCV_DATA[2]), .D(n26), .Y(
        n4) );
  AOI22X1 U9 ( .A(LOAD_DATA[3]), .B(LOAD_RBUF), .C(RCV_DATA[3]), .D(n26), .Y(
        n5) );
  AOI22X1 U11 ( .A(LOAD_DATA[4]), .B(LOAD_RBUF), .C(RCV_DATA[4]), .D(n26), .Y(
        n6) );
  AOI22X1 U13 ( .A(LOAD_DATA[5]), .B(LOAD_RBUF), .C(RCV_DATA[5]), .D(n26), .Y(
        n7) );
  AOI22X1 U15 ( .A(LOAD_DATA[6]), .B(LOAD_RBUF), .C(RCV_DATA[6]), .D(n26), .Y(
        n8) );
  AOI22X1 U18 ( .A(LOAD_DATA[7]), .B(LOAD_RBUF), .C(RCV_DATA[7]), .D(n26), .Y(
        n9) );
  INVX2 U2 ( .A(RST), .Y(n2) );
  INVX2 U4 ( .A(n9), .Y(n11) );
  INVX2 U6 ( .A(n8), .Y(n13) );
  INVX2 U8 ( .A(n7), .Y(n15) );
  INVX2 U10 ( .A(n6), .Y(n17) );
  INVX2 U12 ( .A(n5), .Y(n19) );
  INVX2 U14 ( .A(n4), .Y(n21) );
  INVX2 U16 ( .A(n3), .Y(n23) );
  INVX2 U17 ( .A(n1), .Y(n24) );
  INVX2 U19 ( .A(LOAD_RBUF), .Y(n26) );
endmodule


module uart_rcv_buf_full_1 ( CLK, RST, CLR_RBUF, SET_RBUF_FULL, RBUF_FULL );
  input CLK, RST, CLR_RBUF, SET_RBUF_FULL;
  output RBUF_FULL;
  wire   n1, n3;

  DFFSR Q_int_reg ( .D(n3), .CLK(CLK), .R(n1), .S(1'b1), .Q(RBUF_FULL) );
  NOR2X1 U3 ( .A(RST), .B(CLR_RBUF), .Y(n1) );
  OR2X2 U4 ( .A(RBUF_FULL), .B(SET_RBUF_FULL), .Y(n3) );
endmodule


module uart_sb_check_1 ( RST, CLK, SBC_CLR, SBC_EN, STOP_DATA, SB_DETECT, SBE
 );
  input [1:0] STOP_DATA;
  input RST, CLK, SBC_CLR, SBC_EN;
  output SB_DETECT, SBE;
  wire   SBE_prime, sb_detect_flag, n7, n8, n9, n2, n4, n5, n6;

  DFFSR SB_DETECT_reg ( .D(sb_detect_flag), .CLK(CLK), .R(n2), .S(1'b1), .Q(
        SB_DETECT) );
  DFFSR SBE_reg ( .D(SBE_prime), .CLK(CLK), .R(n2), .S(1'b1), .Q(SBE) );
  OR2X2 U6 ( .A(SBC_CLR), .B(STOP_DATA[0]), .Y(n7) );
  NOR2X1 U10 ( .A(n7), .B(n8), .Y(sb_detect_flag) );
  NAND2X1 U11 ( .A(STOP_DATA[1]), .B(SBC_EN), .Y(n8) );
  NOR2X1 U12 ( .A(n6), .B(n9), .Y(SBE_prime) );
  OAI21X1 U13 ( .A(STOP_DATA[0]), .B(n4), .C(n5), .Y(n9) );
  INVX2 U4 ( .A(RST), .Y(n2) );
  INVX2 U7 ( .A(STOP_DATA[1]), .Y(n4) );
  INVX2 U8 ( .A(SBC_CLR), .Y(n5) );
  INVX2 U9 ( .A(SBC_EN), .Y(n6) );
endmodule


module uart_sr_10bit_1 ( CLK, RST, SHIFT_STROBE, SERIAL_IN, LOAD_DATA, 
        STOP_DATA );
  output [7:0] LOAD_DATA;
  output [1:0] STOP_DATA;
  input CLK, RST, SHIFT_STROBE, SERIAL_IN;
  wire   n3, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n33, n11, n13,
         n15, n17, n19, n21, n23, n25, n27, n29, n31, n34, n35;

  DFFSR \present_val_reg[9]  ( .D(n33), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        STOP_DATA[1]) );
  OAI21X1 U2 ( .A(n35), .B(n17), .C(n3), .Y(n14) );
  NAND2X1 U3 ( .A(LOAD_DATA[0]), .B(n17), .Y(n3) );
  OAI22X1 U4 ( .A(n17), .B(n34), .C(n13), .D(n35), .Y(n16) );
  OAI22X1 U6 ( .A(n17), .B(n31), .C(n13), .D(n34), .Y(n18) );
  OAI22X1 U8 ( .A(n17), .B(n29), .C(n13), .D(n31), .Y(n20) );
  OAI22X1 U10 ( .A(n17), .B(n27), .C(n13), .D(n29), .Y(n22) );
  OAI22X1 U12 ( .A(n17), .B(n25), .C(n13), .D(n27), .Y(n24) );
  OAI22X1 U14 ( .A(n17), .B(n23), .C(n13), .D(n25), .Y(n26) );
  OAI22X1 U16 ( .A(n17), .B(n21), .C(n13), .D(n23), .Y(n28) );
  OAI22X1 U18 ( .A(n17), .B(n19), .C(n13), .D(n21), .Y(n30) );
  OAI21X1 U22 ( .A(n13), .B(n19), .C(n12), .Y(n33) );
  NAND2X1 U23 ( .A(SERIAL_IN), .B(n13), .Y(n12) );
  DFFSR \present_val_reg[8]  ( .D(n30), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        STOP_DATA[0]) );
  DFFSR \present_val_reg[7]  ( .D(n28), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[7]) );
  DFFSR \present_val_reg[6]  ( .D(n26), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[6]) );
  DFFSR \present_val_reg[5]  ( .D(n24), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[5]) );
  DFFSR \present_val_reg[4]  ( .D(n22), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[4]) );
  DFFSR \present_val_reg[3]  ( .D(n20), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[3]) );
  DFFSR \present_val_reg[2]  ( .D(n18), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[2]) );
  DFFSR \present_val_reg[1]  ( .D(n16), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[1]) );
  DFFSR \present_val_reg[0]  ( .D(n14), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[0]) );
  INVX2 U21 ( .A(RST), .Y(n15) );
  INVX2 U24 ( .A(n13), .Y(n17) );
  INVX4 U25 ( .A(n11), .Y(n13) );
  INVX2 U26 ( .A(SHIFT_STROBE), .Y(n11) );
  INVX2 U27 ( .A(STOP_DATA[1]), .Y(n19) );
  INVX2 U28 ( .A(STOP_DATA[0]), .Y(n21) );
  INVX2 U29 ( .A(LOAD_DATA[7]), .Y(n23) );
  INVX2 U30 ( .A(LOAD_DATA[6]), .Y(n25) );
  INVX2 U31 ( .A(LOAD_DATA[5]), .Y(n27) );
  INVX2 U32 ( .A(LOAD_DATA[4]), .Y(n29) );
  INVX2 U33 ( .A(LOAD_DATA[3]), .Y(n31) );
  INVX2 U35 ( .A(LOAD_DATA[2]), .Y(n34) );
  INVX2 U36 ( .A(LOAD_DATA[1]), .Y(n35) );
endmodule


module keyreg_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  AND2X2 U2 ( .A(n21), .B(n17), .Y(n1) );
  XNOR2X1 U3 ( .A(n32), .B(n33), .Y(SUM[3]) );
  XOR2X1 U4 ( .A(n27), .B(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n31), .B(n30), .Y(n2) );
  NAND2X1 U6 ( .A(n35), .B(n36), .Y(n22) );
  INVX2 U7 ( .A(n41), .Y(SUM[0]) );
  XNOR2X1 U8 ( .A(n3), .B(n4), .Y(SUM[7]) );
  XOR2X1 U9 ( .A(B[7]), .B(A[7]), .Y(n4) );
  AOI21X1 U10 ( .A(n5), .B(n6), .C(n7), .Y(n3) );
  NAND2X1 U11 ( .A(n8), .B(n9), .Y(n7) );
  NAND2X1 U12 ( .A(n10), .B(n11), .Y(n8) );
  AND2X2 U13 ( .A(n12), .B(n11), .Y(n5) );
  XNOR2X1 U14 ( .A(n13), .B(n14), .Y(SUM[6]) );
  AND2X2 U15 ( .A(n11), .B(n9), .Y(n14) );
  NAND2X1 U16 ( .A(B[6]), .B(A[6]), .Y(n9) );
  OR2X2 U17 ( .A(A[6]), .B(B[6]), .Y(n11) );
  AOI21X1 U18 ( .A(n6), .B(n12), .C(n10), .Y(n13) );
  INVX2 U19 ( .A(n15), .Y(n10) );
  XNOR2X1 U20 ( .A(n6), .B(n16), .Y(SUM[5]) );
  NAND2X1 U21 ( .A(n12), .B(n15), .Y(n16) );
  NAND2X1 U22 ( .A(B[5]), .B(A[5]), .Y(n15) );
  OR2X2 U23 ( .A(A[5]), .B(B[5]), .Y(n12) );
  NAND3X1 U24 ( .A(n17), .B(n18), .C(n19), .Y(n6) );
  NAND3X1 U25 ( .A(n20), .B(n21), .C(n22), .Y(n19) );
  INVX2 U26 ( .A(n23), .Y(n20) );
  NAND3X1 U27 ( .A(n24), .B(n21), .C(n25), .Y(n18) );
  XOR2X1 U28 ( .A(n26), .B(n1), .Y(SUM[4]) );
  NAND2X1 U29 ( .A(B[4]), .B(A[4]), .Y(n17) );
  OR2X2 U30 ( .A(A[4]), .B(B[4]), .Y(n21) );
  OAI21X1 U31 ( .A(n27), .B(n23), .C(n28), .Y(n26) );
  NAND2X1 U32 ( .A(n24), .B(n25), .Y(n28) );
  NAND2X1 U33 ( .A(n29), .B(n30), .Y(n25) );
  NAND2X1 U34 ( .A(n31), .B(n24), .Y(n23) );
  NAND2X1 U35 ( .A(n24), .B(n29), .Y(n33) );
  NAND2X1 U36 ( .A(B[3]), .B(A[3]), .Y(n29) );
  OR2X2 U37 ( .A(A[3]), .B(B[3]), .Y(n24) );
  NAND2X1 U38 ( .A(n30), .B(n34), .Y(n32) );
  NAND2X1 U39 ( .A(n22), .B(n31), .Y(n34) );
  NAND2X1 U40 ( .A(B[2]), .B(A[2]), .Y(n30) );
  OR2X2 U41 ( .A(A[2]), .B(B[2]), .Y(n31) );
  INVX2 U42 ( .A(n22), .Y(n27) );
  NAND2X1 U43 ( .A(n38), .B(n37), .Y(n35) );
  AND2X2 U44 ( .A(A[0]), .B(B[0]), .Y(n38) );
  XOR2X1 U45 ( .A(n39), .B(n40), .Y(SUM[1]) );
  NAND2X1 U46 ( .A(n37), .B(n36), .Y(n39) );
  NAND2X1 U47 ( .A(B[1]), .B(A[1]), .Y(n36) );
  OR2X2 U48 ( .A(A[1]), .B(B[1]), .Y(n37) );
  OAI21X1 U49 ( .A(A[0]), .B(B[0]), .C(n40), .Y(n41) );
  NAND2X1 U50 ( .A(B[0]), .B(A[0]), .Y(n40) );
endmodule


module keyreg_1 ( CLK, RST, SBE, OE, RBUF_FULL, RCV_DATA, PLAINKEY, KEY_ERROR, 
        PROG_ERROR, CLR_RBUFF, PARITY_ERROR );
  input [7:0] RCV_DATA;
  output [63:0] PLAINKEY;
  input CLK, RST, SBE, OE, RBUF_FULL;
  output KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR;
  wire   parityError, nextParityError, N1792, N1793, N1794, N1795, N1796,
         N1797, N1798, N1799, n12, n13, n15, n18, n22, n24, n26, n28, n30, n32,
         n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60,
         n62, n64, n66, n68, n70, n72, n74, n76, n78, n80, n82, n84, n86, n88,
         n90, n92, n94, n96, n98, n100, n102, n104, n106, n108, n110, n112,
         n114, n116, n118, n120, n122, n124, n126, n128, n130, n132, n134,
         n136, n138, n140, n142, n144, n146, n148, n1178, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1, n2,
         n4, n5, n6, n7, n8, n9, n10, n11, n14, n16, n17, n19, n20, n21, n23,
         n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51,
         n53, n55, n57, n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79,
         n81, n83, n85, n87, n89, n91, n93, n95, n97, n99, n101, n103, n105,
         n107, n109, n111, n113, n115, n117, n119, n121, n123, n125, n127,
         n129, n131, n133, n135, n137, n139, n141, n143, n145, n147, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1267,
         n1268, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695;
  wire   [3:0] state;
  wire   [3:0] keyCount;
  wire   [7:0] address;
  wire   [63:0] currentPlainKey;
  wire   [7:0] parityAccumulator;

  DFFPOSX1 \keyCount_reg[0]  ( .D(n1356), .CLK(CLK), .Q(keyCount[0]) );
  DFFPOSX1 \keyCount_reg[2]  ( .D(n1349), .CLK(CLK), .Q(keyCount[2]) );
  DFFPOSX1 \keyCount_reg[3]  ( .D(n1355), .CLK(CLK), .Q(keyCount[3]) );
  DFFSR \state_reg[0]  ( .D(n1353), .CLK(CLK), .R(n252), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[1]  ( .D(n1351), .CLK(CLK), .R(n252), .S(1'b1), .Q(state[1]) );
  DFFSR \state_reg[2]  ( .D(n1352), .CLK(CLK), .R(n253), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[3]  ( .D(n1354), .CLK(CLK), .R(n252), .S(1'b1), .Q(state[3]) );
  DFFPOSX1 \parityAccumulator_reg[0]  ( .D(n1348), .CLK(CLK), .Q(
        parityAccumulator[0]) );
  DFFPOSX1 \parityAccumulator_reg[1]  ( .D(n1347), .CLK(CLK), .Q(
        parityAccumulator[1]) );
  DFFPOSX1 \parityAccumulator_reg[2]  ( .D(n1346), .CLK(CLK), .Q(
        parityAccumulator[2]) );
  DFFPOSX1 \parityAccumulator_reg[3]  ( .D(n1345), .CLK(CLK), .Q(
        parityAccumulator[3]) );
  DFFPOSX1 \parityAccumulator_reg[4]  ( .D(n1344), .CLK(CLK), .Q(
        parityAccumulator[4]) );
  DFFPOSX1 \parityAccumulator_reg[5]  ( .D(n1343), .CLK(CLK), .Q(
        parityAccumulator[5]) );
  DFFPOSX1 \parityAccumulator_reg[6]  ( .D(n1342), .CLK(CLK), .Q(
        parityAccumulator[6]) );
  DFFPOSX1 \parityAccumulator_reg[7]  ( .D(n1341), .CLK(CLK), .Q(
        parityAccumulator[7]) );
  DFFPOSX1 \keyCount_reg[1]  ( .D(n1350), .CLK(CLK), .Q(keyCount[1]) );
  DFFSR PARITY_ERROR_reg ( .D(nextParityError), .CLK(CLK), .R(n253), .S(1'b1), 
        .Q(PARITY_ERROR) );
  DFFSR parityError_reg ( .D(nextParityError), .CLK(CLK), .R(n253), .S(1'b1), 
        .Q(parityError) );
  DFFPOSX1 \address_reg[7]  ( .D(n1340), .CLK(CLK), .Q(address[7]) );
  DFFPOSX1 \address_reg[6]  ( .D(n1339), .CLK(CLK), .Q(address[6]) );
  DFFPOSX1 \address_reg[5]  ( .D(n1338), .CLK(CLK), .Q(address[5]) );
  DFFPOSX1 \address_reg[4]  ( .D(n1337), .CLK(CLK), .Q(address[4]) );
  DFFPOSX1 \address_reg[3]  ( .D(n1336), .CLK(CLK), .Q(address[3]) );
  DFFPOSX1 \address_reg[2]  ( .D(n1335), .CLK(CLK), .Q(address[2]) );
  DFFPOSX1 \address_reg[1]  ( .D(n1334), .CLK(CLK), .Q(address[1]) );
  DFFPOSX1 \address_reg[0]  ( .D(n1333), .CLK(CLK), .Q(address[0]) );
  DFFPOSX1 \currentPlainKey_reg[63]  ( .D(n1269), .CLK(CLK), .Q(
        currentPlainKey[63]) );
  DFFPOSX1 \currentPlainKey_reg[62]  ( .D(n1270), .CLK(CLK), .Q(
        currentPlainKey[62]) );
  DFFPOSX1 \currentPlainKey_reg[61]  ( .D(n1271), .CLK(CLK), .Q(
        currentPlainKey[61]) );
  DFFPOSX1 \currentPlainKey_reg[60]  ( .D(n1272), .CLK(CLK), .Q(
        currentPlainKey[60]) );
  DFFPOSX1 \currentPlainKey_reg[59]  ( .D(n1273), .CLK(CLK), .Q(
        currentPlainKey[59]) );
  DFFPOSX1 \currentPlainKey_reg[58]  ( .D(n1274), .CLK(CLK), .Q(
        currentPlainKey[58]) );
  DFFPOSX1 \currentPlainKey_reg[57]  ( .D(n1275), .CLK(CLK), .Q(
        currentPlainKey[57]) );
  DFFPOSX1 \currentPlainKey_reg[56]  ( .D(n1276), .CLK(CLK), .Q(
        currentPlainKey[56]) );
  DFFPOSX1 \currentPlainKey_reg[55]  ( .D(n1277), .CLK(CLK), .Q(
        currentPlainKey[55]) );
  DFFPOSX1 \currentPlainKey_reg[54]  ( .D(n1278), .CLK(CLK), .Q(
        currentPlainKey[54]) );
  DFFPOSX1 \currentPlainKey_reg[53]  ( .D(n1279), .CLK(CLK), .Q(
        currentPlainKey[53]) );
  DFFPOSX1 \currentPlainKey_reg[52]  ( .D(n1280), .CLK(CLK), .Q(
        currentPlainKey[52]) );
  DFFPOSX1 \currentPlainKey_reg[51]  ( .D(n1281), .CLK(CLK), .Q(
        currentPlainKey[51]) );
  DFFPOSX1 \currentPlainKey_reg[50]  ( .D(n1282), .CLK(CLK), .Q(
        currentPlainKey[50]) );
  DFFPOSX1 \currentPlainKey_reg[49]  ( .D(n1283), .CLK(CLK), .Q(
        currentPlainKey[49]) );
  DFFPOSX1 \currentPlainKey_reg[48]  ( .D(n1284), .CLK(CLK), .Q(
        currentPlainKey[48]) );
  DFFPOSX1 \currentPlainKey_reg[47]  ( .D(n1285), .CLK(CLK), .Q(
        currentPlainKey[47]) );
  DFFPOSX1 \currentPlainKey_reg[46]  ( .D(n1286), .CLK(CLK), .Q(
        currentPlainKey[46]) );
  DFFPOSX1 \currentPlainKey_reg[45]  ( .D(n1287), .CLK(CLK), .Q(
        currentPlainKey[45]) );
  DFFPOSX1 \currentPlainKey_reg[44]  ( .D(n1288), .CLK(CLK), .Q(
        currentPlainKey[44]) );
  DFFPOSX1 \currentPlainKey_reg[43]  ( .D(n1289), .CLK(CLK), .Q(
        currentPlainKey[43]) );
  DFFPOSX1 \currentPlainKey_reg[42]  ( .D(n1290), .CLK(CLK), .Q(
        currentPlainKey[42]) );
  DFFPOSX1 \currentPlainKey_reg[41]  ( .D(n1291), .CLK(CLK), .Q(
        currentPlainKey[41]) );
  DFFPOSX1 \currentPlainKey_reg[40]  ( .D(n1292), .CLK(CLK), .Q(
        currentPlainKey[40]) );
  DFFPOSX1 \currentPlainKey_reg[39]  ( .D(n1293), .CLK(CLK), .Q(
        currentPlainKey[39]) );
  DFFPOSX1 \currentPlainKey_reg[38]  ( .D(n1294), .CLK(CLK), .Q(
        currentPlainKey[38]) );
  DFFPOSX1 \currentPlainKey_reg[37]  ( .D(n1295), .CLK(CLK), .Q(
        currentPlainKey[37]) );
  DFFPOSX1 \currentPlainKey_reg[36]  ( .D(n1296), .CLK(CLK), .Q(
        currentPlainKey[36]) );
  DFFPOSX1 \currentPlainKey_reg[35]  ( .D(n1297), .CLK(CLK), .Q(
        currentPlainKey[35]) );
  DFFPOSX1 \currentPlainKey_reg[34]  ( .D(n1298), .CLK(CLK), .Q(
        currentPlainKey[34]) );
  DFFPOSX1 \currentPlainKey_reg[33]  ( .D(n1299), .CLK(CLK), .Q(
        currentPlainKey[33]) );
  DFFPOSX1 \currentPlainKey_reg[32]  ( .D(n1300), .CLK(CLK), .Q(
        currentPlainKey[32]) );
  DFFPOSX1 \currentPlainKey_reg[31]  ( .D(n1301), .CLK(CLK), .Q(
        currentPlainKey[31]) );
  DFFPOSX1 \currentPlainKey_reg[30]  ( .D(n1302), .CLK(CLK), .Q(
        currentPlainKey[30]) );
  DFFPOSX1 \currentPlainKey_reg[29]  ( .D(n1303), .CLK(CLK), .Q(
        currentPlainKey[29]) );
  DFFPOSX1 \currentPlainKey_reg[28]  ( .D(n1304), .CLK(CLK), .Q(
        currentPlainKey[28]) );
  DFFPOSX1 \currentPlainKey_reg[27]  ( .D(n1305), .CLK(CLK), .Q(
        currentPlainKey[27]) );
  DFFPOSX1 \currentPlainKey_reg[26]  ( .D(n1306), .CLK(CLK), .Q(
        currentPlainKey[26]) );
  DFFPOSX1 \currentPlainKey_reg[25]  ( .D(n1307), .CLK(CLK), .Q(
        currentPlainKey[25]) );
  DFFPOSX1 \currentPlainKey_reg[24]  ( .D(n1308), .CLK(CLK), .Q(
        currentPlainKey[24]) );
  DFFPOSX1 \currentPlainKey_reg[23]  ( .D(n1309), .CLK(CLK), .Q(
        currentPlainKey[23]) );
  DFFPOSX1 \currentPlainKey_reg[22]  ( .D(n1310), .CLK(CLK), .Q(
        currentPlainKey[22]) );
  DFFPOSX1 \currentPlainKey_reg[21]  ( .D(n1311), .CLK(CLK), .Q(
        currentPlainKey[21]) );
  DFFPOSX1 \currentPlainKey_reg[20]  ( .D(n1312), .CLK(CLK), .Q(
        currentPlainKey[20]) );
  DFFPOSX1 \currentPlainKey_reg[19]  ( .D(n1313), .CLK(CLK), .Q(
        currentPlainKey[19]) );
  DFFPOSX1 \currentPlainKey_reg[18]  ( .D(n1314), .CLK(CLK), .Q(
        currentPlainKey[18]) );
  DFFPOSX1 \currentPlainKey_reg[17]  ( .D(n1315), .CLK(CLK), .Q(
        currentPlainKey[17]) );
  DFFPOSX1 \currentPlainKey_reg[16]  ( .D(n1316), .CLK(CLK), .Q(
        currentPlainKey[16]) );
  DFFPOSX1 \currentPlainKey_reg[15]  ( .D(n1317), .CLK(CLK), .Q(
        currentPlainKey[15]) );
  DFFPOSX1 \currentPlainKey_reg[14]  ( .D(n1318), .CLK(CLK), .Q(
        currentPlainKey[14]) );
  DFFPOSX1 \currentPlainKey_reg[13]  ( .D(n1319), .CLK(CLK), .Q(
        currentPlainKey[13]) );
  DFFPOSX1 \currentPlainKey_reg[12]  ( .D(n1320), .CLK(CLK), .Q(
        currentPlainKey[12]) );
  DFFPOSX1 \currentPlainKey_reg[11]  ( .D(n1321), .CLK(CLK), .Q(
        currentPlainKey[11]) );
  DFFPOSX1 \currentPlainKey_reg[10]  ( .D(n1322), .CLK(CLK), .Q(
        currentPlainKey[10]) );
  DFFPOSX1 \currentPlainKey_reg[9]  ( .D(n1323), .CLK(CLK), .Q(
        currentPlainKey[9]) );
  DFFPOSX1 \currentPlainKey_reg[8]  ( .D(n1324), .CLK(CLK), .Q(
        currentPlainKey[8]) );
  DFFPOSX1 \currentPlainKey_reg[7]  ( .D(n1325), .CLK(CLK), .Q(
        currentPlainKey[7]) );
  DFFPOSX1 \currentPlainKey_reg[6]  ( .D(n1326), .CLK(CLK), .Q(
        currentPlainKey[6]) );
  DFFPOSX1 \currentPlainKey_reg[5]  ( .D(n1327), .CLK(CLK), .Q(
        currentPlainKey[5]) );
  DFFPOSX1 \currentPlainKey_reg[4]  ( .D(n1328), .CLK(CLK), .Q(
        currentPlainKey[4]) );
  DFFPOSX1 \currentPlainKey_reg[3]  ( .D(n1329), .CLK(CLK), .Q(
        currentPlainKey[3]) );
  DFFPOSX1 \currentPlainKey_reg[2]  ( .D(n1330), .CLK(CLK), .Q(
        currentPlainKey[2]) );
  DFFPOSX1 \currentPlainKey_reg[1]  ( .D(n1331), .CLK(CLK), .Q(
        currentPlainKey[1]) );
  DFFPOSX1 \currentPlainKey_reg[0]  ( .D(n1332), .CLK(CLK), .Q(
        currentPlainKey[0]) );
  DFFPOSX1 \PLAINKEY_reg[63]  ( .D(n1260), .CLK(CLK), .Q(PLAINKEY[63]) );
  DFFPOSX1 \PLAINKEY_reg[62]  ( .D(n1259), .CLK(CLK), .Q(PLAINKEY[62]) );
  DFFPOSX1 \PLAINKEY_reg[61]  ( .D(n1258), .CLK(CLK), .Q(PLAINKEY[61]) );
  DFFPOSX1 \PLAINKEY_reg[60]  ( .D(n1257), .CLK(CLK), .Q(PLAINKEY[60]) );
  DFFPOSX1 \PLAINKEY_reg[59]  ( .D(n1256), .CLK(CLK), .Q(PLAINKEY[59]) );
  DFFPOSX1 \PLAINKEY_reg[58]  ( .D(n1255), .CLK(CLK), .Q(PLAINKEY[58]) );
  DFFPOSX1 \PLAINKEY_reg[57]  ( .D(n1254), .CLK(CLK), .Q(PLAINKEY[57]) );
  DFFPOSX1 \PLAINKEY_reg[56]  ( .D(n1253), .CLK(CLK), .Q(PLAINKEY[56]) );
  DFFPOSX1 \PLAINKEY_reg[55]  ( .D(n1252), .CLK(CLK), .Q(PLAINKEY[55]) );
  DFFPOSX1 \PLAINKEY_reg[54]  ( .D(n1251), .CLK(CLK), .Q(PLAINKEY[54]) );
  DFFPOSX1 \PLAINKEY_reg[53]  ( .D(n1250), .CLK(CLK), .Q(PLAINKEY[53]) );
  DFFPOSX1 \PLAINKEY_reg[52]  ( .D(n1249), .CLK(CLK), .Q(PLAINKEY[52]) );
  DFFPOSX1 \PLAINKEY_reg[51]  ( .D(n1248), .CLK(CLK), .Q(PLAINKEY[51]) );
  DFFPOSX1 \PLAINKEY_reg[50]  ( .D(n1247), .CLK(CLK), .Q(PLAINKEY[50]) );
  DFFPOSX1 \PLAINKEY_reg[49]  ( .D(n1246), .CLK(CLK), .Q(PLAINKEY[49]) );
  DFFPOSX1 \PLAINKEY_reg[48]  ( .D(n1245), .CLK(CLK), .Q(PLAINKEY[48]) );
  DFFPOSX1 \PLAINKEY_reg[47]  ( .D(n1244), .CLK(CLK), .Q(PLAINKEY[47]) );
  DFFPOSX1 \PLAINKEY_reg[46]  ( .D(n1243), .CLK(CLK), .Q(PLAINKEY[46]) );
  DFFPOSX1 \PLAINKEY_reg[45]  ( .D(n1242), .CLK(CLK), .Q(PLAINKEY[45]) );
  DFFPOSX1 \PLAINKEY_reg[44]  ( .D(n1241), .CLK(CLK), .Q(PLAINKEY[44]) );
  DFFPOSX1 \PLAINKEY_reg[43]  ( .D(n1240), .CLK(CLK), .Q(PLAINKEY[43]) );
  DFFPOSX1 \PLAINKEY_reg[42]  ( .D(n1239), .CLK(CLK), .Q(PLAINKEY[42]) );
  DFFPOSX1 \PLAINKEY_reg[41]  ( .D(n1238), .CLK(CLK), .Q(PLAINKEY[41]) );
  DFFPOSX1 \PLAINKEY_reg[40]  ( .D(n1237), .CLK(CLK), .Q(PLAINKEY[40]) );
  DFFPOSX1 \PLAINKEY_reg[39]  ( .D(n1236), .CLK(CLK), .Q(PLAINKEY[39]) );
  DFFPOSX1 \PLAINKEY_reg[38]  ( .D(n1235), .CLK(CLK), .Q(PLAINKEY[38]) );
  DFFPOSX1 \PLAINKEY_reg[37]  ( .D(n1234), .CLK(CLK), .Q(PLAINKEY[37]) );
  DFFPOSX1 \PLAINKEY_reg[36]  ( .D(n1233), .CLK(CLK), .Q(PLAINKEY[36]) );
  DFFPOSX1 \PLAINKEY_reg[35]  ( .D(n1232), .CLK(CLK), .Q(PLAINKEY[35]) );
  DFFPOSX1 \PLAINKEY_reg[34]  ( .D(n1231), .CLK(CLK), .Q(PLAINKEY[34]) );
  DFFPOSX1 \PLAINKEY_reg[33]  ( .D(n1230), .CLK(CLK), .Q(PLAINKEY[33]) );
  DFFPOSX1 \PLAINKEY_reg[32]  ( .D(n1229), .CLK(CLK), .Q(PLAINKEY[32]) );
  DFFPOSX1 \PLAINKEY_reg[31]  ( .D(n1228), .CLK(CLK), .Q(PLAINKEY[31]) );
  DFFPOSX1 \PLAINKEY_reg[30]  ( .D(n1227), .CLK(CLK), .Q(PLAINKEY[30]) );
  DFFPOSX1 \PLAINKEY_reg[29]  ( .D(n1226), .CLK(CLK), .Q(PLAINKEY[29]) );
  DFFPOSX1 \PLAINKEY_reg[28]  ( .D(n1225), .CLK(CLK), .Q(PLAINKEY[28]) );
  DFFPOSX1 \PLAINKEY_reg[27]  ( .D(n1224), .CLK(CLK), .Q(PLAINKEY[27]) );
  DFFPOSX1 \PLAINKEY_reg[26]  ( .D(n1223), .CLK(CLK), .Q(PLAINKEY[26]) );
  DFFPOSX1 \PLAINKEY_reg[25]  ( .D(n1222), .CLK(CLK), .Q(PLAINKEY[25]) );
  DFFPOSX1 \PLAINKEY_reg[24]  ( .D(n1221), .CLK(CLK), .Q(PLAINKEY[24]) );
  DFFPOSX1 \PLAINKEY_reg[23]  ( .D(n1220), .CLK(CLK), .Q(PLAINKEY[23]) );
  DFFPOSX1 \PLAINKEY_reg[22]  ( .D(n1219), .CLK(CLK), .Q(PLAINKEY[22]) );
  DFFPOSX1 \PLAINKEY_reg[21]  ( .D(n1218), .CLK(CLK), .Q(PLAINKEY[21]) );
  DFFPOSX1 \PLAINKEY_reg[20]  ( .D(n1217), .CLK(CLK), .Q(PLAINKEY[20]) );
  DFFPOSX1 \PLAINKEY_reg[19]  ( .D(n1216), .CLK(CLK), .Q(PLAINKEY[19]) );
  DFFPOSX1 \PLAINKEY_reg[18]  ( .D(n1215), .CLK(CLK), .Q(PLAINKEY[18]) );
  DFFPOSX1 \PLAINKEY_reg[17]  ( .D(n1214), .CLK(CLK), .Q(PLAINKEY[17]) );
  DFFPOSX1 \PLAINKEY_reg[16]  ( .D(n1213), .CLK(CLK), .Q(PLAINKEY[16]) );
  DFFPOSX1 \PLAINKEY_reg[15]  ( .D(n1212), .CLK(CLK), .Q(PLAINKEY[15]) );
  DFFPOSX1 \PLAINKEY_reg[14]  ( .D(n1211), .CLK(CLK), .Q(PLAINKEY[14]) );
  DFFPOSX1 \PLAINKEY_reg[13]  ( .D(n1210), .CLK(CLK), .Q(PLAINKEY[13]) );
  DFFPOSX1 \PLAINKEY_reg[12]  ( .D(n1209), .CLK(CLK), .Q(PLAINKEY[12]) );
  DFFPOSX1 \PLAINKEY_reg[11]  ( .D(n1208), .CLK(CLK), .Q(PLAINKEY[11]) );
  DFFPOSX1 \PLAINKEY_reg[10]  ( .D(n1207), .CLK(CLK), .Q(PLAINKEY[10]) );
  DFFPOSX1 \PLAINKEY_reg[9]  ( .D(n1206), .CLK(CLK), .Q(PLAINKEY[9]) );
  DFFPOSX1 \PLAINKEY_reg[8]  ( .D(n1205), .CLK(CLK), .Q(PLAINKEY[8]) );
  DFFPOSX1 \PLAINKEY_reg[7]  ( .D(n1204), .CLK(CLK), .Q(PLAINKEY[7]) );
  DFFPOSX1 \PLAINKEY_reg[6]  ( .D(n1203), .CLK(CLK), .Q(PLAINKEY[6]) );
  DFFPOSX1 \PLAINKEY_reg[5]  ( .D(n1202), .CLK(CLK), .Q(PLAINKEY[5]) );
  DFFPOSX1 \PLAINKEY_reg[4]  ( .D(n1201), .CLK(CLK), .Q(PLAINKEY[4]) );
  DFFPOSX1 \PLAINKEY_reg[3]  ( .D(n1200), .CLK(CLK), .Q(PLAINKEY[3]) );
  DFFPOSX1 \PLAINKEY_reg[2]  ( .D(n1199), .CLK(CLK), .Q(PLAINKEY[2]) );
  DFFPOSX1 \PLAINKEY_reg[1]  ( .D(n1198), .CLK(CLK), .Q(PLAINKEY[1]) );
  DFFPOSX1 \PLAINKEY_reg[0]  ( .D(n1197), .CLK(CLK), .Q(PLAINKEY[0]) );
  NAND3X1 U9 ( .A(parityAccumulator[7]), .B(parityAccumulator[6]), .C(n15), 
        .Y(n13) );
  NOR2X1 U10 ( .A(n1627), .B(n1628), .Y(n15) );
  NAND3X1 U11 ( .A(parityAccumulator[3]), .B(parityAccumulator[2]), .C(n18), 
        .Y(n12) );
  NOR2X1 U12 ( .A(n1623), .B(n1624), .Y(n18) );
  OAI21X1 U13 ( .A(n239), .B(n1694), .C(n22), .Y(n1197) );
  NAND2X1 U14 ( .A(PLAINKEY[0]), .B(n244), .Y(n22) );
  OAI21X1 U15 ( .A(n239), .B(n1693), .C(n24), .Y(n1198) );
  NAND2X1 U16 ( .A(PLAINKEY[1]), .B(n247), .Y(n24) );
  OAI21X1 U17 ( .A(n239), .B(n1692), .C(n26), .Y(n1199) );
  NAND2X1 U18 ( .A(PLAINKEY[2]), .B(n247), .Y(n26) );
  OAI21X1 U19 ( .A(n239), .B(n1691), .C(n28), .Y(n1200) );
  NAND2X1 U20 ( .A(PLAINKEY[3]), .B(n247), .Y(n28) );
  OAI21X1 U21 ( .A(n239), .B(n1690), .C(n30), .Y(n1201) );
  NAND2X1 U22 ( .A(PLAINKEY[4]), .B(n247), .Y(n30) );
  OAI21X1 U24 ( .A(n239), .B(n1689), .C(n32), .Y(n1202) );
  NAND2X1 U25 ( .A(PLAINKEY[5]), .B(n247), .Y(n32) );
  OAI21X1 U27 ( .A(n239), .B(n1688), .C(n34), .Y(n1203) );
  NAND2X1 U28 ( .A(PLAINKEY[6]), .B(n247), .Y(n34) );
  OAI21X1 U30 ( .A(n239), .B(n1687), .C(n36), .Y(n1204) );
  NAND2X1 U31 ( .A(PLAINKEY[7]), .B(n247), .Y(n36) );
  OAI21X1 U33 ( .A(n239), .B(n1686), .C(n38), .Y(n1205) );
  NAND2X1 U34 ( .A(PLAINKEY[8]), .B(n247), .Y(n38) );
  OAI21X1 U36 ( .A(n240), .B(n1685), .C(n40), .Y(n1206) );
  NAND2X1 U37 ( .A(PLAINKEY[9]), .B(n247), .Y(n40) );
  OAI21X1 U39 ( .A(n240), .B(n1684), .C(n42), .Y(n1207) );
  NAND2X1 U40 ( .A(PLAINKEY[10]), .B(n247), .Y(n42) );
  OAI21X1 U42 ( .A(n240), .B(n1683), .C(n44), .Y(n1208) );
  NAND2X1 U43 ( .A(PLAINKEY[11]), .B(n246), .Y(n44) );
  OAI21X1 U45 ( .A(n240), .B(n1682), .C(n46), .Y(n1209) );
  NAND2X1 U46 ( .A(PLAINKEY[12]), .B(n246), .Y(n46) );
  OAI21X1 U48 ( .A(n240), .B(n1681), .C(n48), .Y(n1210) );
  NAND2X1 U49 ( .A(PLAINKEY[13]), .B(n246), .Y(n48) );
  OAI21X1 U51 ( .A(n240), .B(n1680), .C(n50), .Y(n1211) );
  NAND2X1 U52 ( .A(PLAINKEY[14]), .B(n246), .Y(n50) );
  OAI21X1 U54 ( .A(n240), .B(n1679), .C(n52), .Y(n1212) );
  NAND2X1 U55 ( .A(PLAINKEY[15]), .B(n246), .Y(n52) );
  OAI21X1 U57 ( .A(n241), .B(n1678), .C(n54), .Y(n1213) );
  NAND2X1 U58 ( .A(PLAINKEY[16]), .B(n246), .Y(n54) );
  OAI21X1 U60 ( .A(n241), .B(n1677), .C(n56), .Y(n1214) );
  NAND2X1 U61 ( .A(PLAINKEY[17]), .B(n246), .Y(n56) );
  OAI21X1 U63 ( .A(n241), .B(n1676), .C(n58), .Y(n1215) );
  NAND2X1 U64 ( .A(PLAINKEY[18]), .B(n246), .Y(n58) );
  OAI21X1 U66 ( .A(n241), .B(n1675), .C(n60), .Y(n1216) );
  NAND2X1 U67 ( .A(PLAINKEY[19]), .B(n246), .Y(n60) );
  OAI21X1 U69 ( .A(n241), .B(n1674), .C(n62), .Y(n1217) );
  NAND2X1 U70 ( .A(PLAINKEY[20]), .B(n246), .Y(n62) );
  OAI21X1 U72 ( .A(n241), .B(n1673), .C(n64), .Y(n1218) );
  NAND2X1 U73 ( .A(PLAINKEY[21]), .B(n246), .Y(n64) );
  OAI21X1 U75 ( .A(n241), .B(n1672), .C(n66), .Y(n1219) );
  NAND2X1 U76 ( .A(PLAINKEY[22]), .B(n246), .Y(n66) );
  OAI21X1 U78 ( .A(n242), .B(n1671), .C(n68), .Y(n1220) );
  NAND2X1 U79 ( .A(PLAINKEY[23]), .B(n246), .Y(n68) );
  OAI21X1 U81 ( .A(n241), .B(n1670), .C(n70), .Y(n1221) );
  NAND2X1 U82 ( .A(PLAINKEY[24]), .B(n246), .Y(n70) );
  OAI21X1 U84 ( .A(n240), .B(n1669), .C(n72), .Y(n1222) );
  NAND2X1 U85 ( .A(PLAINKEY[25]), .B(n246), .Y(n72) );
  OAI21X1 U87 ( .A(n242), .B(n1668), .C(n74), .Y(n1223) );
  NAND2X1 U88 ( .A(PLAINKEY[26]), .B(n246), .Y(n74) );
  OAI21X1 U90 ( .A(n242), .B(n1667), .C(n76), .Y(n1224) );
  NAND2X1 U91 ( .A(PLAINKEY[27]), .B(n246), .Y(n76) );
  OAI21X1 U93 ( .A(n241), .B(n1666), .C(n78), .Y(n1225) );
  NAND2X1 U94 ( .A(PLAINKEY[28]), .B(n246), .Y(n78) );
  OAI21X1 U96 ( .A(n242), .B(n1665), .C(n80), .Y(n1226) );
  NAND2X1 U97 ( .A(PLAINKEY[29]), .B(n245), .Y(n80) );
  OAI21X1 U99 ( .A(n242), .B(n1664), .C(n82), .Y(n1227) );
  NAND2X1 U100 ( .A(PLAINKEY[30]), .B(n245), .Y(n82) );
  OAI21X1 U102 ( .A(n243), .B(n1663), .C(n84), .Y(n1228) );
  NAND2X1 U103 ( .A(PLAINKEY[31]), .B(n245), .Y(n84) );
  OAI21X1 U105 ( .A(n243), .B(n1662), .C(n86), .Y(n1229) );
  NAND2X1 U106 ( .A(PLAINKEY[32]), .B(n245), .Y(n86) );
  OAI21X1 U108 ( .A(n242), .B(n1661), .C(n88), .Y(n1230) );
  NAND2X1 U109 ( .A(PLAINKEY[33]), .B(n245), .Y(n88) );
  OAI21X1 U111 ( .A(n243), .B(n1660), .C(n90), .Y(n1231) );
  NAND2X1 U112 ( .A(PLAINKEY[34]), .B(n245), .Y(n90) );
  OAI21X1 U114 ( .A(n242), .B(n1659), .C(n92), .Y(n1232) );
  NAND2X1 U115 ( .A(PLAINKEY[35]), .B(n245), .Y(n92) );
  OAI21X1 U117 ( .A(n242), .B(n1658), .C(n94), .Y(n1233) );
  NAND2X1 U118 ( .A(PLAINKEY[36]), .B(n245), .Y(n94) );
  OAI21X1 U120 ( .A(n243), .B(n1657), .C(n96), .Y(n1234) );
  NAND2X1 U121 ( .A(PLAINKEY[37]), .B(n245), .Y(n96) );
  OAI21X1 U123 ( .A(n243), .B(n1656), .C(n98), .Y(n1235) );
  NAND2X1 U124 ( .A(PLAINKEY[38]), .B(n245), .Y(n98) );
  OAI21X1 U126 ( .A(n243), .B(n1655), .C(n100), .Y(n1236) );
  NAND2X1 U127 ( .A(PLAINKEY[39]), .B(n245), .Y(n100) );
  OAI21X1 U129 ( .A(n243), .B(n1654), .C(n102), .Y(n1237) );
  NAND2X1 U130 ( .A(PLAINKEY[40]), .B(n245), .Y(n102) );
  OAI21X1 U132 ( .A(n243), .B(n1653), .C(n104), .Y(n1238) );
  NAND2X1 U133 ( .A(PLAINKEY[41]), .B(n245), .Y(n104) );
  OAI21X1 U135 ( .A(n242), .B(n1652), .C(n106), .Y(n1239) );
  NAND2X1 U136 ( .A(PLAINKEY[42]), .B(n245), .Y(n106) );
  OAI21X1 U138 ( .A(n243), .B(n1651), .C(n108), .Y(n1240) );
  NAND2X1 U139 ( .A(PLAINKEY[43]), .B(n245), .Y(n108) );
  OAI21X1 U141 ( .A(n243), .B(n1650), .C(n110), .Y(n1241) );
  NAND2X1 U142 ( .A(PLAINKEY[44]), .B(n244), .Y(n110) );
  OAI21X1 U144 ( .A(n243), .B(n1649), .C(n112), .Y(n1242) );
  NAND2X1 U145 ( .A(PLAINKEY[45]), .B(n244), .Y(n112) );
  OAI21X1 U147 ( .A(n243), .B(n1648), .C(n114), .Y(n1243) );
  NAND2X1 U148 ( .A(PLAINKEY[46]), .B(n245), .Y(n114) );
  OAI21X1 U150 ( .A(n240), .B(n1647), .C(n116), .Y(n1244) );
  NAND2X1 U151 ( .A(PLAINKEY[47]), .B(n244), .Y(n116) );
  OAI21X1 U153 ( .A(n242), .B(n1646), .C(n118), .Y(n1245) );
  NAND2X1 U154 ( .A(PLAINKEY[48]), .B(n244), .Y(n118) );
  OAI21X1 U156 ( .A(n242), .B(n1645), .C(n120), .Y(n1246) );
  NAND2X1 U157 ( .A(PLAINKEY[49]), .B(n244), .Y(n120) );
  OAI21X1 U159 ( .A(n242), .B(n1644), .C(n122), .Y(n1247) );
  NAND2X1 U160 ( .A(PLAINKEY[50]), .B(n244), .Y(n122) );
  OAI21X1 U162 ( .A(n241), .B(n1643), .C(n124), .Y(n1248) );
  NAND2X1 U163 ( .A(PLAINKEY[51]), .B(n244), .Y(n124) );
  OAI21X1 U165 ( .A(n242), .B(n1642), .C(n126), .Y(n1249) );
  NAND2X1 U166 ( .A(PLAINKEY[52]), .B(n244), .Y(n126) );
  OAI21X1 U168 ( .A(n241), .B(n1641), .C(n128), .Y(n1250) );
  NAND2X1 U169 ( .A(PLAINKEY[53]), .B(n244), .Y(n128) );
  OAI21X1 U171 ( .A(n241), .B(n1640), .C(n130), .Y(n1251) );
  NAND2X1 U172 ( .A(PLAINKEY[54]), .B(n244), .Y(n130) );
  OAI21X1 U174 ( .A(n240), .B(n1639), .C(n132), .Y(n1252) );
  NAND2X1 U175 ( .A(PLAINKEY[55]), .B(n245), .Y(n132) );
  OAI21X1 U177 ( .A(n241), .B(n1638), .C(n134), .Y(n1253) );
  NAND2X1 U178 ( .A(PLAINKEY[56]), .B(n244), .Y(n134) );
  OAI21X1 U180 ( .A(n240), .B(n1637), .C(n136), .Y(n1254) );
  NAND2X1 U181 ( .A(PLAINKEY[57]), .B(n244), .Y(n136) );
  OAI21X1 U183 ( .A(n240), .B(n1636), .C(n138), .Y(n1255) );
  NAND2X1 U184 ( .A(PLAINKEY[58]), .B(n244), .Y(n138) );
  OAI21X1 U186 ( .A(n240), .B(n1635), .C(n140), .Y(n1256) );
  NAND2X1 U187 ( .A(PLAINKEY[59]), .B(n244), .Y(n140) );
  OAI21X1 U188 ( .A(n239), .B(n1634), .C(n142), .Y(n1257) );
  NAND2X1 U189 ( .A(PLAINKEY[60]), .B(n244), .Y(n142) );
  OAI21X1 U191 ( .A(n239), .B(n1633), .C(n144), .Y(n1258) );
  NAND2X1 U192 ( .A(PLAINKEY[61]), .B(n244), .Y(n144) );
  OAI21X1 U194 ( .A(n239), .B(n1620), .C(n146), .Y(n1259) );
  NAND2X1 U195 ( .A(PLAINKEY[62]), .B(n244), .Y(n146) );
  OAI21X1 U196 ( .A(n239), .B(n1632), .C(n148), .Y(n1260) );
  NAND2X1 U197 ( .A(PLAINKEY[63]), .B(n245), .Y(n148) );
  NAND2X1 U1305 ( .A(n1584), .B(n1695), .Y(n1178) );
  keyreg_1_DW01_add_1 r577 ( .A(parityAccumulator), .B({RCV_DATA[7:3], n236, 
        n190, n189}), .CI(1'b0), .SUM({N1799, N1798, N1797, N1796, N1795, 
        N1794, N1793, N1792}) );
  INVX2 U3 ( .A(n191), .Y(n193) );
  BUFX2 U4 ( .A(n1503), .Y(n211) );
  INVX4 U5 ( .A(n31), .Y(n143) );
  INVX2 U7 ( .A(n835), .Y(n1080) );
  BUFX2 U8 ( .A(RCV_DATA[1]), .Y(n190) );
  INVX4 U23 ( .A(n67), .Y(n113) );
  INVX2 U26 ( .A(RCV_DATA[1]), .Y(n220) );
  AND2X2 U29 ( .A(n270), .B(n682), .Y(n1) );
  INVX1 U32 ( .A(n167), .Y(n168) );
  INVX1 U35 ( .A(n163), .Y(n164) );
  INVX2 U38 ( .A(n73), .Y(n1118) );
  INVX2 U41 ( .A(n81), .Y(n85) );
  INVX2 U44 ( .A(n169), .Y(n170) );
  INVX2 U47 ( .A(n1400), .Y(n169) );
  AND2X2 U50 ( .A(n1080), .B(n125), .Y(n2) );
  INVX1 U53 ( .A(n1130), .Y(n4) );
  INVX1 U56 ( .A(n894), .Y(n5) );
  INVX1 U59 ( .A(n628), .Y(n6) );
  INVX1 U62 ( .A(n1573), .Y(n7) );
  INVX2 U65 ( .A(n160), .Y(n1573) );
  BUFX2 U68 ( .A(n1394), .Y(n8) );
  INVX2 U71 ( .A(n256), .Y(n9) );
  BUFX4 U74 ( .A(state[2]), .Y(n159) );
  INVX2 U77 ( .A(n397), .Y(n10) );
  NAND2X1 U80 ( .A(n156), .B(n150), .Y(n11) );
  BUFX2 U83 ( .A(n1600), .Y(n14) );
  BUFX2 U86 ( .A(n1511), .Y(n16) );
  OR2X2 U89 ( .A(n139), .B(n1574), .Y(n17) );
  OR2X1 U92 ( .A(n139), .B(n1574), .Y(n1599) );
  OR2X2 U95 ( .A(n159), .B(n1573), .Y(n139) );
  BUFX2 U98 ( .A(n1503), .Y(n19) );
  BUFX2 U101 ( .A(n1503), .Y(n20) );
  NAND2X1 U104 ( .A(RCV_DATA[6]), .B(n223), .Y(n21) );
  BUFX4 U107 ( .A(n1527), .Y(n223) );
  INVX2 U110 ( .A(n378), .Y(n348) );
  NAND3X1 U113 ( .A(n1553), .B(n1593), .C(n267), .Y(n23) );
  OR2X2 U116 ( .A(n1400), .B(n191), .Y(n450) );
  INVX4 U119 ( .A(address[3]), .Y(n191) );
  INVX2 U122 ( .A(n1420), .Y(n25) );
  NOR2X1 U125 ( .A(address[6]), .B(address[7]), .Y(n27) );
  NOR2X1 U128 ( .A(address[6]), .B(address[7]), .Y(n29) );
  AND2X2 U131 ( .A(n266), .B(n1600), .Y(n267) );
  OR2X2 U134 ( .A(n835), .B(n192), .Y(n31) );
  AND2X2 U137 ( .A(n935), .B(n1007), .Y(n33) );
  INVX1 U140 ( .A(n33), .Y(n987) );
  AND2X2 U143 ( .A(n902), .B(n975), .Y(n35) );
  INVX1 U146 ( .A(n35), .Y(n955) );
  AND2X2 U149 ( .A(n438), .B(n510), .Y(n37) );
  INVX1 U152 ( .A(n37), .Y(n490) );
  INVX1 U155 ( .A(n477), .Y(n496) );
  AND2X2 U158 ( .A(n372), .B(n444), .Y(n39) );
  INVX1 U161 ( .A(n39), .Y(n424) );
  AND2X1 U164 ( .A(n1599), .B(n1578), .Y(n41) );
  AND2X2 U167 ( .A(n271), .B(n286), .Y(n43) );
  INVX1 U170 ( .A(n43), .Y(n1081) );
  NAND3X1 U173 ( .A(n1553), .B(n11), .C(n267), .Y(n45) );
  INVX2 U176 ( .A(n1548), .Y(n47) );
  AND2X2 U179 ( .A(n769), .B(n844), .Y(n49) );
  INVX1 U182 ( .A(n49), .Y(n823) );
  INVX4 U185 ( .A(n379), .Y(n51) );
  BUFX2 U190 ( .A(n161), .Y(n235) );
  AND2X2 U193 ( .A(n107), .B(n109), .Y(n53) );
  AND2X2 U198 ( .A(n111), .B(n1405), .Y(n55) );
  INVX1 U199 ( .A(n55), .Y(n1447) );
  AND2X2 U200 ( .A(n1033), .B(n1110), .Y(n57) );
  INVX1 U201 ( .A(n57), .Y(n1089) );
  AND2X2 U202 ( .A(n504), .B(n578), .Y(n59) );
  INVX1 U203 ( .A(n59), .Y(n557) );
  INVX2 U204 ( .A(n1151), .Y(n61) );
  INVX1 U205 ( .A(n61), .Y(n63) );
  INVX4 U206 ( .A(n152), .Y(n166) );
  BUFX4 U207 ( .A(n1503), .Y(n213) );
  INVX1 U208 ( .A(n447), .Y(n65) );
  INVX4 U209 ( .A(n69), .Y(n135) );
  OR2X2 U210 ( .A(n1514), .B(n192), .Y(n67) );
  INVX2 U211 ( .A(n1514), .Y(n1495) );
  OR2X2 U212 ( .A(n268), .B(n45), .Y(n69) );
  INVX1 U213 ( .A(n369), .Y(n107) );
  INVX1 U214 ( .A(n1398), .Y(n1399) );
  INVX4 U215 ( .A(n332), .Y(n415) );
  AND2X2 U216 ( .A(n1067), .B(n1145), .Y(n71) );
  INVX1 U217 ( .A(n71), .Y(n1124) );
  AND2X2 U218 ( .A(n189), .B(n1420), .Y(n73) );
  INVX1 U219 ( .A(n1371), .Y(n1394) );
  AND2X2 U220 ( .A(n803), .B(n876), .Y(n75) );
  INVX1 U221 ( .A(n75), .Y(n856) );
  AND2X2 U222 ( .A(n537), .B(n610), .Y(n77) );
  INVX1 U223 ( .A(n77), .Y(n590) );
  AND2X2 U224 ( .A(n1365), .B(n1383), .Y(n79) );
  INVX1 U225 ( .A(n79), .Y(n1427) );
  INVX4 U226 ( .A(n1438), .Y(n1504) );
  INVX4 U227 ( .A(n372), .Y(n447) );
  MUX2X1 U228 ( .B(n208), .A(n1430), .S(n1380), .Y(n1432) );
  INVX2 U229 ( .A(state[1]), .Y(n81) );
  INVX1 U230 ( .A(n81), .Y(n83) );
  NAND2X1 U231 ( .A(n306), .B(n135), .Y(n87) );
  INVX4 U232 ( .A(n87), .Y(n162) );
  INVX1 U233 ( .A(n204), .Y(n199) );
  OR2X2 U234 ( .A(n1545), .B(n1580), .Y(n1546) );
  INVX2 U235 ( .A(n1545), .Y(n1542) );
  INVX4 U236 ( .A(n1116), .Y(n1420) );
  AND2X2 U237 ( .A(n202), .B(n348), .Y(n303) );
  INVX4 U238 ( .A(n1458), .Y(n1528) );
  INVX1 U239 ( .A(n17), .Y(n1549) );
  INVX8 U240 ( .A(n200), .Y(n198) );
  AND2X2 U241 ( .A(n154), .B(address[0]), .Y(n152) );
  AND2X2 U242 ( .A(n154), .B(n283), .Y(n89) );
  INVX2 U243 ( .A(n89), .Y(n1185) );
  AND2X2 U244 ( .A(n838), .B(n908), .Y(n91) );
  INVX1 U245 ( .A(n91), .Y(n888) );
  INVX1 U246 ( .A(n1545), .Y(n1544) );
  BUFX4 U247 ( .A(n162), .Y(n103) );
  INVX4 U248 ( .A(n119), .Y(n195) );
  INVX4 U249 ( .A(n119), .Y(n196) );
  AND2X2 U250 ( .A(n89), .B(n193), .Y(n93) );
  INVX2 U251 ( .A(n93), .Y(n1513) );
  BUFX2 U252 ( .A(n1608), .Y(n158) );
  BUFX4 U253 ( .A(n1608), .Y(n157) );
  BUFX4 U254 ( .A(n1527), .Y(n222) );
  BUFX4 U255 ( .A(n1527), .Y(n225) );
  AND2X2 U256 ( .A(n83), .B(n159), .Y(n153) );
  INVX4 U257 ( .A(n322), .Y(n1503) );
  INVX1 U258 ( .A(n911), .Y(n95) );
  INVX1 U259 ( .A(n85), .Y(n259) );
  AND2X2 U260 ( .A(n1104), .B(n1179), .Y(n97) );
  INVX1 U261 ( .A(n97), .Y(n1158) );
  AND2X2 U262 ( .A(n572), .B(n642), .Y(n99) );
  INVX1 U263 ( .A(n99), .Y(n622) );
  INVX1 U264 ( .A(n364), .Y(n382) );
  INVX1 U265 ( .A(n14), .Y(n1587) );
  OR2X2 U266 ( .A(n370), .B(n369), .Y(n117) );
  NAND2X1 U267 ( .A(n147), .B(n260), .Y(n101) );
  BUFX2 U268 ( .A(n162), .Y(n105) );
  BUFX4 U269 ( .A(n1503), .Y(n212) );
  AND2X1 U270 ( .A(n41), .B(n302), .Y(n109) );
  INVX2 U271 ( .A(n1), .Y(n165) );
  AND2X1 U272 ( .A(n151), .B(n1101), .Y(n141) );
  INVX4 U273 ( .A(RCV_DATA[2]), .Y(n238) );
  INVX2 U274 ( .A(n249), .Y(n242) );
  INVX2 U275 ( .A(n249), .Y(n241) );
  INVX2 U276 ( .A(n248), .Y(n240) );
  INVX2 U277 ( .A(n248), .Y(n239) );
  INVX2 U278 ( .A(n250), .Y(n243) );
  INVX2 U279 ( .A(n251), .Y(n244) );
  INVX2 U280 ( .A(n251), .Y(n245) );
  INVX2 U281 ( .A(n252), .Y(n246) );
  INVX2 U282 ( .A(n250), .Y(n247) );
  BUFX2 U283 ( .A(n1510), .Y(n219) );
  AND2X2 U284 ( .A(n1399), .B(n223), .Y(n111) );
  BUFX2 U285 ( .A(n255), .Y(n250) );
  BUFX2 U286 ( .A(n254), .Y(n251) );
  BUFX2 U287 ( .A(n255), .Y(n249) );
  BUFX2 U288 ( .A(n255), .Y(n248) );
  BUFX2 U289 ( .A(n254), .Y(n252) );
  BUFX2 U290 ( .A(n254), .Y(n253) );
  INVX2 U291 ( .A(n275), .Y(n360) );
  INVX2 U292 ( .A(n117), .Y(n205) );
  INVX2 U293 ( .A(n117), .Y(n206) );
  AND2X2 U294 ( .A(n125), .B(n1495), .Y(n115) );
  INVX2 U295 ( .A(n117), .Y(n207) );
  INVX2 U296 ( .A(RST), .Y(n254) );
  INVX2 U297 ( .A(RST), .Y(n255) );
  BUFX2 U298 ( .A(n162), .Y(n209) );
  BUFX2 U299 ( .A(n162), .Y(n210) );
  AND2X2 U300 ( .A(n367), .B(n135), .Y(n119) );
  AND2X2 U301 ( .A(n1420), .B(n193), .Y(n121) );
  AND2X2 U302 ( .A(n61), .B(n193), .Y(n123) );
  AND2X2 U303 ( .A(n167), .B(n193), .Y(n125) );
  AND2X2 U304 ( .A(n163), .B(n193), .Y(n127) );
  INVX2 U305 ( .A(RCV_DATA[1]), .Y(n221) );
  AND2X2 U306 ( .A(n550), .B(n1101), .Y(n129) );
  AND2X2 U307 ( .A(n193), .B(n43), .Y(n131) );
  AND2X2 U308 ( .A(n152), .B(n193), .Y(n133) );
  INVX2 U309 ( .A(n171), .Y(n172) );
  INVX2 U310 ( .A(n171), .Y(n173) );
  AND2X2 U311 ( .A(n284), .B(n121), .Y(n137) );
  INVX2 U312 ( .A(n141), .Y(n186) );
  INVX2 U313 ( .A(n141), .Y(n187) );
  BUFX2 U314 ( .A(n1503), .Y(n214) );
  INVX2 U315 ( .A(n238), .Y(n236) );
  INVX2 U316 ( .A(n533), .Y(n171) );
  AND2X2 U317 ( .A(n816), .B(n1101), .Y(n145) );
  AND2X2 U318 ( .A(n159), .B(n81), .Y(n147) );
  INVX2 U319 ( .A(n174), .Y(n175) );
  INVX2 U320 ( .A(n174), .Y(n176) );
  INVX2 U321 ( .A(n180), .Y(n181) );
  INVX2 U322 ( .A(n180), .Y(n182) );
  INVX2 U323 ( .A(n177), .Y(n178) );
  INVX2 U324 ( .A(n183), .Y(n184) );
  INVX2 U325 ( .A(n177), .Y(n179) );
  INVX2 U326 ( .A(n183), .Y(n185) );
  INVX2 U327 ( .A(n238), .Y(n237) );
  NOR2X1 U328 ( .A(n160), .B(n194), .Y(n149) );
  AND2X2 U329 ( .A(n194), .B(n1573), .Y(n150) );
  INVX2 U330 ( .A(n191), .Y(n192) );
  INVX2 U331 ( .A(n1476), .Y(n167) );
  INVX2 U332 ( .A(n1440), .Y(n163) );
  INVX2 U333 ( .A(n665), .Y(n174) );
  INVX2 U334 ( .A(n931), .Y(n180) );
  INVX2 U335 ( .A(n799), .Y(n177) );
  INVX2 U336 ( .A(n1063), .Y(n183) );
  AND2X2 U337 ( .A(address[4]), .B(address[5]), .Y(n151) );
  INVX4 U338 ( .A(n188), .Y(n189) );
  INVX2 U339 ( .A(RCV_DATA[0]), .Y(n188) );
  AND2X2 U340 ( .A(address[1]), .B(address[2]), .Y(n154) );
  NOR2X1 U341 ( .A(address[6]), .B(address[7]), .Y(n155) );
  NOR2X1 U342 ( .A(n85), .B(n159), .Y(n156) );
  BUFX4 U343 ( .A(state[0]), .Y(n194) );
  BUFX4 U344 ( .A(state[3]), .Y(n160) );
  INVX4 U345 ( .A(n333), .Y(n1527) );
  BUFX2 U346 ( .A(n53), .Y(n204) );
  BUFX2 U347 ( .A(n53), .Y(n203) );
  BUFX2 U348 ( .A(n53), .Y(n201) );
  AND2X2 U349 ( .A(RCV_DATA[7]), .B(n223), .Y(n161) );
  INVX1 U350 ( .A(n161), .Y(n379) );
  INVX2 U351 ( .A(n162), .Y(n1439) );
  INVX1 U352 ( .A(n1593), .Y(n1548) );
  MUX2X1 U353 ( .B(n1439), .A(n307), .S(n275), .Y(n308) );
  INVX4 U354 ( .A(n298), .Y(n550) );
  INVX4 U355 ( .A(n569), .Y(n816) );
  INVX8 U356 ( .A(n202), .Y(n197) );
  BUFX4 U357 ( .A(n53), .Y(n200) );
  BUFX4 U358 ( .A(n53), .Y(n202) );
  BUFX4 U359 ( .A(n162), .Y(n208) );
  BUFX4 U360 ( .A(n1510), .Y(n215) );
  BUFX4 U361 ( .A(n1510), .Y(n216) );
  BUFX4 U362 ( .A(n1510), .Y(n217) );
  BUFX4 U363 ( .A(n1510), .Y(n218) );
  BUFX4 U364 ( .A(n1527), .Y(n224) );
  INVX8 U365 ( .A(n228), .Y(n226) );
  INVX8 U366 ( .A(n228), .Y(n227) );
  BUFX4 U367 ( .A(n1529), .Y(n228) );
  BUFX4 U368 ( .A(n21), .Y(n229) );
  BUFX4 U369 ( .A(n21), .Y(n230) );
  BUFX4 U370 ( .A(n161), .Y(n231) );
  BUFX4 U371 ( .A(n161), .Y(n232) );
  BUFX4 U372 ( .A(n161), .Y(n233) );
  BUFX4 U373 ( .A(n161), .Y(n234) );
  NOR2X1 U374 ( .A(n160), .B(n194), .Y(n257) );
  INVX2 U375 ( .A(n159), .Y(n256) );
  NAND3X1 U376 ( .A(n257), .B(n85), .C(n256), .Y(n1608) );
  NOR2X1 U377 ( .A(n160), .B(n259), .Y(n258) );
  NAND3X1 U378 ( .A(n9), .B(n194), .C(n258), .Y(n1578) );
  NAND2X1 U379 ( .A(n158), .B(n1578), .Y(CLR_RBUFF) );
  NOR2X1 U380 ( .A(n160), .B(n194), .Y(n260) );
  NAND2X1 U381 ( .A(n147), .B(n260), .Y(n1553) );
  INVX2 U382 ( .A(n101), .Y(PROG_ERROR) );
  NAND2X1 U383 ( .A(n153), .B(n260), .Y(n1597) );
  NAND2X1 U384 ( .A(n1597), .B(n1553), .Y(n264) );
  INVX2 U385 ( .A(n194), .Y(n261) );
  NAND2X1 U386 ( .A(n156), .B(n261), .Y(n1598) );
  NOR2X1 U387 ( .A(n160), .B(n159), .Y(n262) );
  NAND3X1 U388 ( .A(n85), .B(n194), .C(n262), .Y(n1600) );
  OAI21X1 U389 ( .A(n7), .B(n1598), .C(n1600), .Y(n263) );
  NOR3X1 U390 ( .A(n264), .B(CLR_RBUFF), .C(n263), .Y(n1535) );
  OR2X2 U391 ( .A(n83), .B(n194), .Y(n1574) );
  NAND2X1 U392 ( .A(n150), .B(n147), .Y(n1605) );
  INVX2 U393 ( .A(n1605), .Y(n1583) );
  NAND2X1 U394 ( .A(n156), .B(n150), .Y(n1593) );
  AOI21X1 U395 ( .A(n1583), .B(parityError), .C(n1548), .Y(n265) );
  NAND3X1 U396 ( .A(n1535), .B(n17), .C(n265), .Y(KEY_ERROR) );
  INVX2 U397 ( .A(currentPlainKey[63]), .Y(n1632) );
  INVX2 U398 ( .A(currentPlainKey[62]), .Y(n1620) );
  INVX2 U399 ( .A(currentPlainKey[3]), .Y(n1691) );
  INVX2 U400 ( .A(currentPlainKey[2]), .Y(n1692) );
  INVX2 U401 ( .A(currentPlainKey[1]), .Y(n1693) );
  INVX2 U402 ( .A(currentPlainKey[0]), .Y(n1694) );
  INVX2 U403 ( .A(parityAccumulator[4]), .Y(n1627) );
  INVX2 U404 ( .A(parityAccumulator[5]), .Y(n1628) );
  NAND2X1 U405 ( .A(n1599), .B(n1578), .Y(n268) );
  AOI21X1 U406 ( .A(n149), .B(n153), .C(n243), .Y(n266) );
  NAND3X1 U407 ( .A(n1593), .B(n1553), .C(n267), .Y(n369) );
  NAND2X1 U408 ( .A(n135), .B(n1605), .Y(n1510) );
  NAND2X1 U409 ( .A(n219), .B(currentPlainKey[0]), .Y(n292) );
  NAND3X1 U410 ( .A(address[6]), .B(address[7]), .C(n151), .Y(n288) );
  INVX2 U411 ( .A(n288), .Y(n284) );
  INVX2 U412 ( .A(address[0]), .Y(n283) );
  INVX2 U413 ( .A(address[1]), .Y(n287) );
  NAND3X1 U414 ( .A(address[2]), .B(n283), .C(n287), .Y(n1151) );
  NAND2X1 U415 ( .A(n284), .B(n123), .Y(n269) );
  INVX2 U416 ( .A(n269), .Y(n344) );
  INVX2 U417 ( .A(RCV_DATA[4]), .Y(n305) );
  NAND2X1 U418 ( .A(n344), .B(n305), .Y(n282) );
  NAND2X1 U419 ( .A(n284), .B(n93), .Y(n378) );
  INVX2 U420 ( .A(address[2]), .Y(n286) );
  NAND3X1 U421 ( .A(address[0]), .B(address[1]), .C(n286), .Y(n1440) );
  NAND2X1 U422 ( .A(n284), .B(n127), .Y(n294) );
  NAND2X1 U423 ( .A(n294), .B(n269), .Y(n296) );
  AOI21X1 U424 ( .A(n348), .B(n236), .C(n296), .Y(n278) );
  NOR2X1 U425 ( .A(address[4]), .B(n192), .Y(n270) );
  INVX2 U426 ( .A(address[5]), .Y(n682) );
  INVX2 U427 ( .A(n165), .Y(n314) );
  NOR2X1 U428 ( .A(address[1]), .B(address[0]), .Y(n271) );
  NAND2X1 U429 ( .A(n314), .B(n43), .Y(n272) );
  NAND2X1 U430 ( .A(n189), .B(n43), .Y(n1083) );
  INVX2 U431 ( .A(n1083), .Y(n1378) );
  AOI22X1 U432 ( .A(n272), .B(currentPlainKey[0]), .C(n314), .D(n1378), .Y(
        n274) );
  NAND2X1 U433 ( .A(n284), .B(n133), .Y(n331) );
  NAND2X1 U434 ( .A(n378), .B(n331), .Y(n364) );
  INVX2 U435 ( .A(n331), .Y(n397) );
  NAND2X1 U436 ( .A(n397), .B(n190), .Y(n273) );
  OAI21X1 U437 ( .A(n274), .B(n364), .C(n273), .Y(n276) );
  NAND3X1 U438 ( .A(address[0]), .B(address[2]), .C(n287), .Y(n1476) );
  NAND2X1 U439 ( .A(n284), .B(n125), .Y(n275) );
  MUX2X1 U440 ( .B(n276), .A(RCV_DATA[3]), .S(n360), .Y(n277) );
  NAND2X1 U441 ( .A(n278), .B(n277), .Y(n281) );
  INVX2 U442 ( .A(n294), .Y(n327) );
  OR2X2 U443 ( .A(n23), .B(n158), .Y(n333) );
  INVX2 U444 ( .A(n158), .Y(n1596) );
  NAND2X1 U445 ( .A(n1596), .B(RCV_DATA[5]), .Y(n279) );
  OR2X2 U446 ( .A(n369), .B(n279), .Y(n322) );
  OAI21X1 U447 ( .A(n327), .B(n333), .C(n322), .Y(n280) );
  NAND3X1 U448 ( .A(n282), .B(n281), .C(n280), .Y(n285) );
  NAND2X1 U449 ( .A(RCV_DATA[6]), .B(n223), .Y(n1529) );
  NAND3X1 U450 ( .A(address[1]), .B(n283), .C(n286), .Y(n1116) );
  MUX2X1 U451 ( .B(n285), .A(n229), .S(n137), .Y(n290) );
  NAND3X1 U452 ( .A(address[0]), .B(n287), .C(n286), .Y(n1400) );
  NOR2X1 U453 ( .A(n450), .B(n288), .Y(n289) );
  MUX2X1 U454 ( .B(n290), .A(n232), .S(n289), .Y(n291) );
  NAND2X1 U455 ( .A(n292), .B(n291), .Y(n1332) );
  NAND2X1 U456 ( .A(n219), .B(currentPlainKey[1]), .Y(n313) );
  INVX2 U457 ( .A(RCV_DATA[6]), .Y(n293) );
  NOR2X1 U458 ( .A(n294), .B(n293), .Y(n295) );
  AOI22X1 U459 ( .A(n344), .B(n214), .C(n295), .D(n222), .Y(n310) );
  INVX2 U460 ( .A(n296), .Y(n324) );
  NAND2X1 U461 ( .A(n189), .B(n169), .Y(n1402) );
  OAI21X1 U462 ( .A(n170), .B(n165), .C(currentPlainKey[1]), .Y(n297) );
  OAI21X1 U463 ( .A(n1402), .B(n165), .C(n297), .Y(n299) );
  INVX2 U464 ( .A(address[4]), .Y(n948) );
  NAND3X1 U465 ( .A(n27), .B(n948), .C(n682), .Y(n298) );
  INVX2 U466 ( .A(n192), .Y(n1101) );
  NAND2X1 U467 ( .A(n129), .B(n43), .Y(n332) );
  MUX2X1 U468 ( .B(n299), .A(n190), .S(n415), .Y(n301) );
  NAND2X1 U469 ( .A(n397), .B(n236), .Y(n300) );
  OAI21X1 U470 ( .A(n364), .B(n301), .C(n300), .Y(n304) );
  INVX2 U471 ( .A(RCV_DATA[3]), .Y(n1520) );
  NOR2X1 U472 ( .A(n1520), .B(n157), .Y(n302) );
  AOI21X1 U473 ( .A(n222), .B(n304), .C(n303), .Y(n307) );
  NOR2X1 U474 ( .A(n305), .B(n157), .Y(n306) );
  NAND2X1 U475 ( .A(n324), .B(n308), .Y(n309) );
  NAND2X1 U476 ( .A(n310), .B(n309), .Y(n311) );
  MUX2X1 U477 ( .B(n311), .A(n234), .S(n137), .Y(n312) );
  NAND2X1 U478 ( .A(n312), .B(n313), .Y(n1331) );
  NOR2X1 U479 ( .A(n1439), .B(n378), .Y(n326) );
  NAND2X1 U480 ( .A(n314), .B(n1420), .Y(n315) );
  AOI22X1 U481 ( .A(n315), .B(currentPlainKey[2]), .C(n314), .D(n73), .Y(n317)
         );
  NAND2X1 U482 ( .A(n129), .B(n169), .Y(n411) );
  NAND2X1 U483 ( .A(n332), .B(n411), .Y(n391) );
  INVX2 U484 ( .A(n411), .Y(n430) );
  NAND2X1 U485 ( .A(n430), .B(n190), .Y(n316) );
  OAI21X1 U486 ( .A(n317), .B(n391), .C(n316), .Y(n319) );
  NOR2X1 U487 ( .A(n238), .B(n332), .Y(n318) );
  AOI21X1 U488 ( .A(n319), .B(n10), .C(n318), .Y(n320) );
  OAI22X1 U489 ( .A(n320), .B(n333), .C(n197), .D(n10), .Y(n321) );
  NAND2X1 U490 ( .A(n321), .B(n378), .Y(n323) );
  MUX2X1 U491 ( .B(n323), .A(n322), .S(n360), .Y(n325) );
  OAI21X1 U492 ( .A(n326), .B(n325), .C(n324), .Y(n330) );
  NAND2X1 U493 ( .A(n344), .B(n227), .Y(n329) );
  AOI22X1 U494 ( .A(n327), .B(n231), .C(n219), .D(currentPlainKey[2]), .Y(n328) );
  NAND3X1 U495 ( .A(n330), .B(n329), .C(n328), .Y(n1330) );
  NAND2X1 U496 ( .A(n219), .B(currentPlainKey[3]), .Y(n347) );
  NOR2X1 U497 ( .A(n1439), .B(n10), .Y(n342) );
  NAND2X1 U498 ( .A(n189), .B(n163), .Y(n1135) );
  OAI21X1 U499 ( .A(n164), .B(n165), .C(currentPlainKey[3]), .Y(n334) );
  OAI21X1 U500 ( .A(n1135), .B(n165), .C(n334), .Y(n335) );
  NAND2X1 U501 ( .A(n129), .B(n1420), .Y(n372) );
  MUX2X1 U502 ( .B(n335), .A(n190), .S(n447), .Y(n337) );
  NAND2X1 U503 ( .A(n430), .B(n237), .Y(n336) );
  OAI21X1 U504 ( .A(n337), .B(n391), .C(n336), .Y(n338) );
  AOI22X1 U505 ( .A(n415), .B(n203), .C(n338), .D(n225), .Y(n340) );
  NAND2X1 U506 ( .A(n348), .B(n211), .Y(n339) );
  OAI21X1 U507 ( .A(n340), .B(n364), .C(n339), .Y(n341) );
  NOR2X1 U508 ( .A(n342), .B(n341), .Y(n343) );
  MUX2X1 U509 ( .B(n343), .A(n229), .S(n360), .Y(n345) );
  MUX2X1 U510 ( .B(n345), .A(n233), .S(n344), .Y(n346) );
  NAND2X1 U511 ( .A(n347), .B(n346), .Y(n1329) );
  AOI22X1 U512 ( .A(n348), .B(n227), .C(currentPlainKey[4]), .D(n219), .Y(n363) );
  NAND2X1 U513 ( .A(n129), .B(n163), .Y(n444) );
  NAND2X1 U514 ( .A(n189), .B(n61), .Y(n1455) );
  OAI21X1 U515 ( .A(n63), .B(n165), .C(currentPlainKey[4]), .Y(n349) );
  OAI21X1 U516 ( .A(n1455), .B(n165), .C(n349), .Y(n351) );
  NOR2X1 U517 ( .A(n221), .B(n444), .Y(n350) );
  AOI21X1 U518 ( .A(n39), .B(n351), .C(n350), .Y(n353) );
  NAND2X1 U519 ( .A(n447), .B(n237), .Y(n352) );
  OAI21X1 U520 ( .A(n430), .B(n353), .C(n352), .Y(n354) );
  NAND2X1 U521 ( .A(n222), .B(n354), .Y(n356) );
  NAND2X1 U522 ( .A(n430), .B(n201), .Y(n355) );
  AOI21X1 U523 ( .A(n356), .B(n355), .C(n364), .Y(n357) );
  MUX2X1 U524 ( .B(n357), .A(n208), .S(n415), .Y(n359) );
  NAND2X1 U525 ( .A(n397), .B(n20), .Y(n358) );
  NAND2X1 U526 ( .A(n359), .B(n358), .Y(n361) );
  MUX2X1 U527 ( .B(n361), .A(n51), .S(n360), .Y(n362) );
  NAND2X1 U528 ( .A(n362), .B(n363), .Y(n1328) );
  NAND2X1 U529 ( .A(n430), .B(n210), .Y(n377) );
  NAND2X1 U530 ( .A(n189), .B(n167), .Y(n1478) );
  OAI21X1 U531 ( .A(n168), .B(n165), .C(currentPlainKey[5]), .Y(n365) );
  OAI21X1 U532 ( .A(n1478), .B(n165), .C(n365), .Y(n366) );
  NAND3X1 U533 ( .A(n39), .B(n222), .C(n366), .Y(n368) );
  NOR2X1 U534 ( .A(n220), .B(n157), .Y(n367) );
  NAND2X1 U535 ( .A(n129), .B(n61), .Y(n405) );
  INVX2 U536 ( .A(n405), .Y(n481) );
  MUX2X1 U537 ( .B(n368), .A(n195), .S(n481), .Y(n374) );
  INVX2 U538 ( .A(n444), .Y(n463) );
  NAND2X1 U539 ( .A(n1596), .B(n237), .Y(n370) );
  NAND2X1 U540 ( .A(n463), .B(n205), .Y(n371) );
  OAI21X1 U541 ( .A(n199), .B(n65), .C(n371), .Y(n373) );
  INVX2 U542 ( .A(n391), .Y(n414) );
  OAI21X1 U543 ( .A(n374), .B(n373), .C(n414), .Y(n376) );
  NAND2X1 U544 ( .A(n415), .B(n212), .Y(n375) );
  NAND3X1 U545 ( .A(n377), .B(n376), .C(n375), .Y(n381) );
  NOR2X1 U546 ( .A(n379), .B(n378), .Y(n380) );
  AOI21X1 U547 ( .A(n382), .B(n381), .C(n380), .Y(n384) );
  AOI22X1 U548 ( .A(n397), .B(n226), .C(currentPlainKey[5]), .D(n219), .Y(n383) );
  NAND2X1 U549 ( .A(n384), .B(n383), .Y(n1327) );
  AOI22X1 U550 ( .A(n415), .B(n226), .C(currentPlainKey[6]), .D(n219), .Y(n400) );
  NAND2X1 U551 ( .A(n129), .B(n167), .Y(n477) );
  NAND2X1 U552 ( .A(n405), .B(n477), .Y(n457) );
  INVX2 U553 ( .A(n457), .Y(n480) );
  NAND2X1 U554 ( .A(n189), .B(n89), .Y(n1490) );
  OAI21X1 U555 ( .A(n1185), .B(n165), .C(currentPlainKey[6]), .Y(n385) );
  OAI21X1 U556 ( .A(n1490), .B(n165), .C(n385), .Y(n387) );
  NOR2X1 U557 ( .A(n220), .B(n477), .Y(n386) );
  AOI21X1 U558 ( .A(n480), .B(n387), .C(n386), .Y(n389) );
  NAND2X1 U559 ( .A(n481), .B(n237), .Y(n388) );
  OAI21X1 U560 ( .A(n463), .B(n389), .C(n388), .Y(n390) );
  NAND2X1 U561 ( .A(n222), .B(n390), .Y(n393) );
  NAND2X1 U562 ( .A(n463), .B(n200), .Y(n392) );
  AOI21X1 U563 ( .A(n393), .B(n392), .C(n391), .Y(n394) );
  MUX2X1 U564 ( .B(n394), .A(n209), .S(n447), .Y(n396) );
  NAND2X1 U565 ( .A(n430), .B(n214), .Y(n395) );
  NAND2X1 U566 ( .A(n396), .B(n395), .Y(n398) );
  MUX2X1 U567 ( .B(n398), .A(n234), .S(n397), .Y(n399) );
  NAND2X1 U568 ( .A(n400), .B(n399), .Y(n1326) );
  NAND2X1 U569 ( .A(n463), .B(n210), .Y(n410) );
  NAND2X1 U570 ( .A(n189), .B(n152), .Y(n1361) );
  OAI21X1 U571 ( .A(n166), .B(n165), .C(currentPlainKey[7]), .Y(n401) );
  OAI21X1 U572 ( .A(n1361), .B(n165), .C(n401), .Y(n402) );
  NAND3X1 U573 ( .A(n480), .B(n225), .C(n402), .Y(n403) );
  NAND2X1 U574 ( .A(n129), .B(n89), .Y(n438) );
  INVX2 U575 ( .A(n438), .Y(n513) );
  MUX2X1 U576 ( .B(n403), .A(n195), .S(n513), .Y(n407) );
  NAND2X1 U577 ( .A(n496), .B(n205), .Y(n404) );
  OAI21X1 U578 ( .A(n198), .B(n405), .C(n404), .Y(n406) );
  OAI21X1 U579 ( .A(n407), .B(n406), .C(n39), .Y(n409) );
  NAND2X1 U580 ( .A(n447), .B(n20), .Y(n408) );
  NAND3X1 U581 ( .A(n410), .B(n409), .C(n408), .Y(n413) );
  NOR2X1 U582 ( .A(n230), .B(n411), .Y(n412) );
  AOI21X1 U583 ( .A(n414), .B(n413), .C(n412), .Y(n417) );
  AOI22X1 U584 ( .A(n415), .B(n235), .C(currentPlainKey[7]), .D(n219), .Y(n416) );
  NAND2X1 U585 ( .A(n417), .B(n416), .Y(n1325) );
  AOI22X1 U586 ( .A(n447), .B(n227), .C(currentPlainKey[8]), .D(n219), .Y(n433) );
  NAND2X1 U587 ( .A(n129), .B(n152), .Y(n510) );
  NAND3X1 U588 ( .A(n192), .B(n948), .C(n682), .Y(n533) );
  OAI21X1 U589 ( .A(n1081), .B(n172), .C(currentPlainKey[8]), .Y(n418) );
  OAI21X1 U590 ( .A(n1083), .B(n173), .C(n418), .Y(n420) );
  NOR2X1 U591 ( .A(n220), .B(n510), .Y(n419) );
  AOI21X1 U592 ( .A(n37), .B(n420), .C(n419), .Y(n422) );
  NAND2X1 U593 ( .A(n513), .B(n237), .Y(n421) );
  OAI21X1 U594 ( .A(n496), .B(n422), .C(n421), .Y(n423) );
  NAND2X1 U595 ( .A(n222), .B(n423), .Y(n426) );
  NAND2X1 U596 ( .A(n496), .B(n201), .Y(n425) );
  AOI21X1 U597 ( .A(n426), .B(n425), .C(n424), .Y(n427) );
  MUX2X1 U598 ( .B(n427), .A(n210), .S(n481), .Y(n429) );
  NAND2X1 U599 ( .A(n463), .B(n20), .Y(n428) );
  NAND2X1 U600 ( .A(n429), .B(n428), .Y(n431) );
  MUX2X1 U601 ( .B(n431), .A(n233), .S(n430), .Y(n432) );
  NAND2X1 U602 ( .A(n433), .B(n432), .Y(n1324) );
  NAND2X1 U603 ( .A(n496), .B(n105), .Y(n443) );
  OAI21X1 U604 ( .A(n170), .B(n172), .C(currentPlainKey[9]), .Y(n434) );
  OAI21X1 U605 ( .A(n1402), .B(n173), .C(n434), .Y(n435) );
  NAND3X1 U606 ( .A(n37), .B(n224), .C(n435), .Y(n436) );
  NAND2X1 U607 ( .A(n550), .B(n131), .Y(n471) );
  INVX2 U608 ( .A(n471), .Y(n547) );
  MUX2X1 U609 ( .B(n436), .A(n196), .S(n547), .Y(n440) );
  INVX2 U610 ( .A(n510), .Y(n528) );
  NAND2X1 U611 ( .A(n528), .B(n205), .Y(n437) );
  OAI21X1 U612 ( .A(n198), .B(n438), .C(n437), .Y(n439) );
  OAI21X1 U613 ( .A(n440), .B(n439), .C(n480), .Y(n442) );
  NAND2X1 U614 ( .A(n481), .B(n212), .Y(n441) );
  NAND3X1 U615 ( .A(n443), .B(n442), .C(n441), .Y(n446) );
  NOR2X1 U616 ( .A(n230), .B(n444), .Y(n445) );
  AOI21X1 U617 ( .A(n39), .B(n446), .C(n445), .Y(n449) );
  AOI22X1 U618 ( .A(n447), .B(n235), .C(currentPlainKey[9]), .D(n218), .Y(n448) );
  NAND2X1 U619 ( .A(n449), .B(n448), .Y(n1323) );
  AOI22X1 U620 ( .A(n481), .B(n227), .C(currentPlainKey[10]), .D(n219), .Y(
        n466) );
  INVX2 U621 ( .A(n450), .Y(n1422) );
  NAND2X1 U622 ( .A(n550), .B(n1422), .Y(n543) );
  NAND2X1 U623 ( .A(n471), .B(n543), .Y(n522) );
  INVX2 U624 ( .A(n522), .Y(n546) );
  OAI21X1 U625 ( .A(n25), .B(n172), .C(currentPlainKey[10]), .Y(n451) );
  OAI21X1 U626 ( .A(n1118), .B(n173), .C(n451), .Y(n453) );
  NOR2X1 U627 ( .A(n220), .B(n543), .Y(n452) );
  AOI21X1 U628 ( .A(n546), .B(n453), .C(n452), .Y(n455) );
  NAND2X1 U629 ( .A(n547), .B(n237), .Y(n454) );
  OAI21X1 U630 ( .A(n528), .B(n455), .C(n454), .Y(n456) );
  NAND2X1 U631 ( .A(n224), .B(n456), .Y(n459) );
  NAND2X1 U632 ( .A(n528), .B(n200), .Y(n458) );
  AOI21X1 U633 ( .A(n459), .B(n458), .C(n457), .Y(n460) );
  MUX2X1 U634 ( .B(n460), .A(n210), .S(n513), .Y(n462) );
  NAND2X1 U635 ( .A(n496), .B(n19), .Y(n461) );
  NAND2X1 U636 ( .A(n462), .B(n461), .Y(n464) );
  MUX2X1 U637 ( .B(n464), .A(n232), .S(n463), .Y(n465) );
  NAND2X1 U638 ( .A(n466), .B(n465), .Y(n1322) );
  NAND2X1 U639 ( .A(n528), .B(n209), .Y(n476) );
  OAI21X1 U640 ( .A(n164), .B(n172), .C(currentPlainKey[11]), .Y(n467) );
  OAI21X1 U641 ( .A(n1135), .B(n173), .C(n467), .Y(n468) );
  NAND3X1 U642 ( .A(n546), .B(n222), .C(n468), .Y(n469) );
  NAND2X1 U643 ( .A(n550), .B(n121), .Y(n504) );
  INVX2 U644 ( .A(n504), .Y(n581) );
  MUX2X1 U645 ( .B(n469), .A(n196), .S(n581), .Y(n473) );
  INVX2 U646 ( .A(n543), .Y(n563) );
  NAND2X1 U647 ( .A(n563), .B(n205), .Y(n470) );
  OAI21X1 U648 ( .A(n198), .B(n471), .C(n470), .Y(n472) );
  OAI21X1 U649 ( .A(n473), .B(n472), .C(n37), .Y(n475) );
  NAND2X1 U650 ( .A(n513), .B(n212), .Y(n474) );
  NAND3X1 U651 ( .A(n476), .B(n475), .C(n474), .Y(n479) );
  NOR2X1 U652 ( .A(n230), .B(n477), .Y(n478) );
  AOI21X1 U653 ( .A(n480), .B(n479), .C(n478), .Y(n483) );
  AOI22X1 U654 ( .A(n481), .B(n234), .C(currentPlainKey[11]), .D(n218), .Y(
        n482) );
  NAND2X1 U655 ( .A(n483), .B(n482), .Y(n1321) );
  AOI22X1 U656 ( .A(n513), .B(n227), .C(currentPlainKey[12]), .D(n218), .Y(
        n499) );
  NAND2X1 U657 ( .A(n550), .B(n127), .Y(n578) );
  OAI21X1 U658 ( .A(n63), .B(n172), .C(currentPlainKey[12]), .Y(n484) );
  OAI21X1 U659 ( .A(n1455), .B(n173), .C(n484), .Y(n486) );
  NOR2X1 U660 ( .A(n220), .B(n578), .Y(n485) );
  AOI21X1 U661 ( .A(n59), .B(n486), .C(n485), .Y(n488) );
  NAND2X1 U662 ( .A(n581), .B(n237), .Y(n487) );
  OAI21X1 U663 ( .A(n563), .B(n488), .C(n487), .Y(n489) );
  NAND2X1 U664 ( .A(n224), .B(n489), .Y(n492) );
  NAND2X1 U665 ( .A(n563), .B(n200), .Y(n491) );
  AOI21X1 U666 ( .A(n492), .B(n491), .C(n490), .Y(n493) );
  MUX2X1 U667 ( .B(n493), .A(n208), .S(n547), .Y(n495) );
  NAND2X1 U668 ( .A(n528), .B(n19), .Y(n494) );
  NAND2X1 U669 ( .A(n495), .B(n494), .Y(n497) );
  MUX2X1 U670 ( .B(n497), .A(n51), .S(n496), .Y(n498) );
  NAND2X1 U671 ( .A(n499), .B(n498), .Y(n1320) );
  NAND2X1 U672 ( .A(n563), .B(n103), .Y(n509) );
  OAI21X1 U673 ( .A(n168), .B(n172), .C(currentPlainKey[13]), .Y(n500) );
  OAI21X1 U674 ( .A(n1478), .B(n173), .C(n500), .Y(n501) );
  NAND3X1 U675 ( .A(n59), .B(n225), .C(n501), .Y(n502) );
  NAND2X1 U676 ( .A(n550), .B(n123), .Y(n537) );
  INVX2 U677 ( .A(n537), .Y(n613) );
  MUX2X1 U678 ( .B(n502), .A(n196), .S(n613), .Y(n506) );
  INVX2 U679 ( .A(n578), .Y(n596) );
  NAND2X1 U680 ( .A(n596), .B(n205), .Y(n503) );
  OAI21X1 U681 ( .A(n198), .B(n504), .C(n503), .Y(n505) );
  OAI21X1 U682 ( .A(n506), .B(n505), .C(n546), .Y(n508) );
  NAND2X1 U683 ( .A(n547), .B(n214), .Y(n507) );
  NAND3X1 U684 ( .A(n509), .B(n508), .C(n507), .Y(n512) );
  NOR2X1 U685 ( .A(n229), .B(n510), .Y(n511) );
  AOI21X1 U686 ( .A(n37), .B(n512), .C(n511), .Y(n515) );
  AOI22X1 U687 ( .A(n513), .B(n233), .C(currentPlainKey[13]), .D(n218), .Y(
        n514) );
  NAND2X1 U688 ( .A(n515), .B(n514), .Y(n1319) );
  AOI22X1 U689 ( .A(n547), .B(n227), .C(currentPlainKey[14]), .D(n218), .Y(
        n531) );
  NAND2X1 U690 ( .A(n550), .B(n125), .Y(n610) );
  OAI21X1 U691 ( .A(n1185), .B(n172), .C(currentPlainKey[14]), .Y(n516) );
  OAI21X1 U692 ( .A(n1490), .B(n173), .C(n516), .Y(n518) );
  NOR2X1 U693 ( .A(n220), .B(n610), .Y(n517) );
  AOI21X1 U694 ( .A(n77), .B(n518), .C(n517), .Y(n520) );
  NAND2X1 U695 ( .A(n613), .B(n237), .Y(n519) );
  OAI21X1 U696 ( .A(n596), .B(n520), .C(n519), .Y(n521) );
  NAND2X1 U697 ( .A(n225), .B(n521), .Y(n524) );
  NAND2X1 U698 ( .A(n596), .B(n201), .Y(n523) );
  AOI21X1 U699 ( .A(n524), .B(n523), .C(n522), .Y(n525) );
  MUX2X1 U700 ( .B(n525), .A(n208), .S(n581), .Y(n527) );
  NAND2X1 U701 ( .A(n563), .B(n214), .Y(n526) );
  NAND2X1 U702 ( .A(n527), .B(n526), .Y(n529) );
  MUX2X1 U703 ( .B(n529), .A(n234), .S(n528), .Y(n530) );
  NAND2X1 U704 ( .A(n531), .B(n530), .Y(n1318) );
  NAND2X1 U705 ( .A(n596), .B(n209), .Y(n542) );
  OAI21X1 U706 ( .A(n166), .B(n172), .C(currentPlainKey[15]), .Y(n532) );
  OAI21X1 U707 ( .A(n1361), .B(n173), .C(n532), .Y(n534) );
  NAND3X1 U708 ( .A(n77), .B(n225), .C(n534), .Y(n535) );
  NAND2X1 U709 ( .A(n550), .B(n93), .Y(n572) );
  INVX2 U710 ( .A(n572), .Y(n645) );
  MUX2X1 U711 ( .B(n535), .A(n195), .S(n645), .Y(n539) );
  INVX2 U712 ( .A(n610), .Y(n628) );
  NAND2X1 U713 ( .A(n628), .B(n205), .Y(n536) );
  OAI21X1 U714 ( .A(n198), .B(n537), .C(n536), .Y(n538) );
  OAI21X1 U715 ( .A(n539), .B(n538), .C(n59), .Y(n541) );
  NAND2X1 U716 ( .A(n581), .B(n19), .Y(n540) );
  NAND3X1 U717 ( .A(n542), .B(n541), .C(n540), .Y(n545) );
  NOR2X1 U718 ( .A(n229), .B(n543), .Y(n544) );
  AOI21X1 U719 ( .A(n546), .B(n545), .C(n544), .Y(n549) );
  AOI22X1 U720 ( .A(n547), .B(n231), .C(currentPlainKey[15]), .D(n218), .Y(
        n548) );
  NAND2X1 U721 ( .A(n549), .B(n548), .Y(n1317) );
  AOI22X1 U722 ( .A(n581), .B(n227), .C(currentPlainKey[16]), .D(n218), .Y(
        n566) );
  NAND2X1 U723 ( .A(n550), .B(n133), .Y(n642) );
  NAND3X1 U724 ( .A(address[4]), .B(n1101), .C(n682), .Y(n665) );
  OAI21X1 U725 ( .A(n1081), .B(n175), .C(currentPlainKey[16]), .Y(n551) );
  OAI21X1 U726 ( .A(n1083), .B(n176), .C(n551), .Y(n553) );
  NOR2X1 U727 ( .A(n220), .B(n642), .Y(n552) );
  AOI21X1 U728 ( .A(n99), .B(n553), .C(n552), .Y(n555) );
  NAND2X1 U729 ( .A(n645), .B(n237), .Y(n554) );
  OAI21X1 U730 ( .A(n628), .B(n555), .C(n554), .Y(n556) );
  NAND2X1 U731 ( .A(n225), .B(n556), .Y(n559) );
  NAND2X1 U732 ( .A(n628), .B(n204), .Y(n558) );
  AOI21X1 U733 ( .A(n559), .B(n558), .C(n557), .Y(n560) );
  MUX2X1 U734 ( .B(n560), .A(n105), .S(n613), .Y(n562) );
  NAND2X1 U735 ( .A(n596), .B(n213), .Y(n561) );
  NAND2X1 U736 ( .A(n562), .B(n561), .Y(n564) );
  MUX2X1 U737 ( .B(n564), .A(n232), .S(n563), .Y(n565) );
  NAND2X1 U738 ( .A(n566), .B(n565), .Y(n1316) );
  NAND2X1 U739 ( .A(n628), .B(n105), .Y(n577) );
  OAI21X1 U740 ( .A(n170), .B(n175), .C(currentPlainKey[17]), .Y(n567) );
  OAI21X1 U741 ( .A(n1402), .B(n176), .C(n567), .Y(n568) );
  NAND3X1 U742 ( .A(n99), .B(n222), .C(n568), .Y(n570) );
  NAND3X1 U743 ( .A(n155), .B(address[4]), .C(n682), .Y(n569) );
  NAND2X1 U744 ( .A(n145), .B(n43), .Y(n604) );
  INVX2 U745 ( .A(n604), .Y(n679) );
  MUX2X1 U746 ( .B(n570), .A(n196), .S(n679), .Y(n574) );
  INVX2 U747 ( .A(n642), .Y(n660) );
  NAND2X1 U748 ( .A(n660), .B(n205), .Y(n571) );
  OAI21X1 U749 ( .A(n198), .B(n572), .C(n571), .Y(n573) );
  OAI21X1 U750 ( .A(n574), .B(n573), .C(n77), .Y(n576) );
  NAND2X1 U751 ( .A(n613), .B(n20), .Y(n575) );
  NAND3X1 U752 ( .A(n577), .B(n576), .C(n575), .Y(n580) );
  NOR2X1 U753 ( .A(n229), .B(n578), .Y(n579) );
  AOI21X1 U754 ( .A(n59), .B(n580), .C(n579), .Y(n583) );
  AOI22X1 U755 ( .A(n581), .B(n231), .C(currentPlainKey[17]), .D(n218), .Y(
        n582) );
  NAND2X1 U756 ( .A(n583), .B(n582), .Y(n1315) );
  AOI22X1 U757 ( .A(n613), .B(n227), .C(currentPlainKey[18]), .D(n218), .Y(
        n599) );
  NAND2X1 U758 ( .A(n145), .B(n169), .Y(n675) );
  NAND2X1 U759 ( .A(n604), .B(n675), .Y(n654) );
  INVX2 U760 ( .A(n654), .Y(n678) );
  OAI21X1 U761 ( .A(n25), .B(n175), .C(currentPlainKey[18]), .Y(n584) );
  OAI21X1 U762 ( .A(n1118), .B(n176), .C(n584), .Y(n586) );
  NOR2X1 U763 ( .A(n220), .B(n675), .Y(n585) );
  AOI21X1 U764 ( .A(n678), .B(n586), .C(n585), .Y(n588) );
  NAND2X1 U765 ( .A(n679), .B(n237), .Y(n587) );
  OAI21X1 U766 ( .A(n660), .B(n588), .C(n587), .Y(n589) );
  NAND2X1 U767 ( .A(n224), .B(n589), .Y(n592) );
  NAND2X1 U768 ( .A(n660), .B(n204), .Y(n591) );
  AOI21X1 U769 ( .A(n592), .B(n591), .C(n590), .Y(n593) );
  MUX2X1 U770 ( .B(n593), .A(n209), .S(n645), .Y(n595) );
  NAND2X1 U771 ( .A(n628), .B(n213), .Y(n594) );
  NAND2X1 U772 ( .A(n595), .B(n594), .Y(n597) );
  MUX2X1 U773 ( .B(n597), .A(n51), .S(n596), .Y(n598) );
  NAND2X1 U774 ( .A(n599), .B(n598), .Y(n1314) );
  NAND2X1 U775 ( .A(n660), .B(n103), .Y(n609) );
  OAI21X1 U776 ( .A(n164), .B(n175), .C(currentPlainKey[19]), .Y(n600) );
  OAI21X1 U777 ( .A(n1135), .B(n176), .C(n600), .Y(n601) );
  NAND3X1 U778 ( .A(n678), .B(n224), .C(n601), .Y(n602) );
  NAND2X1 U779 ( .A(n145), .B(n1420), .Y(n636) );
  INVX2 U780 ( .A(n636), .Y(n713) );
  MUX2X1 U781 ( .B(n602), .A(n195), .S(n713), .Y(n606) );
  INVX2 U782 ( .A(n675), .Y(n695) );
  NAND2X1 U783 ( .A(n695), .B(n205), .Y(n603) );
  OAI21X1 U784 ( .A(n198), .B(n604), .C(n603), .Y(n605) );
  OAI21X1 U785 ( .A(n606), .B(n605), .C(n99), .Y(n608) );
  NAND2X1 U786 ( .A(n645), .B(n213), .Y(n607) );
  NAND3X1 U787 ( .A(n609), .B(n608), .C(n607), .Y(n612) );
  NOR2X1 U788 ( .A(n230), .B(n6), .Y(n611) );
  AOI21X1 U789 ( .A(n77), .B(n612), .C(n611), .Y(n615) );
  AOI22X1 U790 ( .A(n613), .B(n235), .C(currentPlainKey[19]), .D(n218), .Y(
        n614) );
  NAND2X1 U791 ( .A(n615), .B(n614), .Y(n1313) );
  AOI22X1 U792 ( .A(n645), .B(n227), .C(currentPlainKey[20]), .D(n218), .Y(
        n631) );
  NAND2X1 U793 ( .A(n145), .B(n163), .Y(n709) );
  NAND2X1 U794 ( .A(n636), .B(n709), .Y(n689) );
  INVX2 U795 ( .A(n689), .Y(n712) );
  OAI21X1 U796 ( .A(n63), .B(n175), .C(currentPlainKey[20]), .Y(n616) );
  OAI21X1 U797 ( .A(n1455), .B(n176), .C(n616), .Y(n618) );
  NOR2X1 U798 ( .A(n220), .B(n709), .Y(n617) );
  AOI21X1 U799 ( .A(n712), .B(n618), .C(n617), .Y(n620) );
  NAND2X1 U800 ( .A(n713), .B(n236), .Y(n619) );
  OAI21X1 U801 ( .A(n695), .B(n620), .C(n619), .Y(n621) );
  NAND2X1 U802 ( .A(n224), .B(n621), .Y(n624) );
  NAND2X1 U803 ( .A(n695), .B(n201), .Y(n623) );
  AOI21X1 U804 ( .A(n624), .B(n623), .C(n622), .Y(n625) );
  MUX2X1 U805 ( .B(n625), .A(n103), .S(n679), .Y(n627) );
  NAND2X1 U806 ( .A(n660), .B(n19), .Y(n626) );
  NAND2X1 U807 ( .A(n627), .B(n626), .Y(n629) );
  MUX2X1 U808 ( .B(n629), .A(n234), .S(n628), .Y(n630) );
  NAND2X1 U809 ( .A(n631), .B(n630), .Y(n1312) );
  NAND2X1 U810 ( .A(n695), .B(n208), .Y(n641) );
  OAI21X1 U811 ( .A(n168), .B(n175), .C(currentPlainKey[21]), .Y(n632) );
  OAI21X1 U812 ( .A(n1478), .B(n176), .C(n632), .Y(n633) );
  NAND3X1 U813 ( .A(n712), .B(n225), .C(n633), .Y(n634) );
  NAND2X1 U814 ( .A(n145), .B(n61), .Y(n669) );
  INVX2 U815 ( .A(n669), .Y(n746) );
  MUX2X1 U816 ( .B(n634), .A(n195), .S(n746), .Y(n638) );
  INVX2 U817 ( .A(n709), .Y(n728) );
  NAND2X1 U818 ( .A(n728), .B(n205), .Y(n635) );
  OAI21X1 U819 ( .A(n198), .B(n636), .C(n635), .Y(n637) );
  OAI21X1 U820 ( .A(n638), .B(n637), .C(n678), .Y(n640) );
  NAND2X1 U821 ( .A(n679), .B(n212), .Y(n639) );
  NAND3X1 U822 ( .A(n641), .B(n640), .C(n639), .Y(n644) );
  NOR2X1 U823 ( .A(n229), .B(n642), .Y(n643) );
  AOI21X1 U824 ( .A(n99), .B(n644), .C(n643), .Y(n647) );
  AOI22X1 U825 ( .A(n645), .B(n234), .C(currentPlainKey[21]), .D(n218), .Y(
        n646) );
  NAND2X1 U826 ( .A(n647), .B(n646), .Y(n1311) );
  AOI22X1 U827 ( .A(n679), .B(n227), .C(currentPlainKey[22]), .D(n218), .Y(
        n663) );
  NAND2X1 U828 ( .A(n145), .B(n167), .Y(n742) );
  NAND2X1 U829 ( .A(n669), .B(n742), .Y(n722) );
  INVX2 U830 ( .A(n722), .Y(n745) );
  OAI21X1 U831 ( .A(n1185), .B(n175), .C(currentPlainKey[22]), .Y(n648) );
  OAI21X1 U832 ( .A(n1490), .B(n176), .C(n648), .Y(n650) );
  NOR2X1 U833 ( .A(n221), .B(n742), .Y(n649) );
  AOI21X1 U834 ( .A(n745), .B(n650), .C(n649), .Y(n652) );
  NAND2X1 U835 ( .A(n746), .B(n236), .Y(n651) );
  OAI21X1 U836 ( .A(n728), .B(n652), .C(n651), .Y(n653) );
  NAND2X1 U837 ( .A(n224), .B(n653), .Y(n656) );
  NAND2X1 U838 ( .A(n728), .B(n200), .Y(n655) );
  AOI21X1 U839 ( .A(n656), .B(n655), .C(n654), .Y(n657) );
  MUX2X1 U840 ( .B(n657), .A(n103), .S(n713), .Y(n659) );
  NAND2X1 U841 ( .A(n695), .B(n19), .Y(n658) );
  NAND2X1 U842 ( .A(n659), .B(n658), .Y(n661) );
  MUX2X1 U843 ( .B(n661), .A(n233), .S(n660), .Y(n662) );
  NAND2X1 U844 ( .A(n663), .B(n662), .Y(n1310) );
  NAND2X1 U845 ( .A(n728), .B(n208), .Y(n674) );
  OAI21X1 U846 ( .A(n166), .B(n175), .C(currentPlainKey[23]), .Y(n664) );
  OAI21X1 U847 ( .A(n1361), .B(n176), .C(n664), .Y(n666) );
  NAND3X1 U848 ( .A(n745), .B(n225), .C(n666), .Y(n667) );
  NAND2X1 U849 ( .A(n145), .B(n89), .Y(n703) );
  INVX2 U850 ( .A(n703), .Y(n779) );
  MUX2X1 U851 ( .B(n667), .A(n195), .S(n779), .Y(n671) );
  INVX2 U852 ( .A(n742), .Y(n761) );
  NAND2X1 U853 ( .A(n761), .B(n205), .Y(n668) );
  OAI21X1 U854 ( .A(n198), .B(n669), .C(n668), .Y(n670) );
  OAI21X1 U855 ( .A(n671), .B(n670), .C(n712), .Y(n673) );
  NAND2X1 U856 ( .A(n713), .B(n213), .Y(n672) );
  NAND3X1 U857 ( .A(n674), .B(n673), .C(n672), .Y(n677) );
  NOR2X1 U858 ( .A(n229), .B(n675), .Y(n676) );
  AOI21X1 U859 ( .A(n678), .B(n677), .C(n676), .Y(n681) );
  AOI22X1 U860 ( .A(n679), .B(n233), .C(currentPlainKey[23]), .D(n217), .Y(
        n680) );
  NAND2X1 U861 ( .A(n681), .B(n680), .Y(n1309) );
  AOI22X1 U862 ( .A(n713), .B(n227), .C(currentPlainKey[24]), .D(n217), .Y(
        n698) );
  NAND2X1 U863 ( .A(n145), .B(n152), .Y(n775) );
  NAND2X1 U864 ( .A(n703), .B(n775), .Y(n755) );
  INVX2 U865 ( .A(n755), .Y(n778) );
  NAND3X1 U866 ( .A(n192), .B(address[4]), .C(n682), .Y(n799) );
  OAI21X1 U867 ( .A(n1081), .B(n178), .C(currentPlainKey[24]), .Y(n683) );
  OAI21X1 U868 ( .A(n1083), .B(n179), .C(n683), .Y(n685) );
  NOR2X1 U869 ( .A(n221), .B(n775), .Y(n684) );
  AOI21X1 U870 ( .A(n778), .B(n685), .C(n684), .Y(n687) );
  NAND2X1 U871 ( .A(n779), .B(n236), .Y(n686) );
  OAI21X1 U872 ( .A(n761), .B(n687), .C(n686), .Y(n688) );
  NAND2X1 U873 ( .A(n225), .B(n688), .Y(n691) );
  NAND2X1 U874 ( .A(n761), .B(n203), .Y(n690) );
  AOI21X1 U875 ( .A(n691), .B(n690), .C(n689), .Y(n692) );
  MUX2X1 U876 ( .B(n692), .A(n105), .S(n746), .Y(n694) );
  NAND2X1 U877 ( .A(n728), .B(n214), .Y(n693) );
  NAND2X1 U878 ( .A(n694), .B(n693), .Y(n696) );
  MUX2X1 U879 ( .B(n696), .A(n51), .S(n695), .Y(n697) );
  NAND2X1 U880 ( .A(n698), .B(n697), .Y(n1308) );
  NAND2X1 U881 ( .A(n761), .B(n208), .Y(n708) );
  OAI21X1 U882 ( .A(n170), .B(n178), .C(currentPlainKey[25]), .Y(n699) );
  OAI21X1 U883 ( .A(n1402), .B(n179), .C(n699), .Y(n700) );
  NAND3X1 U884 ( .A(n778), .B(n222), .C(n700), .Y(n701) );
  NAND2X1 U885 ( .A(n816), .B(n131), .Y(n736) );
  INVX2 U886 ( .A(n736), .Y(n813) );
  MUX2X1 U887 ( .B(n701), .A(n195), .S(n813), .Y(n705) );
  INVX2 U888 ( .A(n775), .Y(n794) );
  NAND2X1 U889 ( .A(n794), .B(n205), .Y(n702) );
  OAI21X1 U890 ( .A(n198), .B(n703), .C(n702), .Y(n704) );
  OAI21X1 U891 ( .A(n705), .B(n704), .C(n745), .Y(n707) );
  NAND2X1 U892 ( .A(n746), .B(n213), .Y(n706) );
  NAND3X1 U893 ( .A(n708), .B(n707), .C(n706), .Y(n711) );
  NOR2X1 U894 ( .A(n229), .B(n709), .Y(n710) );
  AOI21X1 U895 ( .A(n712), .B(n711), .C(n710), .Y(n715) );
  AOI22X1 U896 ( .A(n713), .B(n235), .C(currentPlainKey[25]), .D(n217), .Y(
        n714) );
  NAND2X1 U897 ( .A(n715), .B(n714), .Y(n1307) );
  AOI22X1 U898 ( .A(n746), .B(n227), .C(currentPlainKey[26]), .D(n217), .Y(
        n731) );
  NAND2X1 U899 ( .A(n816), .B(n1422), .Y(n809) );
  NAND2X1 U900 ( .A(n736), .B(n809), .Y(n788) );
  INVX2 U901 ( .A(n788), .Y(n812) );
  OAI21X1 U902 ( .A(n25), .B(n178), .C(currentPlainKey[26]), .Y(n716) );
  OAI21X1 U903 ( .A(n1118), .B(n179), .C(n716), .Y(n718) );
  NOR2X1 U904 ( .A(n221), .B(n809), .Y(n717) );
  AOI21X1 U905 ( .A(n812), .B(n718), .C(n717), .Y(n720) );
  NAND2X1 U906 ( .A(n813), .B(n236), .Y(n719) );
  OAI21X1 U907 ( .A(n794), .B(n720), .C(n719), .Y(n721) );
  NAND2X1 U908 ( .A(n225), .B(n721), .Y(n724) );
  NAND2X1 U909 ( .A(n794), .B(n204), .Y(n723) );
  AOI21X1 U910 ( .A(n724), .B(n723), .C(n722), .Y(n725) );
  MUX2X1 U911 ( .B(n725), .A(n105), .S(n779), .Y(n727) );
  NAND2X1 U912 ( .A(n761), .B(n213), .Y(n726) );
  NAND2X1 U913 ( .A(n727), .B(n726), .Y(n729) );
  MUX2X1 U914 ( .B(n729), .A(n232), .S(n728), .Y(n730) );
  NAND2X1 U915 ( .A(n731), .B(n730), .Y(n1306) );
  NAND2X1 U916 ( .A(n794), .B(n208), .Y(n741) );
  OAI21X1 U917 ( .A(n164), .B(n178), .C(currentPlainKey[27]), .Y(n732) );
  OAI21X1 U918 ( .A(n1135), .B(n179), .C(n732), .Y(n733) );
  NAND3X1 U919 ( .A(n812), .B(n222), .C(n733), .Y(n734) );
  NAND2X1 U920 ( .A(n816), .B(n121), .Y(n769) );
  INVX2 U921 ( .A(n769), .Y(n847) );
  MUX2X1 U922 ( .B(n734), .A(n195), .S(n847), .Y(n738) );
  INVX2 U923 ( .A(n809), .Y(n829) );
  NAND2X1 U924 ( .A(n829), .B(n205), .Y(n735) );
  OAI21X1 U925 ( .A(n198), .B(n736), .C(n735), .Y(n737) );
  OAI21X1 U926 ( .A(n738), .B(n737), .C(n778), .Y(n740) );
  NAND2X1 U927 ( .A(n779), .B(n212), .Y(n739) );
  NAND3X1 U928 ( .A(n741), .B(n740), .C(n739), .Y(n744) );
  NOR2X1 U929 ( .A(n229), .B(n742), .Y(n743) );
  AOI21X1 U930 ( .A(n745), .B(n744), .C(n743), .Y(n748) );
  AOI22X1 U931 ( .A(n746), .B(n232), .C(currentPlainKey[27]), .D(n217), .Y(
        n747) );
  NAND2X1 U932 ( .A(n748), .B(n747), .Y(n1305) );
  AOI22X1 U933 ( .A(n779), .B(n227), .C(currentPlainKey[28]), .D(n217), .Y(
        n764) );
  NAND2X1 U934 ( .A(n816), .B(n127), .Y(n844) );
  OAI21X1 U935 ( .A(n63), .B(n178), .C(currentPlainKey[28]), .Y(n749) );
  OAI21X1 U936 ( .A(n1455), .B(n179), .C(n749), .Y(n751) );
  NOR2X1 U937 ( .A(n221), .B(n844), .Y(n750) );
  AOI21X1 U938 ( .A(n49), .B(n751), .C(n750), .Y(n753) );
  NAND2X1 U939 ( .A(n847), .B(n236), .Y(n752) );
  OAI21X1 U940 ( .A(n829), .B(n753), .C(n752), .Y(n754) );
  NAND2X1 U941 ( .A(n224), .B(n754), .Y(n757) );
  NAND2X1 U942 ( .A(n829), .B(n201), .Y(n756) );
  AOI21X1 U943 ( .A(n757), .B(n756), .C(n755), .Y(n758) );
  MUX2X1 U944 ( .B(n758), .A(n103), .S(n813), .Y(n760) );
  NAND2X1 U945 ( .A(n794), .B(n20), .Y(n759) );
  NAND2X1 U946 ( .A(n760), .B(n759), .Y(n762) );
  MUX2X1 U947 ( .B(n762), .A(n234), .S(n761), .Y(n763) );
  NAND2X1 U948 ( .A(n764), .B(n763), .Y(n1304) );
  NAND2X1 U949 ( .A(n829), .B(n208), .Y(n774) );
  OAI21X1 U950 ( .A(n168), .B(n178), .C(currentPlainKey[29]), .Y(n765) );
  OAI21X1 U951 ( .A(n1478), .B(n179), .C(n765), .Y(n766) );
  NAND3X1 U952 ( .A(n49), .B(n224), .C(n766), .Y(n767) );
  NAND2X1 U953 ( .A(n816), .B(n123), .Y(n803) );
  INVX2 U954 ( .A(n803), .Y(n879) );
  MUX2X1 U955 ( .B(n767), .A(n196), .S(n879), .Y(n771) );
  INVX2 U956 ( .A(n844), .Y(n862) );
  NAND2X1 U957 ( .A(n862), .B(n206), .Y(n768) );
  OAI21X1 U958 ( .A(n198), .B(n769), .C(n768), .Y(n770) );
  OAI21X1 U959 ( .A(n771), .B(n770), .C(n812), .Y(n773) );
  NAND2X1 U960 ( .A(n813), .B(n19), .Y(n772) );
  NAND3X1 U961 ( .A(n774), .B(n773), .C(n772), .Y(n777) );
  NOR2X1 U962 ( .A(n230), .B(n775), .Y(n776) );
  AOI21X1 U963 ( .A(n778), .B(n777), .C(n776), .Y(n781) );
  AOI22X1 U964 ( .A(n779), .B(n234), .C(currentPlainKey[29]), .D(n217), .Y(
        n780) );
  NAND2X1 U965 ( .A(n781), .B(n780), .Y(n1303) );
  AOI22X1 U966 ( .A(n813), .B(n227), .C(currentPlainKey[30]), .D(n217), .Y(
        n797) );
  NAND2X1 U967 ( .A(n816), .B(n125), .Y(n876) );
  OAI21X1 U968 ( .A(n1185), .B(n178), .C(currentPlainKey[30]), .Y(n782) );
  OAI21X1 U969 ( .A(n1490), .B(n179), .C(n782), .Y(n784) );
  NOR2X1 U970 ( .A(n221), .B(n876), .Y(n783) );
  AOI21X1 U971 ( .A(n75), .B(n784), .C(n783), .Y(n786) );
  NAND2X1 U972 ( .A(n879), .B(n236), .Y(n785) );
  OAI21X1 U973 ( .A(n862), .B(n786), .C(n785), .Y(n787) );
  NAND2X1 U974 ( .A(n224), .B(n787), .Y(n790) );
  NAND2X1 U975 ( .A(n862), .B(n200), .Y(n789) );
  AOI21X1 U976 ( .A(n790), .B(n789), .C(n788), .Y(n791) );
  MUX2X1 U977 ( .B(n791), .A(n208), .S(n847), .Y(n793) );
  NAND2X1 U978 ( .A(n829), .B(n212), .Y(n792) );
  NAND2X1 U979 ( .A(n793), .B(n792), .Y(n795) );
  MUX2X1 U980 ( .B(n795), .A(n232), .S(n794), .Y(n796) );
  NAND2X1 U981 ( .A(n797), .B(n796), .Y(n1302) );
  NAND2X1 U982 ( .A(n862), .B(n210), .Y(n808) );
  OAI21X1 U983 ( .A(n166), .B(n178), .C(currentPlainKey[31]), .Y(n798) );
  OAI21X1 U984 ( .A(n1361), .B(n179), .C(n798), .Y(n800) );
  NAND3X1 U985 ( .A(n75), .B(n222), .C(n800), .Y(n801) );
  NAND2X1 U986 ( .A(n816), .B(n93), .Y(n838) );
  INVX2 U987 ( .A(n838), .Y(n911) );
  MUX2X1 U988 ( .B(n801), .A(n196), .S(n911), .Y(n805) );
  INVX2 U989 ( .A(n876), .Y(n894) );
  NAND2X1 U990 ( .A(n894), .B(n206), .Y(n802) );
  OAI21X1 U991 ( .A(n197), .B(n803), .C(n802), .Y(n804) );
  OAI21X1 U992 ( .A(n805), .B(n804), .C(n49), .Y(n807) );
  NAND2X1 U993 ( .A(n847), .B(n212), .Y(n806) );
  NAND3X1 U994 ( .A(n808), .B(n807), .C(n806), .Y(n811) );
  NOR2X1 U995 ( .A(n229), .B(n809), .Y(n810) );
  AOI21X1 U996 ( .A(n812), .B(n811), .C(n810), .Y(n815) );
  AOI22X1 U997 ( .A(n813), .B(n232), .C(currentPlainKey[31]), .D(n217), .Y(
        n814) );
  NAND2X1 U998 ( .A(n815), .B(n814), .Y(n1301) );
  AOI22X1 U999 ( .A(n847), .B(n227), .C(currentPlainKey[32]), .D(n217), .Y(
        n832) );
  NAND2X1 U1000 ( .A(n816), .B(n133), .Y(n908) );
  NAND3X1 U1001 ( .A(address[5]), .B(n1101), .C(n948), .Y(n931) );
  OAI21X1 U1002 ( .A(n1081), .B(n181), .C(currentPlainKey[32]), .Y(n817) );
  OAI21X1 U1003 ( .A(n1083), .B(n182), .C(n817), .Y(n819) );
  NOR2X1 U1004 ( .A(n221), .B(n908), .Y(n818) );
  AOI21X1 U1005 ( .A(n91), .B(n819), .C(n818), .Y(n821) );
  NAND2X1 U1006 ( .A(n911), .B(n236), .Y(n820) );
  OAI21X1 U1007 ( .A(n821), .B(n894), .C(n820), .Y(n822) );
  NAND2X1 U1008 ( .A(n225), .B(n822), .Y(n825) );
  NAND2X1 U1009 ( .A(n894), .B(n203), .Y(n824) );
  AOI21X1 U1010 ( .A(n825), .B(n824), .C(n823), .Y(n826) );
  MUX2X1 U1011 ( .B(n826), .A(n103), .S(n879), .Y(n828) );
  NAND2X1 U1012 ( .A(n862), .B(n213), .Y(n827) );
  NAND2X1 U1013 ( .A(n828), .B(n827), .Y(n830) );
  MUX2X1 U1014 ( .B(n830), .A(n234), .S(n829), .Y(n831) );
  NAND2X1 U1015 ( .A(n832), .B(n831), .Y(n1300) );
  NAND2X1 U1016 ( .A(n894), .B(n105), .Y(n843) );
  OAI21X1 U1017 ( .A(n170), .B(n181), .C(currentPlainKey[33]), .Y(n833) );
  OAI21X1 U1018 ( .A(n1402), .B(n182), .C(n833), .Y(n834) );
  NAND3X1 U1019 ( .A(n91), .B(n224), .C(n834), .Y(n836) );
  NAND3X1 U1020 ( .A(n29), .B(address[5]), .C(n948), .Y(n835) );
  NAND2X1 U1021 ( .A(n143), .B(n43), .Y(n870) );
  INVX2 U1022 ( .A(n870), .Y(n945) );
  MUX2X1 U1023 ( .B(n836), .A(n196), .S(n945), .Y(n840) );
  INVX2 U1024 ( .A(n908), .Y(n926) );
  NAND2X1 U1025 ( .A(n926), .B(n206), .Y(n837) );
  OAI21X1 U1026 ( .A(n197), .B(n95), .C(n837), .Y(n839) );
  OAI21X1 U1027 ( .A(n840), .B(n839), .C(n75), .Y(n842) );
  NAND2X1 U1028 ( .A(n879), .B(n213), .Y(n841) );
  NAND3X1 U1029 ( .A(n843), .B(n842), .C(n841), .Y(n846) );
  NOR2X1 U1030 ( .A(n230), .B(n844), .Y(n845) );
  AOI21X1 U1031 ( .A(n49), .B(n846), .C(n845), .Y(n849) );
  AOI22X1 U1032 ( .A(n847), .B(n233), .C(currentPlainKey[33]), .D(n217), .Y(
        n848) );
  NAND2X1 U1033 ( .A(n849), .B(n848), .Y(n1299) );
  AOI22X1 U1034 ( .A(n879), .B(n226), .C(currentPlainKey[34]), .D(n217), .Y(
        n865) );
  NAND2X1 U1035 ( .A(n143), .B(n169), .Y(n941) );
  NAND2X1 U1036 ( .A(n870), .B(n941), .Y(n920) );
  INVX2 U1037 ( .A(n920), .Y(n944) );
  OAI21X1 U1038 ( .A(n25), .B(n181), .C(currentPlainKey[34]), .Y(n850) );
  OAI21X1 U1039 ( .A(n1118), .B(n182), .C(n850), .Y(n852) );
  NOR2X1 U1040 ( .A(n221), .B(n941), .Y(n851) );
  AOI21X1 U1041 ( .A(n944), .B(n852), .C(n851), .Y(n854) );
  NAND2X1 U1042 ( .A(n945), .B(n236), .Y(n853) );
  OAI21X1 U1043 ( .A(n926), .B(n854), .C(n853), .Y(n855) );
  NAND2X1 U1044 ( .A(n222), .B(n855), .Y(n858) );
  NAND2X1 U1045 ( .A(n926), .B(n203), .Y(n857) );
  AOI21X1 U1046 ( .A(n858), .B(n857), .C(n856), .Y(n859) );
  MUX2X1 U1047 ( .B(n859), .A(n105), .S(n911), .Y(n861) );
  NAND2X1 U1048 ( .A(n894), .B(n212), .Y(n860) );
  NAND2X1 U1049 ( .A(n861), .B(n860), .Y(n863) );
  MUX2X1 U1050 ( .B(n863), .A(n233), .S(n862), .Y(n864) );
  NAND2X1 U1051 ( .A(n865), .B(n864), .Y(n1298) );
  NAND2X1 U1052 ( .A(n926), .B(n105), .Y(n875) );
  OAI21X1 U1053 ( .A(n164), .B(n181), .C(currentPlainKey[35]), .Y(n866) );
  OAI21X1 U1054 ( .A(n1135), .B(n182), .C(n866), .Y(n867) );
  NAND3X1 U1055 ( .A(n944), .B(n224), .C(n867), .Y(n868) );
  NAND2X1 U1056 ( .A(n143), .B(n1420), .Y(n902) );
  INVX2 U1057 ( .A(n902), .Y(n978) );
  MUX2X1 U1058 ( .B(n868), .A(n195), .S(n978), .Y(n872) );
  INVX2 U1059 ( .A(n941), .Y(n961) );
  NAND2X1 U1060 ( .A(n961), .B(n206), .Y(n869) );
  OAI21X1 U1061 ( .A(n197), .B(n870), .C(n869), .Y(n871) );
  OAI21X1 U1062 ( .A(n872), .B(n871), .C(n91), .Y(n874) );
  NAND2X1 U1063 ( .A(n911), .B(n20), .Y(n873) );
  NAND3X1 U1064 ( .A(n875), .B(n874), .C(n873), .Y(n878) );
  NOR2X1 U1065 ( .A(n230), .B(n5), .Y(n877) );
  AOI21X1 U1066 ( .A(n75), .B(n878), .C(n877), .Y(n881) );
  AOI22X1 U1067 ( .A(n879), .B(n233), .C(currentPlainKey[35]), .D(n216), .Y(
        n880) );
  NAND2X1 U1068 ( .A(n881), .B(n880), .Y(n1297) );
  AOI22X1 U1069 ( .A(n911), .B(n226), .C(currentPlainKey[36]), .D(n216), .Y(
        n897) );
  NAND2X1 U1070 ( .A(n143), .B(n163), .Y(n975) );
  OAI21X1 U1071 ( .A(n63), .B(n181), .C(currentPlainKey[36]), .Y(n882) );
  OAI21X1 U1072 ( .A(n1455), .B(n182), .C(n882), .Y(n884) );
  NOR2X1 U1073 ( .A(n221), .B(n975), .Y(n883) );
  AOI21X1 U1074 ( .A(n35), .B(n884), .C(n883), .Y(n886) );
  NAND2X1 U1075 ( .A(n978), .B(n236), .Y(n885) );
  OAI21X1 U1076 ( .A(n961), .B(n886), .C(n885), .Y(n887) );
  NAND2X1 U1077 ( .A(n224), .B(n887), .Y(n890) );
  NAND2X1 U1078 ( .A(n961), .B(n200), .Y(n889) );
  AOI21X1 U1079 ( .A(n890), .B(n889), .C(n888), .Y(n891) );
  MUX2X1 U1080 ( .B(n891), .A(n208), .S(n945), .Y(n893) );
  NAND2X1 U1081 ( .A(n926), .B(n213), .Y(n892) );
  NAND2X1 U1082 ( .A(n893), .B(n892), .Y(n895) );
  MUX2X1 U1083 ( .B(n895), .A(n234), .S(n894), .Y(n896) );
  NAND2X1 U1084 ( .A(n897), .B(n896), .Y(n1296) );
  NAND2X1 U1085 ( .A(n961), .B(n162), .Y(n907) );
  OAI21X1 U1086 ( .A(n168), .B(n181), .C(currentPlainKey[37]), .Y(n898) );
  OAI21X1 U1087 ( .A(n1478), .B(n182), .C(n898), .Y(n899) );
  NAND3X1 U1088 ( .A(n35), .B(n222), .C(n899), .Y(n900) );
  NAND2X1 U1089 ( .A(n143), .B(n61), .Y(n935) );
  INVX2 U1090 ( .A(n935), .Y(n1010) );
  MUX2X1 U1091 ( .B(n900), .A(n195), .S(n1010), .Y(n904) );
  INVX2 U1092 ( .A(n975), .Y(n993) );
  NAND2X1 U1093 ( .A(n993), .B(n206), .Y(n901) );
  OAI21X1 U1094 ( .A(n197), .B(n902), .C(n901), .Y(n903) );
  OAI21X1 U1095 ( .A(n904), .B(n903), .C(n944), .Y(n906) );
  NAND2X1 U1096 ( .A(n945), .B(n20), .Y(n905) );
  NAND3X1 U1097 ( .A(n907), .B(n906), .C(n905), .Y(n910) );
  NOR2X1 U1098 ( .A(n230), .B(n908), .Y(n909) );
  AOI21X1 U1099 ( .A(n91), .B(n910), .C(n909), .Y(n913) );
  AOI22X1 U1100 ( .A(n911), .B(n235), .C(currentPlainKey[37]), .D(n216), .Y(
        n912) );
  NAND2X1 U1101 ( .A(n913), .B(n912), .Y(n1295) );
  AOI22X1 U1102 ( .A(n945), .B(n226), .C(currentPlainKey[38]), .D(n216), .Y(
        n929) );
  NAND2X1 U1103 ( .A(n143), .B(n167), .Y(n1007) );
  OAI21X1 U1104 ( .A(n1185), .B(n181), .C(currentPlainKey[38]), .Y(n914) );
  OAI21X1 U1105 ( .A(n1490), .B(n182), .C(n914), .Y(n916) );
  NOR2X1 U1106 ( .A(n221), .B(n1007), .Y(n915) );
  AOI21X1 U1107 ( .A(n33), .B(n916), .C(n915), .Y(n918) );
  NAND2X1 U1108 ( .A(n1010), .B(n236), .Y(n917) );
  OAI21X1 U1109 ( .A(n993), .B(n918), .C(n917), .Y(n919) );
  NAND2X1 U1110 ( .A(n224), .B(n919), .Y(n922) );
  NAND2X1 U1111 ( .A(n993), .B(n200), .Y(n921) );
  AOI21X1 U1112 ( .A(n922), .B(n921), .C(n920), .Y(n923) );
  MUX2X1 U1113 ( .B(n923), .A(n210), .S(n978), .Y(n925) );
  NAND2X1 U1114 ( .A(n961), .B(n212), .Y(n924) );
  NAND2X1 U1115 ( .A(n925), .B(n924), .Y(n927) );
  MUX2X1 U1116 ( .B(n927), .A(n232), .S(n926), .Y(n928) );
  NAND2X1 U1117 ( .A(n929), .B(n928), .Y(n1294) );
  NAND2X1 U1118 ( .A(n993), .B(n208), .Y(n940) );
  OAI21X1 U1119 ( .A(n166), .B(n181), .C(currentPlainKey[39]), .Y(n930) );
  OAI21X1 U1120 ( .A(n1361), .B(n182), .C(n930), .Y(n932) );
  NAND3X1 U1121 ( .A(n33), .B(n225), .C(n932), .Y(n933) );
  NAND2X1 U1122 ( .A(n143), .B(n89), .Y(n969) );
  INVX2 U1123 ( .A(n969), .Y(n1043) );
  MUX2X1 U1124 ( .B(n933), .A(n195), .S(n1043), .Y(n937) );
  INVX2 U1125 ( .A(n1007), .Y(n1025) );
  NAND2X1 U1126 ( .A(n1025), .B(n206), .Y(n934) );
  OAI21X1 U1127 ( .A(n197), .B(n935), .C(n934), .Y(n936) );
  OAI21X1 U1128 ( .A(n937), .B(n936), .C(n35), .Y(n939) );
  NAND2X1 U1129 ( .A(n978), .B(n213), .Y(n938) );
  NAND3X1 U1130 ( .A(n940), .B(n939), .C(n938), .Y(n943) );
  NOR2X1 U1131 ( .A(n230), .B(n941), .Y(n942) );
  AOI21X1 U1132 ( .A(n944), .B(n943), .C(n942), .Y(n947) );
  AOI22X1 U1133 ( .A(n945), .B(n232), .C(currentPlainKey[39]), .D(n216), .Y(
        n946) );
  NAND2X1 U1134 ( .A(n947), .B(n946), .Y(n1293) );
  AOI22X1 U1135 ( .A(n978), .B(n226), .C(currentPlainKey[40]), .D(n216), .Y(
        n964) );
  NAND2X1 U1136 ( .A(n143), .B(n152), .Y(n1039) );
  NAND2X1 U1137 ( .A(n969), .B(n1039), .Y(n1019) );
  INVX2 U1138 ( .A(n1019), .Y(n1042) );
  NAND3X1 U1139 ( .A(n192), .B(address[5]), .C(n948), .Y(n1063) );
  OAI21X1 U1140 ( .A(n1081), .B(n184), .C(currentPlainKey[40]), .Y(n949) );
  OAI21X1 U1141 ( .A(n1083), .B(n185), .C(n949), .Y(n951) );
  NOR2X1 U1142 ( .A(n221), .B(n1039), .Y(n950) );
  AOI21X1 U1143 ( .A(n1042), .B(n951), .C(n950), .Y(n953) );
  NAND2X1 U1144 ( .A(n1043), .B(n236), .Y(n952) );
  OAI21X1 U1145 ( .A(n1025), .B(n953), .C(n952), .Y(n954) );
  NAND2X1 U1146 ( .A(n225), .B(n954), .Y(n957) );
  NAND2X1 U1147 ( .A(n1025), .B(n201), .Y(n956) );
  AOI21X1 U1148 ( .A(n957), .B(n956), .C(n955), .Y(n958) );
  MUX2X1 U1149 ( .B(n958), .A(n209), .S(n1010), .Y(n960) );
  NAND2X1 U1150 ( .A(n993), .B(n212), .Y(n959) );
  NAND2X1 U1151 ( .A(n960), .B(n959), .Y(n962) );
  MUX2X1 U1152 ( .B(n962), .A(n234), .S(n961), .Y(n963) );
  NAND2X1 U1153 ( .A(n964), .B(n963), .Y(n1292) );
  NAND2X1 U1154 ( .A(n1025), .B(n209), .Y(n974) );
  OAI21X1 U1155 ( .A(n170), .B(n184), .C(currentPlainKey[41]), .Y(n965) );
  OAI21X1 U1156 ( .A(n1402), .B(n185), .C(n965), .Y(n966) );
  NAND3X1 U1157 ( .A(n1042), .B(n225), .C(n966), .Y(n967) );
  NAND2X1 U1158 ( .A(n1080), .B(n131), .Y(n1001) );
  INVX2 U1159 ( .A(n1001), .Y(n1077) );
  MUX2X1 U1160 ( .B(n967), .A(n196), .S(n1077), .Y(n971) );
  INVX2 U1161 ( .A(n1039), .Y(n1058) );
  NAND2X1 U1162 ( .A(n1058), .B(n206), .Y(n968) );
  OAI21X1 U1163 ( .A(n197), .B(n969), .C(n968), .Y(n970) );
  OAI21X1 U1164 ( .A(n971), .B(n970), .C(n33), .Y(n973) );
  NAND2X1 U1165 ( .A(n1010), .B(n212), .Y(n972) );
  NAND3X1 U1166 ( .A(n974), .B(n973), .C(n972), .Y(n977) );
  NOR2X1 U1167 ( .A(n229), .B(n975), .Y(n976) );
  AOI21X1 U1168 ( .A(n35), .B(n977), .C(n976), .Y(n980) );
  AOI22X1 U1169 ( .A(n978), .B(n234), .C(currentPlainKey[41]), .D(n216), .Y(
        n979) );
  NAND2X1 U1170 ( .A(n980), .B(n979), .Y(n1291) );
  AOI22X1 U1171 ( .A(n1010), .B(n226), .C(currentPlainKey[42]), .D(n216), .Y(
        n996) );
  NAND2X1 U1172 ( .A(n1080), .B(n1422), .Y(n1073) );
  NAND2X1 U1173 ( .A(n1001), .B(n1073), .Y(n1052) );
  INVX2 U1174 ( .A(n1052), .Y(n1076) );
  OAI21X1 U1175 ( .A(n25), .B(n184), .C(currentPlainKey[42]), .Y(n981) );
  OAI21X1 U1176 ( .A(n1118), .B(n185), .C(n981), .Y(n983) );
  NOR2X1 U1177 ( .A(n221), .B(n1073), .Y(n982) );
  AOI21X1 U1178 ( .A(n1076), .B(n983), .C(n982), .Y(n985) );
  NAND2X1 U1179 ( .A(n1077), .B(n236), .Y(n984) );
  OAI21X1 U1180 ( .A(n1058), .B(n985), .C(n984), .Y(n986) );
  NAND2X1 U1181 ( .A(n222), .B(n986), .Y(n989) );
  NAND2X1 U1182 ( .A(n1058), .B(n202), .Y(n988) );
  AOI21X1 U1183 ( .A(n989), .B(n988), .C(n987), .Y(n990) );
  MUX2X1 U1184 ( .B(n990), .A(n208), .S(n1043), .Y(n992) );
  NAND2X1 U1185 ( .A(n1025), .B(n212), .Y(n991) );
  NAND2X1 U1186 ( .A(n992), .B(n991), .Y(n994) );
  MUX2X1 U1187 ( .B(n994), .A(n51), .S(n993), .Y(n995) );
  NAND2X1 U1188 ( .A(n996), .B(n995), .Y(n1290) );
  NAND2X1 U1189 ( .A(n1058), .B(n210), .Y(n1006) );
  OAI21X1 U1190 ( .A(n164), .B(n184), .C(currentPlainKey[43]), .Y(n997) );
  OAI21X1 U1191 ( .A(n1135), .B(n185), .C(n997), .Y(n998) );
  NAND3X1 U1192 ( .A(n1076), .B(n225), .C(n998), .Y(n999) );
  NAND2X1 U1193 ( .A(n1080), .B(n121), .Y(n1033) );
  INVX2 U1194 ( .A(n1033), .Y(n1113) );
  MUX2X1 U1195 ( .B(n999), .A(n195), .S(n1113), .Y(n1003) );
  INVX2 U1196 ( .A(n1073), .Y(n1095) );
  NAND2X1 U1197 ( .A(n1095), .B(n206), .Y(n1000) );
  OAI21X1 U1198 ( .A(n198), .B(n1001), .C(n1000), .Y(n1002) );
  OAI21X1 U1199 ( .A(n1003), .B(n1002), .C(n1042), .Y(n1005) );
  NAND2X1 U1200 ( .A(n1043), .B(n212), .Y(n1004) );
  NAND3X1 U1201 ( .A(n1006), .B(n1005), .C(n1004), .Y(n1009) );
  NOR2X1 U1202 ( .A(n230), .B(n1007), .Y(n1008) );
  AOI21X1 U1203 ( .A(n33), .B(n1009), .C(n1008), .Y(n1012) );
  AOI22X1 U1204 ( .A(n1010), .B(n234), .C(currentPlainKey[43]), .D(n216), .Y(
        n1011) );
  NAND2X1 U1205 ( .A(n1012), .B(n1011), .Y(n1289) );
  AOI22X1 U1206 ( .A(n1043), .B(n226), .C(currentPlainKey[44]), .D(n216), .Y(
        n1028) );
  NAND2X1 U1207 ( .A(n1080), .B(n127), .Y(n1110) );
  OAI21X1 U1208 ( .A(n63), .B(n184), .C(currentPlainKey[44]), .Y(n1013) );
  OAI21X1 U1209 ( .A(n1455), .B(n185), .C(n1013), .Y(n1015) );
  NOR2X1 U1210 ( .A(n221), .B(n1110), .Y(n1014) );
  AOI21X1 U1211 ( .A(n57), .B(n1015), .C(n1014), .Y(n1017) );
  NAND2X1 U1212 ( .A(n1113), .B(n236), .Y(n1016) );
  OAI21X1 U1213 ( .A(n1095), .B(n1017), .C(n1016), .Y(n1018) );
  NAND2X1 U1214 ( .A(n224), .B(n1018), .Y(n1021) );
  NAND2X1 U1215 ( .A(n1095), .B(n203), .Y(n1020) );
  AOI21X1 U1216 ( .A(n1021), .B(n1020), .C(n1019), .Y(n1022) );
  MUX2X1 U1217 ( .B(n1022), .A(n208), .S(n1077), .Y(n1024) );
  NAND2X1 U1218 ( .A(n1058), .B(n20), .Y(n1023) );
  NAND2X1 U1219 ( .A(n1024), .B(n1023), .Y(n1026) );
  MUX2X1 U1220 ( .B(n1026), .A(n233), .S(n1025), .Y(n1027) );
  NAND2X1 U1221 ( .A(n1028), .B(n1027), .Y(n1288) );
  NAND2X1 U1222 ( .A(n1095), .B(n162), .Y(n1038) );
  OAI21X1 U1223 ( .A(n168), .B(n184), .C(currentPlainKey[45]), .Y(n1029) );
  OAI21X1 U1224 ( .A(n1478), .B(n185), .C(n1029), .Y(n1030) );
  NAND3X1 U1225 ( .A(n57), .B(n224), .C(n1030), .Y(n1031) );
  NAND2X1 U1226 ( .A(n1080), .B(n123), .Y(n1067) );
  INVX2 U1227 ( .A(n1067), .Y(n1148) );
  MUX2X1 U1228 ( .B(n1031), .A(n195), .S(n1148), .Y(n1035) );
  INVX2 U1229 ( .A(n1110), .Y(n1130) );
  NAND2X1 U1230 ( .A(n1130), .B(n206), .Y(n1032) );
  OAI21X1 U1231 ( .A(n197), .B(n1033), .C(n1032), .Y(n1034) );
  OAI21X1 U1232 ( .A(n1035), .B(n1034), .C(n1076), .Y(n1037) );
  NAND2X1 U1233 ( .A(n1077), .B(n212), .Y(n1036) );
  NAND3X1 U1234 ( .A(n1038), .B(n1037), .C(n1036), .Y(n1041) );
  NOR2X1 U1235 ( .A(n229), .B(n1039), .Y(n1040) );
  AOI21X1 U1236 ( .A(n1042), .B(n1041), .C(n1040), .Y(n1045) );
  AOI22X1 U1237 ( .A(n1043), .B(n232), .C(currentPlainKey[45]), .D(n216), .Y(
        n1044) );
  NAND2X1 U1238 ( .A(n1045), .B(n1044), .Y(n1287) );
  AOI22X1 U1239 ( .A(n1077), .B(n226), .C(currentPlainKey[46]), .D(n216), .Y(
        n1061) );
  NAND2X1 U1240 ( .A(n1080), .B(n125), .Y(n1145) );
  OAI21X1 U1241 ( .A(n1185), .B(n184), .C(currentPlainKey[46]), .Y(n1046) );
  OAI21X1 U1242 ( .A(n1490), .B(n185), .C(n1046), .Y(n1048) );
  NOR2X1 U1243 ( .A(n221), .B(n1145), .Y(n1047) );
  AOI21X1 U1244 ( .A(n71), .B(n1048), .C(n1047), .Y(n1050) );
  NAND2X1 U1245 ( .A(n1148), .B(n236), .Y(n1049) );
  OAI21X1 U1246 ( .A(n1130), .B(n1050), .C(n1049), .Y(n1051) );
  NAND2X1 U1247 ( .A(n225), .B(n1051), .Y(n1054) );
  NAND2X1 U1248 ( .A(n1130), .B(n204), .Y(n1053) );
  AOI21X1 U1249 ( .A(n1054), .B(n1053), .C(n1052), .Y(n1055) );
  MUX2X1 U1250 ( .B(n1055), .A(n103), .S(n1113), .Y(n1057) );
  NAND2X1 U1251 ( .A(n1095), .B(n213), .Y(n1056) );
  NAND2X1 U1252 ( .A(n1057), .B(n1056), .Y(n1059) );
  MUX2X1 U1253 ( .B(n1059), .A(n233), .S(n1058), .Y(n1060) );
  NAND2X1 U1254 ( .A(n1061), .B(n1060), .Y(n1286) );
  NAND2X1 U1255 ( .A(n1130), .B(n209), .Y(n1072) );
  OAI21X1 U1256 ( .A(n166), .B(n184), .C(currentPlainKey[47]), .Y(n1062) );
  OAI21X1 U1257 ( .A(n1361), .B(n185), .C(n1062), .Y(n1064) );
  NAND3X1 U1258 ( .A(n71), .B(n224), .C(n1064), .Y(n1065) );
  NAND2X1 U1259 ( .A(n1080), .B(n93), .Y(n1104) );
  INVX2 U1260 ( .A(n1104), .Y(n1182) );
  MUX2X1 U1261 ( .B(n1065), .A(n196), .S(n1182), .Y(n1069) );
  NAND2X1 U1262 ( .A(n2), .B(n206), .Y(n1066) );
  OAI21X1 U1263 ( .A(n197), .B(n1067), .C(n1066), .Y(n1068) );
  OAI21X1 U1264 ( .A(n1069), .B(n1068), .C(n57), .Y(n1071) );
  NAND2X1 U1265 ( .A(n1113), .B(n213), .Y(n1070) );
  NAND3X1 U1266 ( .A(n1072), .B(n1071), .C(n1070), .Y(n1075) );
  NOR2X1 U1267 ( .A(n230), .B(n1073), .Y(n1074) );
  AOI21X1 U1268 ( .A(n1076), .B(n1075), .C(n1074), .Y(n1079) );
  AOI22X1 U1269 ( .A(n1077), .B(n235), .C(currentPlainKey[47]), .D(n217), .Y(
        n1078) );
  NAND2X1 U1270 ( .A(n1079), .B(n1078), .Y(n1285) );
  AOI22X1 U1271 ( .A(n1113), .B(n226), .C(currentPlainKey[48]), .D(n216), .Y(
        n1098) );
  NAND2X1 U1272 ( .A(n1080), .B(n133), .Y(n1179) );
  OAI21X1 U1273 ( .A(n1081), .B(n186), .C(currentPlainKey[48]), .Y(n1082) );
  OAI21X1 U1274 ( .A(n1083), .B(n187), .C(n1082), .Y(n1085) );
  NOR2X1 U1275 ( .A(n221), .B(n1179), .Y(n1084) );
  AOI21X1 U1276 ( .A(n97), .B(n1085), .C(n1084), .Y(n1087) );
  NAND2X1 U1277 ( .A(n1182), .B(n236), .Y(n1086) );
  OAI21X1 U1278 ( .A(n2), .B(n1087), .C(n1086), .Y(n1088) );
  NAND2X1 U1279 ( .A(n222), .B(n1088), .Y(n1091) );
  NAND2X1 U1280 ( .A(n2), .B(n200), .Y(n1090) );
  AOI21X1 U1281 ( .A(n1091), .B(n1090), .C(n1089), .Y(n1092) );
  MUX2X1 U1282 ( .B(n1092), .A(n210), .S(n1148), .Y(n1094) );
  NAND2X1 U1283 ( .A(n1130), .B(n212), .Y(n1093) );
  NAND2X1 U1284 ( .A(n1094), .B(n1093), .Y(n1096) );
  MUX2X1 U1285 ( .B(n1096), .A(n232), .S(n1095), .Y(n1097) );
  NAND2X1 U1286 ( .A(n1098), .B(n1097), .Y(n1284) );
  NAND2X1 U1287 ( .A(n2), .B(n208), .Y(n1109) );
  OAI21X1 U1288 ( .A(n170), .B(n186), .C(currentPlainKey[49]), .Y(n1099) );
  OAI21X1 U1289 ( .A(n1402), .B(n187), .C(n1099), .Y(n1100) );
  NAND3X1 U1290 ( .A(n97), .B(n224), .C(n1100), .Y(n1102) );
  NAND2X1 U1291 ( .A(n27), .B(n151), .Y(n1514) );
  NAND2X1 U1292 ( .A(n113), .B(n43), .Y(n1139) );
  INVX2 U1293 ( .A(n1139), .Y(n1375) );
  MUX2X1 U1294 ( .B(n1102), .A(n196), .S(n1375), .Y(n1106) );
  INVX2 U1295 ( .A(n1179), .Y(n1268) );
  NAND2X1 U1296 ( .A(n1268), .B(n206), .Y(n1103) );
  OAI21X1 U1297 ( .A(n197), .B(n1104), .C(n1103), .Y(n1105) );
  OAI21X1 U1298 ( .A(n1106), .B(n1105), .C(n71), .Y(n1108) );
  NAND2X1 U1299 ( .A(n1148), .B(n20), .Y(n1107) );
  NAND3X1 U1300 ( .A(n1109), .B(n1108), .C(n1107), .Y(n1112) );
  NOR2X1 U1301 ( .A(n229), .B(n4), .Y(n1111) );
  AOI21X1 U1302 ( .A(n57), .B(n1112), .C(n1111), .Y(n1115) );
  AOI22X1 U1303 ( .A(n1113), .B(n232), .C(currentPlainKey[49]), .D(n215), .Y(
        n1114) );
  NAND2X1 U1304 ( .A(n1115), .B(n1114), .Y(n1283) );
  AOI22X1 U1306 ( .A(n1148), .B(n226), .C(currentPlainKey[50]), .D(n215), .Y(
        n1133) );
  NAND2X1 U1307 ( .A(n113), .B(n169), .Y(n1371) );
  NAND2X1 U1308 ( .A(n1139), .B(n1371), .Y(n1192) );
  INVX2 U1309 ( .A(n1192), .Y(n1374) );
  OAI21X1 U1310 ( .A(n25), .B(n186), .C(currentPlainKey[50]), .Y(n1117) );
  OAI21X1 U1311 ( .A(n1118), .B(n187), .C(n1117), .Y(n1120) );
  NOR2X1 U1312 ( .A(n220), .B(n1371), .Y(n1119) );
  AOI21X1 U1313 ( .A(n1374), .B(n1120), .C(n1119), .Y(n1122) );
  NAND2X1 U1314 ( .A(n1375), .B(n236), .Y(n1121) );
  OAI21X1 U1315 ( .A(n1268), .B(n1122), .C(n1121), .Y(n1123) );
  NAND2X1 U1316 ( .A(n222), .B(n1123), .Y(n1126) );
  NAND2X1 U1317 ( .A(n1268), .B(n204), .Y(n1125) );
  AOI21X1 U1318 ( .A(n1126), .B(n1125), .C(n1124), .Y(n1127) );
  MUX2X1 U1319 ( .B(n1127), .A(n209), .S(n1182), .Y(n1129) );
  NAND2X1 U1320 ( .A(n2), .B(n214), .Y(n1128) );
  NAND2X1 U1321 ( .A(n1129), .B(n1128), .Y(n1131) );
  MUX2X1 U1322 ( .B(n1131), .A(n51), .S(n1130), .Y(n1132) );
  NAND2X1 U1323 ( .A(n1133), .B(n1132), .Y(n1282) );
  NAND2X1 U1324 ( .A(n1268), .B(n209), .Y(n1144) );
  OAI21X1 U1325 ( .A(n164), .B(n186), .C(currentPlainKey[51]), .Y(n1134) );
  OAI21X1 U1326 ( .A(n187), .B(n1135), .C(n1134), .Y(n1136) );
  NAND3X1 U1327 ( .A(n1374), .B(n222), .C(n1136), .Y(n1137) );
  NAND2X1 U1328 ( .A(n113), .B(n1420), .Y(n1172) );
  INVX2 U1329 ( .A(n1172), .Y(n1416) );
  MUX2X1 U1330 ( .B(n1137), .A(n196), .S(n1416), .Y(n1141) );
  NAND2X1 U1331 ( .A(n1394), .B(n206), .Y(n1138) );
  OAI21X1 U1332 ( .A(n197), .B(n1139), .C(n1138), .Y(n1140) );
  OAI21X1 U1333 ( .A(n1141), .B(n1140), .C(n97), .Y(n1143) );
  NAND2X1 U1334 ( .A(n1182), .B(n213), .Y(n1142) );
  NAND3X1 U1335 ( .A(n1144), .B(n1143), .C(n1142), .Y(n1147) );
  NOR2X1 U1336 ( .A(n230), .B(n1145), .Y(n1146) );
  AOI21X1 U1337 ( .A(n71), .B(n1147), .C(n1146), .Y(n1150) );
  AOI22X1 U1338 ( .A(n1148), .B(n231), .C(currentPlainKey[51]), .D(n215), .Y(
        n1149) );
  NAND2X1 U1339 ( .A(n1150), .B(n1149), .Y(n1281) );
  AOI22X1 U1340 ( .A(n1182), .B(n227), .C(currentPlainKey[52]), .D(n215), .Y(
        n1166) );
  NAND2X1 U1341 ( .A(n113), .B(n163), .Y(n1170) );
  NAND2X1 U1342 ( .A(n1172), .B(n1170), .Y(n1388) );
  INVX2 U1343 ( .A(n1388), .Y(n1412) );
  OAI21X1 U1344 ( .A(n63), .B(n187), .C(currentPlainKey[52]), .Y(n1152) );
  OAI21X1 U1345 ( .A(n1455), .B(n186), .C(n1152), .Y(n1154) );
  NOR2X1 U1346 ( .A(n220), .B(n1170), .Y(n1153) );
  AOI21X1 U1347 ( .A(n1412), .B(n1154), .C(n1153), .Y(n1156) );
  NAND2X1 U1348 ( .A(n1416), .B(n236), .Y(n1155) );
  OAI21X1 U1349 ( .A(n1394), .B(n1156), .C(n1155), .Y(n1157) );
  NAND2X1 U1350 ( .A(n225), .B(n1157), .Y(n1160) );
  NAND2X1 U1351 ( .A(n1394), .B(n203), .Y(n1159) );
  AOI21X1 U1358 ( .A(n1160), .B(n1159), .C(n1158), .Y(n1161) );
  MUX2X1 U1359 ( .B(n1161), .A(n208), .S(n1375), .Y(n1163) );
  NAND2X1 U1360 ( .A(n1268), .B(n19), .Y(n1162) );
  NAND2X1 U1361 ( .A(n1163), .B(n1162), .Y(n1164) );
  MUX2X1 U1362 ( .B(n1164), .A(n233), .S(n2), .Y(n1165) );
  NAND2X1 U1363 ( .A(n1166), .B(n1165), .Y(n1280) );
  NAND2X1 U1364 ( .A(n1394), .B(n105), .Y(n1177) );
  OAI21X1 U1365 ( .A(n168), .B(n187), .C(currentPlainKey[53]), .Y(n1167) );
  OAI21X1 U1366 ( .A(n1478), .B(n186), .C(n1167), .Y(n1168) );
  NAND3X1 U1367 ( .A(n1412), .B(n224), .C(n1168), .Y(n1169) );
  NAND2X1 U1368 ( .A(n113), .B(n61), .Y(n1365) );
  INVX2 U1369 ( .A(n1365), .Y(n1451) );
  MUX2X1 U1370 ( .B(n1169), .A(n196), .S(n1451), .Y(n1174) );
  INVX2 U1371 ( .A(n1170), .Y(n1433) );
  NAND2X1 U1372 ( .A(n1433), .B(n207), .Y(n1171) );
  OAI21X1 U1373 ( .A(n197), .B(n1172), .C(n1171), .Y(n1173) );
  OAI21X1 U1374 ( .A(n1174), .B(n1173), .C(n1374), .Y(n1176) );
  NAND2X1 U1375 ( .A(n1375), .B(n213), .Y(n1175) );
  NAND3X1 U1376 ( .A(n1177), .B(n1176), .C(n1175), .Y(n1181) );
  NOR2X1 U1377 ( .A(n230), .B(n1179), .Y(n1180) );
  AOI21X1 U1378 ( .A(n97), .B(n1181), .C(n1180), .Y(n1184) );
  AOI22X1 U1379 ( .A(n1182), .B(n231), .C(currentPlainKey[53]), .D(n215), .Y(
        n1183) );
  NAND2X1 U1380 ( .A(n1184), .B(n1183), .Y(n1279) );
  AOI22X1 U1381 ( .A(n1375), .B(n226), .C(currentPlainKey[54]), .D(n215), .Y(
        n1359) );
  NAND2X1 U1382 ( .A(n113), .B(n167), .Y(n1383) );
  OAI21X1 U1383 ( .A(n1185), .B(n187), .C(currentPlainKey[54]), .Y(n1186) );
  OAI21X1 U1384 ( .A(n186), .B(n1490), .C(n1186), .Y(n1188) );
  NOR2X1 U1385 ( .A(n220), .B(n1383), .Y(n1187) );
  AOI21X1 U1386 ( .A(n79), .B(n1188), .C(n1187), .Y(n1190) );
  NAND2X1 U1387 ( .A(n1451), .B(n236), .Y(n1189) );
  OAI21X1 U1388 ( .A(n1433), .B(n1190), .C(n1189), .Y(n1191) );
  NAND2X1 U1389 ( .A(n222), .B(n1191), .Y(n1194) );
  NAND2X1 U1390 ( .A(n1433), .B(n200), .Y(n1193) );
  AOI21X1 U1391 ( .A(n1194), .B(n1193), .C(n1192), .Y(n1195) );
  MUX2X1 U1392 ( .B(n1195), .A(n103), .S(n1416), .Y(n1267) );
  NAND2X1 U1393 ( .A(n1394), .B(n214), .Y(n1196) );
  NAND2X1 U1394 ( .A(n1267), .B(n1196), .Y(n1357) );
  MUX2X1 U1395 ( .B(n1357), .A(n232), .S(n1268), .Y(n1358) );
  NAND2X1 U1396 ( .A(n1359), .B(n1358), .Y(n1278) );
  NAND2X1 U1397 ( .A(n1433), .B(n210), .Y(n1370) );
  OAI21X1 U1398 ( .A(n166), .B(n186), .C(currentPlainKey[55]), .Y(n1360) );
  OAI21X1 U1399 ( .A(n187), .B(n1361), .C(n1360), .Y(n1362) );
  NAND3X1 U1400 ( .A(n79), .B(n222), .C(n1362), .Y(n1363) );
  NAND2X1 U1401 ( .A(n113), .B(n89), .Y(n1380) );
  INVX2 U1402 ( .A(n1380), .Y(n1486) );
  MUX2X1 U1403 ( .B(n1363), .A(n196), .S(n1486), .Y(n1367) );
  INVX2 U1404 ( .A(n1383), .Y(n1468) );
  NAND2X1 U1405 ( .A(n207), .B(n1468), .Y(n1364) );
  OAI21X1 U1406 ( .A(n1365), .B(n197), .C(n1364), .Y(n1366) );
  OAI21X1 U1407 ( .A(n1367), .B(n1366), .C(n1412), .Y(n1369) );
  NAND2X1 U1408 ( .A(n1416), .B(n214), .Y(n1368) );
  NAND3X1 U1409 ( .A(n1370), .B(n1369), .C(n1368), .Y(n1373) );
  NOR2X1 U1410 ( .A(n229), .B(n1371), .Y(n1372) );
  AOI21X1 U1411 ( .A(n1374), .B(n1373), .C(n1372), .Y(n1377) );
  AOI22X1 U1412 ( .A(n1375), .B(n231), .C(currentPlainKey[55]), .D(n215), .Y(
        n1376) );
  NAND2X1 U1413 ( .A(n1377), .B(n1376), .Y(n1277) );
  AOI22X1 U1414 ( .A(n1416), .B(n226), .C(currentPlainKey[56]), .D(n215), .Y(
        n1397) );
  NAND2X1 U1415 ( .A(n1486), .B(n236), .Y(n1386) );
  NAND2X1 U1416 ( .A(n193), .B(n151), .Y(n1511) );
  INVX2 U1417 ( .A(n1511), .Y(n1491) );
  NAND2X1 U1418 ( .A(n1491), .B(n43), .Y(n1379) );
  AOI22X1 U1419 ( .A(currentPlainKey[56]), .B(n1379), .C(n1378), .D(n1491), 
        .Y(n1382) );
  NAND2X1 U1420 ( .A(n113), .B(n152), .Y(n1438) );
  NAND2X1 U1421 ( .A(n1380), .B(n1438), .Y(n1398) );
  NAND2X1 U1422 ( .A(n1504), .B(n190), .Y(n1381) );
  OAI21X1 U1423 ( .A(n1382), .B(n1398), .C(n1381), .Y(n1384) );
  NAND2X1 U1424 ( .A(n1384), .B(n1383), .Y(n1385) );
  NAND2X1 U1425 ( .A(n1386), .B(n1385), .Y(n1387) );
  NAND2X1 U1426 ( .A(n225), .B(n1387), .Y(n1390) );
  NAND2X1 U1427 ( .A(n203), .B(n1468), .Y(n1389) );
  AOI21X1 U1428 ( .A(n1390), .B(n1389), .C(n1388), .Y(n1391) );
  MUX2X1 U1429 ( .B(n1391), .A(n103), .S(n1451), .Y(n1393) );
  NAND2X1 U1430 ( .A(n1433), .B(n212), .Y(n1392) );
  NAND2X1 U1431 ( .A(n1393), .B(n1392), .Y(n1395) );
  MUX2X1 U1432 ( .B(n1395), .A(n51), .S(n8), .Y(n1396) );
  NAND2X1 U1433 ( .A(n1396), .B(n1397), .Y(n1276) );
  NAND2X1 U1434 ( .A(n1433), .B(n226), .Y(n1419) );
  NAND2X1 U1435 ( .A(n1495), .B(n131), .Y(n1405) );
  OAI21X1 U1436 ( .A(n170), .B(n16), .C(currentPlainKey[57]), .Y(n1401) );
  OAI21X1 U1437 ( .A(n16), .B(n1402), .C(n1401), .Y(n1403) );
  NAND2X1 U1438 ( .A(n55), .B(n1403), .Y(n1404) );
  NAND2X1 U1439 ( .A(n1468), .B(n162), .Y(n1409) );
  NAND2X1 U1440 ( .A(n1451), .B(n211), .Y(n1410) );
  NAND3X1 U1441 ( .A(n1404), .B(n1409), .C(n1410), .Y(n1415) );
  NAND2X1 U1442 ( .A(n207), .B(n1504), .Y(n1408) );
  INVX2 U1443 ( .A(n1405), .Y(n1531) );
  NAND2X1 U1444 ( .A(n1531), .B(n111), .Y(n1446) );
  INVX2 U1445 ( .A(n1446), .Y(n1485) );
  NAND2X1 U1446 ( .A(n1485), .B(n190), .Y(n1407) );
  NAND2X1 U1447 ( .A(n201), .B(n1486), .Y(n1406) );
  NAND3X1 U1448 ( .A(n1408), .B(n1407), .C(n1406), .Y(n1414) );
  NAND3X1 U1449 ( .A(n1410), .B(n1409), .C(n1427), .Y(n1411) );
  AND2X2 U1450 ( .A(n1412), .B(n1411), .Y(n1413) );
  OAI21X1 U1451 ( .A(n1415), .B(n1414), .C(n1413), .Y(n1418) );
  AOI22X1 U1452 ( .A(n1416), .B(n231), .C(currentPlainKey[57]), .D(n215), .Y(
        n1417) );
  NAND3X1 U1453 ( .A(n1419), .B(n1418), .C(n1417), .Y(n1275) );
  AOI22X1 U1454 ( .A(n1451), .B(n226), .C(currentPlainKey[58]), .D(n215), .Y(
        n1436) );
  NAND2X1 U1455 ( .A(n204), .B(n1504), .Y(n1429) );
  NAND2X1 U1456 ( .A(n1420), .B(n1491), .Y(n1421) );
  AOI22X1 U1457 ( .A(currentPlainKey[58]), .B(n1421), .C(n73), .D(n1491), .Y(
        n1423) );
  NAND2X1 U1458 ( .A(n1422), .B(n1495), .Y(n1458) );
  MUX2X1 U1459 ( .B(n1423), .A(n220), .S(n1528), .Y(n1424) );
  NAND2X1 U1460 ( .A(n1424), .B(n1438), .Y(n1425) );
  MUX2X1 U1461 ( .B(n1425), .A(n238), .S(n1531), .Y(n1426) );
  NAND2X1 U1462 ( .A(n225), .B(n1426), .Y(n1428) );
  AOI21X1 U1463 ( .A(n1429), .B(n1428), .C(n1427), .Y(n1430) );
  NAND2X1 U1464 ( .A(n1468), .B(n213), .Y(n1431) );
  NAND2X1 U1465 ( .A(n1432), .B(n1431), .Y(n1434) );
  MUX2X1 U1466 ( .B(n1434), .A(n234), .S(n1433), .Y(n1435) );
  NAND2X1 U1467 ( .A(n1435), .B(n1436), .Y(n1274) );
  NAND2X1 U1468 ( .A(n1468), .B(n226), .Y(n1454) );
  NAND2X1 U1469 ( .A(n1486), .B(n213), .Y(n1437) );
  OAI21X1 U1470 ( .A(n1439), .B(n1438), .C(n1437), .Y(n1450) );
  NOR2X1 U1471 ( .A(n238), .B(n1458), .Y(n1445) );
  NOR2X1 U1472 ( .A(n16), .B(n164), .Y(n1441) );
  MUX2X1 U1473 ( .B(n1635), .A(n188), .S(n1441), .Y(n1442) );
  NAND2X1 U1474 ( .A(n1442), .B(n1458), .Y(n1443) );
  NAND2X1 U1475 ( .A(n121), .B(n1495), .Y(n1459) );
  INVX2 U1476 ( .A(n1459), .Y(n1523) );
  MUX2X1 U1477 ( .B(n1443), .A(n220), .S(n1523), .Y(n1444) );
  NOR2X1 U1478 ( .A(n1445), .B(n1444), .Y(n1448) );
  OAI22X1 U1479 ( .A(n1448), .B(n1447), .C(n1520), .D(n1446), .Y(n1449) );
  OAI21X1 U1480 ( .A(n1450), .B(n1449), .C(n79), .Y(n1453) );
  AOI22X1 U1481 ( .A(n1451), .B(n231), .C(currentPlainKey[59]), .D(n215), .Y(
        n1452) );
  NAND3X1 U1482 ( .A(n1454), .B(n1453), .C(n1452), .Y(n1273) );
  AOI22X1 U1483 ( .A(n1486), .B(n226), .C(currentPlainKey[60]), .D(n215), .Y(
        n1471) );
  NAND2X1 U1484 ( .A(n1531), .B(n103), .Y(n1467) );
  AOI22X1 U1485 ( .A(n1523), .B(n236), .C(n1528), .D(RCV_DATA[3]), .Y(n1463)
         );
  NAND2X1 U1486 ( .A(n61), .B(n1491), .Y(n1457) );
  INVX2 U1487 ( .A(n1455), .Y(n1456) );
  AOI22X1 U1488 ( .A(currentPlainKey[60]), .B(n1457), .C(n1456), .D(n1491), 
        .Y(n1460) );
  NAND2X1 U1489 ( .A(n1459), .B(n1458), .Y(n1472) );
  NOR2X1 U1490 ( .A(n1460), .B(n1472), .Y(n1461) );
  NAND2X1 U1491 ( .A(n127), .B(n1495), .Y(n1474) );
  INVX2 U1492 ( .A(n1474), .Y(n1521) );
  MUX2X1 U1493 ( .B(n1461), .A(n190), .S(n1521), .Y(n1462) );
  NAND2X1 U1494 ( .A(n1463), .B(n1462), .Y(n1464) );
  NAND2X1 U1495 ( .A(n55), .B(n1464), .Y(n1466) );
  NAND2X1 U1496 ( .A(n214), .B(n1504), .Y(n1465) );
  NAND3X1 U1497 ( .A(n1467), .B(n1466), .C(n1465), .Y(n1469) );
  MUX2X1 U1498 ( .B(n1469), .A(n233), .S(n1468), .Y(n1470) );
  NAND2X1 U1499 ( .A(n1471), .B(n1470), .Y(n1272) );
  NAND2X1 U1500 ( .A(n123), .B(n1495), .Y(n1518) );
  INVX2 U1501 ( .A(n1472), .Y(n1473) );
  NAND3X1 U1502 ( .A(n1518), .B(n1474), .C(n1473), .Y(n1475) );
  INVX2 U1503 ( .A(n1475), .Y(n1499) );
  OAI21X1 U1504 ( .A(n16), .B(n168), .C(currentPlainKey[61]), .Y(n1477) );
  OAI21X1 U1505 ( .A(n16), .B(n1478), .C(n1477), .Y(n1480) );
  NOR2X1 U1506 ( .A(n220), .B(n1518), .Y(n1479) );
  AOI21X1 U1507 ( .A(n1499), .B(n1480), .C(n1479), .Y(n1483) );
  NAND2X1 U1508 ( .A(n1521), .B(n236), .Y(n1482) );
  AOI22X1 U1509 ( .A(n1523), .B(RCV_DATA[3]), .C(n1528), .D(RCV_DATA[4]), .Y(
        n1481) );
  NAND3X1 U1510 ( .A(n1483), .B(n1482), .C(n1481), .Y(n1484) );
  AOI22X1 U1511 ( .A(n1485), .B(RCV_DATA[5]), .C(n55), .D(n1484), .Y(n1489) );
  NAND2X1 U1512 ( .A(n227), .B(n1504), .Y(n1488) );
  AOI22X1 U1513 ( .A(n1486), .B(n231), .C(currentPlainKey[61]), .D(n215), .Y(
        n1487) );
  NAND3X1 U1514 ( .A(n1489), .B(n1488), .C(n1487), .Y(n1271) );
  AOI22X1 U1515 ( .A(n233), .B(n1504), .C(n219), .D(currentPlainKey[62]), .Y(
        n1509) );
  INVX2 U1516 ( .A(n1490), .Y(n1494) );
  AOI21X1 U1517 ( .A(n89), .B(n1491), .C(n1620), .Y(n1493) );
  NAND2X1 U1518 ( .A(n16), .B(n1620), .Y(n1492) );
  OAI21X1 U1519 ( .A(n1494), .B(n1493), .C(n1492), .Y(n1496) );
  MUX2X1 U1520 ( .B(n1496), .A(n220), .S(n115), .Y(n1498) );
  NOR2X1 U1521 ( .A(n238), .B(n1518), .Y(n1497) );
  AOI21X1 U1522 ( .A(n1499), .B(n1498), .C(n1497), .Y(n1501) );
  NAND2X1 U1523 ( .A(n1521), .B(RCV_DATA[3]), .Y(n1500) );
  NAND2X1 U1524 ( .A(n1501), .B(n1500), .Y(n1502) );
  AOI22X1 U1525 ( .A(n225), .B(n1502), .C(n1523), .D(n103), .Y(n1506) );
  NAND2X1 U1526 ( .A(n1528), .B(n19), .Y(n1505) );
  AOI21X1 U1527 ( .A(n1506), .B(n1505), .C(n1504), .Y(n1507) );
  MUX2X1 U1528 ( .B(n1507), .A(n226), .S(n1531), .Y(n1508) );
  NAND2X1 U1529 ( .A(n1509), .B(n1508), .Y(n1270) );
  NAND2X1 U1530 ( .A(n219), .B(currentPlainKey[63]), .Y(n1534) );
  NOR2X1 U1531 ( .A(n1511), .B(n166), .Y(n1512) );
  MUX2X1 U1532 ( .B(currentPlainKey[63]), .A(n189), .S(n1512), .Y(n1516) );
  NOR2X1 U1533 ( .A(n1514), .B(n1513), .Y(n1515) );
  MUX2X1 U1534 ( .B(n1516), .A(n220), .S(n1515), .Y(n1517) );
  MUX2X1 U1535 ( .B(n1517), .A(n236), .S(n115), .Y(n1519) );
  MUX2X1 U1536 ( .B(n1520), .A(n1519), .S(n1518), .Y(n1522) );
  MUX2X1 U1537 ( .B(n1522), .A(RCV_DATA[4]), .S(n1521), .Y(n1525) );
  INVX2 U1538 ( .A(RCV_DATA[5]), .Y(n1524) );
  MUX2X1 U1539 ( .B(n1525), .A(n1524), .S(n1523), .Y(n1526) );
  NAND2X1 U1540 ( .A(n224), .B(n1526), .Y(n1530) );
  MUX2X1 U1541 ( .B(n1530), .A(n230), .S(n1528), .Y(n1532) );
  MUX2X1 U1542 ( .B(n1532), .A(n51), .S(n1531), .Y(n1533) );
  NAND2X1 U1543 ( .A(n1534), .B(n1533), .Y(n1269) );
  NAND2X1 U1544 ( .A(n1535), .B(n1605), .Y(n1547) );
  INVX2 U1545 ( .A(n1547), .Y(n1536) );
  NAND3X1 U1546 ( .A(n17), .B(n253), .C(n1536), .Y(n1545) );
  NAND2X1 U1547 ( .A(address[0]), .B(n1545), .Y(n1537) );
  NAND2X1 U1548 ( .A(n1546), .B(n1537), .Y(n1333) );
  NAND2X1 U1549 ( .A(address[1]), .B(n1545), .Y(n1538) );
  NAND2X1 U1550 ( .A(n1546), .B(n1538), .Y(n1334) );
  NAND2X1 U1551 ( .A(address[2]), .B(n1545), .Y(n1539) );
  NAND2X1 U1552 ( .A(n1546), .B(n1539), .Y(n1335) );
  MUX2X1 U1553 ( .B(n192), .A(keyCount[0]), .S(n1542), .Y(n1540) );
  NAND2X1 U1554 ( .A(n1546), .B(n1540), .Y(n1336) );
  MUX2X1 U1555 ( .B(address[4]), .A(keyCount[1]), .S(n1542), .Y(n1541) );
  NAND2X1 U1556 ( .A(n1546), .B(n1541), .Y(n1337) );
  MUX2X1 U1557 ( .B(address[5]), .A(keyCount[2]), .S(n1542), .Y(n1543) );
  NAND2X1 U1558 ( .A(n1546), .B(n1543), .Y(n1338) );
  OAI21X1 U1559 ( .A(n1631), .B(n1544), .C(n1546), .Y(n1339) );
  OAI21X1 U1560 ( .A(n1630), .B(n1544), .C(n1546), .Y(n1340) );
  OAI21X1 U1561 ( .A(n1548), .B(n1547), .C(parityError), .Y(n1551) );
  OAI21X1 U1562 ( .A(n12), .B(n13), .C(n1549), .Y(n1550) );
  NAND2X1 U1563 ( .A(n1551), .B(n1550), .Y(nextParityError) );
  OAI21X1 U1564 ( .A(keyCount[0]), .B(n157), .C(n135), .Y(n1552) );
  INVX2 U1565 ( .A(n1552), .Y(n1607) );
  NAND2X1 U1566 ( .A(n1596), .B(n135), .Y(n1619) );
  INVX2 U1567 ( .A(n1619), .Y(n1610) );
  NAND2X1 U1568 ( .A(keyCount[0]), .B(n1610), .Y(n1615) );
  MUX2X1 U1569 ( .B(n1607), .A(n1615), .S(n1629), .Y(n1350) );
  NAND3X1 U1570 ( .A(n1597), .B(n14), .C(n17), .Y(n1555) );
  NAND3X1 U1571 ( .A(n101), .B(n253), .C(n11), .Y(n1554) );
  OR2X2 U1572 ( .A(n1555), .B(n1554), .Y(n1569) );
  NAND2X1 U1573 ( .A(n1565), .B(CLR_RBUFF), .Y(n1571) );
  INVX2 U1574 ( .A(n1571), .Y(n1566) );
  NAND2X1 U1575 ( .A(N1799), .B(n1566), .Y(n1557) );
  NAND2X1 U1576 ( .A(parityAccumulator[7]), .B(n1569), .Y(n1556) );
  NAND2X1 U1577 ( .A(n1557), .B(n1556), .Y(n1341) );
  NAND2X1 U1578 ( .A(N1798), .B(n1566), .Y(n1559) );
  NAND2X1 U1579 ( .A(parityAccumulator[6]), .B(n1569), .Y(n1558) );
  NAND2X1 U1580 ( .A(n1559), .B(n1558), .Y(n1342) );
  NAND2X1 U1581 ( .A(N1797), .B(n1566), .Y(n1561) );
  NAND2X1 U1582 ( .A(n1569), .B(parityAccumulator[5]), .Y(n1560) );
  NAND2X1 U1583 ( .A(n1561), .B(n1560), .Y(n1343) );
  NAND2X1 U1584 ( .A(N1796), .B(n1566), .Y(n1563) );
  NAND2X1 U1585 ( .A(n1569), .B(parityAccumulator[4]), .Y(n1562) );
  NAND2X1 U1586 ( .A(n1563), .B(n1562), .Y(n1344) );
  INVX2 U1587 ( .A(n1569), .Y(n1565) );
  NAND2X1 U1588 ( .A(N1795), .B(n1566), .Y(n1564) );
  OAI21X1 U1589 ( .A(n1626), .B(n1565), .C(n1564), .Y(n1345) );
  NAND2X1 U1590 ( .A(N1794), .B(n1566), .Y(n1567) );
  OAI21X1 U1591 ( .A(n1625), .B(n1565), .C(n1567), .Y(n1346) );
  INVX2 U1592 ( .A(N1793), .Y(n1568) );
  OAI22X1 U1593 ( .A(n1624), .B(n1565), .C(n1571), .D(n1568), .Y(n1347) );
  INVX2 U1594 ( .A(N1792), .Y(n1570) );
  OAI22X1 U1595 ( .A(n1623), .B(n1565), .C(n1571), .D(n1570), .Y(n1348) );
  AOI21X1 U1596 ( .A(n1580), .B(RBUF_FULL), .C(n1178), .Y(n1572) );
  NAND2X1 U1597 ( .A(n1572), .B(n1587), .Y(n1576) );
  NAND2X1 U1598 ( .A(n1574), .B(n1573), .Y(n1575) );
  NAND2X1 U1599 ( .A(n1575), .B(n1598), .Y(n1581) );
  NAND2X1 U1600 ( .A(n1576), .B(n1581), .Y(n1591) );
  NAND2X1 U1601 ( .A(n7), .B(n1591), .Y(n1577) );
  NAND2X1 U1602 ( .A(n1578), .B(n1577), .Y(n1354) );
  INVX2 U1603 ( .A(keyCount[3]), .Y(n1580) );
  AND2X2 U1604 ( .A(keyCount[2]), .B(keyCount[0]), .Y(n1579) );
  NAND3X1 U1605 ( .A(keyCount[1]), .B(n1580), .C(n1579), .Y(n1595) );
  INVX2 U1606 ( .A(n1595), .Y(n1611) );
  INVX2 U1607 ( .A(n1581), .Y(n1594) );
  AOI22X1 U1608 ( .A(n1611), .B(n1596), .C(n1594), .D(n9), .Y(n1590) );
  INVX2 U1609 ( .A(RBUF_FULL), .Y(n1582) );
  NAND2X1 U1610 ( .A(n1583), .B(n1582), .Y(n1589) );
  INVX2 U1611 ( .A(OE), .Y(n1584) );
  NAND2X1 U1612 ( .A(n1695), .B(n1584), .Y(n1586) );
  NAND2X1 U1613 ( .A(n1597), .B(n17), .Y(n1585) );
  AOI21X1 U1614 ( .A(n1587), .B(n1586), .C(n1585), .Y(n1588) );
  NAND3X1 U1615 ( .A(n1590), .B(n1589), .C(n1588), .Y(n1352) );
  AOI21X1 U1616 ( .A(n85), .B(n1591), .C(n1596), .Y(n1592) );
  NAND3X1 U1617 ( .A(n1597), .B(n47), .C(n1592), .Y(n1351) );
  AOI22X1 U1618 ( .A(n1596), .B(n1595), .C(n1594), .D(n194), .Y(n1606) );
  NAND2X1 U1619 ( .A(n1598), .B(n1597), .Y(n1603) );
  NAND2X1 U1620 ( .A(n1695), .B(n1584), .Y(n1601) );
  OAI21X1 U1621 ( .A(n1601), .B(n14), .C(n17), .Y(n1602) );
  AOI21X1 U1622 ( .A(RBUF_FULL), .B(n1603), .C(n1602), .Y(n1604) );
  NAND3X1 U1623 ( .A(n1606), .B(n1605), .C(n1604), .Y(n1353) );
  NOR2X1 U1624 ( .A(keyCount[2]), .B(n157), .Y(n1609) );
  OAI21X1 U1625 ( .A(keyCount[1]), .B(n157), .C(n1607), .Y(n1614) );
  OAI21X1 U1626 ( .A(n1609), .B(n1614), .C(keyCount[3]), .Y(n1613) );
  NAND2X1 U1627 ( .A(n1611), .B(n1610), .Y(n1612) );
  NAND2X1 U1628 ( .A(n1613), .B(n1612), .Y(n1355) );
  INVX2 U1629 ( .A(n1614), .Y(n1618) );
  INVX2 U1630 ( .A(n1615), .Y(n1616) );
  NAND2X1 U1631 ( .A(n1616), .B(keyCount[1]), .Y(n1617) );
  MUX2X1 U1632 ( .B(n1618), .A(n1617), .S(n1621), .Y(n1349) );
  MUX2X1 U1633 ( .B(n1619), .A(n135), .S(keyCount[0]), .Y(n1356) );
  INVX2 U1634 ( .A(keyCount[2]), .Y(n1621) );
  INVX2 U1635 ( .A(parityAccumulator[0]), .Y(n1623) );
  INVX2 U1636 ( .A(parityAccumulator[1]), .Y(n1624) );
  INVX2 U1637 ( .A(parityAccumulator[2]), .Y(n1625) );
  INVX2 U1638 ( .A(parityAccumulator[3]), .Y(n1626) );
  INVX2 U1639 ( .A(keyCount[1]), .Y(n1629) );
  INVX2 U1640 ( .A(address[7]), .Y(n1630) );
  INVX2 U1641 ( .A(address[6]), .Y(n1631) );
  INVX2 U1642 ( .A(currentPlainKey[61]), .Y(n1633) );
  INVX2 U1643 ( .A(currentPlainKey[60]), .Y(n1634) );
  INVX2 U1644 ( .A(currentPlainKey[59]), .Y(n1635) );
  INVX2 U1645 ( .A(currentPlainKey[58]), .Y(n1636) );
  INVX2 U1646 ( .A(currentPlainKey[57]), .Y(n1637) );
  INVX2 U1647 ( .A(currentPlainKey[56]), .Y(n1638) );
  INVX2 U1648 ( .A(currentPlainKey[55]), .Y(n1639) );
  INVX2 U1649 ( .A(currentPlainKey[54]), .Y(n1640) );
  INVX2 U1650 ( .A(currentPlainKey[53]), .Y(n1641) );
  INVX2 U1651 ( .A(currentPlainKey[52]), .Y(n1642) );
  INVX2 U1652 ( .A(currentPlainKey[51]), .Y(n1643) );
  INVX2 U1653 ( .A(currentPlainKey[50]), .Y(n1644) );
  INVX2 U1654 ( .A(currentPlainKey[49]), .Y(n1645) );
  INVX2 U1655 ( .A(currentPlainKey[48]), .Y(n1646) );
  INVX2 U1656 ( .A(currentPlainKey[47]), .Y(n1647) );
  INVX2 U1657 ( .A(currentPlainKey[46]), .Y(n1648) );
  INVX2 U1658 ( .A(currentPlainKey[45]), .Y(n1649) );
  INVX2 U1659 ( .A(currentPlainKey[44]), .Y(n1650) );
  INVX2 U1660 ( .A(currentPlainKey[43]), .Y(n1651) );
  INVX2 U1661 ( .A(currentPlainKey[42]), .Y(n1652) );
  INVX2 U1662 ( .A(currentPlainKey[41]), .Y(n1653) );
  INVX2 U1663 ( .A(currentPlainKey[40]), .Y(n1654) );
  INVX2 U1664 ( .A(currentPlainKey[39]), .Y(n1655) );
  INVX2 U1665 ( .A(currentPlainKey[38]), .Y(n1656) );
  INVX2 U1666 ( .A(currentPlainKey[37]), .Y(n1657) );
  INVX2 U1667 ( .A(currentPlainKey[36]), .Y(n1658) );
  INVX2 U1668 ( .A(currentPlainKey[35]), .Y(n1659) );
  INVX2 U1669 ( .A(currentPlainKey[34]), .Y(n1660) );
  INVX2 U1670 ( .A(currentPlainKey[33]), .Y(n1661) );
  INVX2 U1671 ( .A(currentPlainKey[32]), .Y(n1662) );
  INVX2 U1672 ( .A(currentPlainKey[31]), .Y(n1663) );
  INVX2 U1673 ( .A(currentPlainKey[30]), .Y(n1664) );
  INVX2 U1674 ( .A(currentPlainKey[29]), .Y(n1665) );
  INVX2 U1675 ( .A(currentPlainKey[28]), .Y(n1666) );
  INVX2 U1676 ( .A(currentPlainKey[27]), .Y(n1667) );
  INVX2 U1677 ( .A(currentPlainKey[26]), .Y(n1668) );
  INVX2 U1678 ( .A(currentPlainKey[25]), .Y(n1669) );
  INVX2 U1679 ( .A(currentPlainKey[24]), .Y(n1670) );
  INVX2 U1680 ( .A(currentPlainKey[23]), .Y(n1671) );
  INVX2 U1681 ( .A(currentPlainKey[22]), .Y(n1672) );
  INVX2 U1682 ( .A(currentPlainKey[21]), .Y(n1673) );
  INVX2 U1683 ( .A(currentPlainKey[20]), .Y(n1674) );
  INVX2 U1684 ( .A(currentPlainKey[19]), .Y(n1675) );
  INVX2 U1685 ( .A(currentPlainKey[18]), .Y(n1676) );
  INVX2 U1686 ( .A(currentPlainKey[17]), .Y(n1677) );
  INVX2 U1687 ( .A(currentPlainKey[16]), .Y(n1678) );
  INVX2 U1688 ( .A(currentPlainKey[15]), .Y(n1679) );
  INVX2 U1689 ( .A(currentPlainKey[14]), .Y(n1680) );
  INVX2 U1690 ( .A(currentPlainKey[13]), .Y(n1681) );
  INVX2 U1691 ( .A(currentPlainKey[12]), .Y(n1682) );
  INVX2 U1692 ( .A(currentPlainKey[11]), .Y(n1683) );
  INVX2 U1693 ( .A(currentPlainKey[10]), .Y(n1684) );
  INVX2 U1694 ( .A(currentPlainKey[9]), .Y(n1685) );
  INVX2 U1695 ( .A(currentPlainKey[8]), .Y(n1686) );
  INVX2 U1696 ( .A(currentPlainKey[7]), .Y(n1687) );
  INVX2 U1697 ( .A(currentPlainKey[6]), .Y(n1688) );
  INVX2 U1698 ( .A(currentPlainKey[5]), .Y(n1689) );
  INVX2 U1699 ( .A(currentPlainKey[4]), .Y(n1690) );
  INVX2 U1700 ( .A(SBE), .Y(n1695) );
endmodule


module uart_timer_1_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module uart_timer_1 ( CLK, RST, TIMER_TRIG, STOP_RCVING, SHIFT_STROBE );
  input CLK, RST, TIMER_TRIG;
  output STOP_RCVING, SHIFT_STROBE;
  wire   N26, N27, N28, N29, N30, N31, N32, N33, N60, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n17, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34;
  wire   [7:0] state;
  wire   [7:0] nextState;
  assign SHIFT_STROBE = N60;

  DFFSR \nextState_reg[0]  ( .D(n71), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[0]) );
  DFFSR \nextState_reg[1]  ( .D(n70), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[1]) );
  DFFSR \nextState_reg[2]  ( .D(n69), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[2]) );
  DFFSR \nextState_reg[3]  ( .D(n68), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[3]) );
  DFFSR \nextState_reg[4]  ( .D(n67), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[4]) );
  DFFSR \nextState_reg[5]  ( .D(n66), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[5]) );
  DFFSR \nextState_reg[6]  ( .D(n65), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[6]) );
  DFFSR STOP_RCVING_reg ( .D(n72), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        STOP_RCVING) );
  DFFSR \state_reg[7]  ( .D(nextState[7]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[7]) );
  DFFSR \state_reg[6]  ( .D(nextState[6]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[6]) );
  DFFSR \state_reg[5]  ( .D(nextState[5]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[5]) );
  DFFSR \state_reg[4]  ( .D(nextState[4]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[3]  ( .D(nextState[3]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[0]) );
  OR2X2 U21 ( .A(state[7]), .B(n50), .Y(n49) );
  OAI21X1 U38 ( .A(n20), .B(n27), .C(n35), .Y(n64) );
  NAND2X1 U39 ( .A(N33), .B(n36), .Y(n35) );
  OAI21X1 U40 ( .A(n26), .B(n20), .C(n37), .Y(n65) );
  NAND2X1 U41 ( .A(N32), .B(n36), .Y(n37) );
  OAI21X1 U42 ( .A(n25), .B(n20), .C(n38), .Y(n66) );
  NAND2X1 U43 ( .A(N31), .B(n36), .Y(n38) );
  OAI21X1 U44 ( .A(n20), .B(n24), .C(n39), .Y(n67) );
  NAND2X1 U45 ( .A(N30), .B(n36), .Y(n39) );
  OAI21X1 U46 ( .A(n23), .B(n20), .C(n40), .Y(n68) );
  NAND2X1 U47 ( .A(N29), .B(n36), .Y(n40) );
  OAI21X1 U48 ( .A(n22), .B(n20), .C(n41), .Y(n69) );
  NAND2X1 U49 ( .A(N28), .B(n36), .Y(n41) );
  OAI21X1 U50 ( .A(n20), .B(n21), .C(n42), .Y(n70) );
  NAND2X1 U51 ( .A(N27), .B(n36), .Y(n42) );
  OAI21X1 U52 ( .A(n19), .B(n20), .C(n43), .Y(n71) );
  NAND2X1 U53 ( .A(N26), .B(n36), .Y(n43) );
  NOR2X1 U54 ( .A(n44), .B(n72), .Y(n36) );
  NOR2X1 U55 ( .A(n72), .B(TIMER_TRIG), .Y(n44) );
  NOR2X1 U56 ( .A(n45), .B(n46), .Y(n72) );
  NAND3X1 U57 ( .A(nextState[6]), .B(nextState[5]), .C(n47), .Y(n46) );
  NOR2X1 U58 ( .A(n22), .B(n23), .Y(n47) );
  NAND3X1 U59 ( .A(nextState[0]), .B(n21), .C(n48), .Y(n45) );
  NOR2X1 U60 ( .A(nextState[7]), .B(nextState[4]), .Y(n48) );
  NOR2X1 U61 ( .A(state[0]), .B(n49), .Y(N60) );
  AOI21X1 U62 ( .A(n51), .B(n32), .C(n52), .Y(n50) );
  OAI21X1 U63 ( .A(n33), .B(n53), .C(n54), .Y(n52) );
  NAND3X1 U64 ( .A(state[6]), .B(state[1]), .C(n55), .Y(n54) );
  AOI21X1 U65 ( .A(n56), .B(n57), .C(state[3]), .Y(n55) );
  NAND3X1 U66 ( .A(n33), .B(n31), .C(state[4]), .Y(n57) );
  NAND3X1 U67 ( .A(state[2]), .B(n32), .C(state[5]), .Y(n56) );
  NAND2X1 U68 ( .A(state[4]), .B(n58), .Y(n53) );
  OAI21X1 U69 ( .A(state[2]), .B(n28), .C(n59), .Y(n51) );
  NAND3X1 U70 ( .A(state[2]), .B(n29), .C(n30), .Y(n59) );
  OAI22X1 U71 ( .A(state[6]), .B(n61), .C(n29), .D(n60), .Y(n58) );
  NAND3X1 U72 ( .A(n34), .B(n31), .C(state[3]), .Y(n60) );
  AOI22X1 U73 ( .A(n62), .B(state[1]), .C(n63), .D(state[5]), .Y(n61) );
  XOR2X1 U74 ( .A(n34), .B(state[3]), .Y(n63) );
  NOR2X1 U75 ( .A(state[5]), .B(state[3]), .Y(n62) );
  uart_timer_1_DW01_inc_0 add_39 ( .A(nextState), .SUM({N33, N32, N31, N30, 
        N29, N28, N27, N26}) );
  DFFSR \nextState_reg[7]  ( .D(n64), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[7]) );
  INVX2 U19 ( .A(RST), .Y(n17) );
  INVX2 U22 ( .A(nextState[0]), .Y(n19) );
  INVX2 U23 ( .A(n44), .Y(n20) );
  INVX2 U24 ( .A(nextState[1]), .Y(n21) );
  INVX2 U25 ( .A(nextState[2]), .Y(n22) );
  INVX2 U26 ( .A(nextState[3]), .Y(n23) );
  INVX2 U27 ( .A(nextState[4]), .Y(n24) );
  INVX2 U28 ( .A(nextState[5]), .Y(n25) );
  INVX2 U29 ( .A(nextState[6]), .Y(n26) );
  INVX2 U30 ( .A(nextState[7]), .Y(n27) );
  INVX2 U31 ( .A(n58), .Y(n28) );
  INVX2 U32 ( .A(state[6]), .Y(n29) );
  INVX2 U33 ( .A(n60), .Y(n30) );
  INVX2 U34 ( .A(state[5]), .Y(n31) );
  INVX2 U35 ( .A(state[4]), .Y(n32) );
  INVX2 U36 ( .A(state[2]), .Y(n33) );
  INVX2 U37 ( .A(state[1]), .Y(n34) );
endmodule


module uart_rcv_block_1 ( CLK, RST, SERIAL_IN, KEY_ERROR, PROG_ERROR, PLAINKEY, 
        RBUF_FULL, PARITY_ERROR );
  output [63:0] PLAINKEY;
  input CLK, RST, SERIAL_IN;
  output KEY_ERROR, PROG_ERROR, RBUF_FULL, PARITY_ERROR;
  wire   START_BIT, CHK_ERROR, OE, SB_DETECT, STOP_RCVING, RBUF_LOAD, SBC_CLR,
         SBC_EN, SET_RBUF_FULL, TIMER_TRIG, CLR_RBUF, SBE, SHIFT_STROBE, n1,
         n2;
  wire   [7:0] LOAD_DATA;
  wire   [7:0] RCV_DATA;
  wire   [1:0] STOP_DATA;

  uart_edge_detector_1 U_0 ( .CLK(CLK), .RST(n1), .SERIAL_IN(SERIAL_IN), 
        .START_BIT(START_BIT) );
  uart_error_1 U_1 ( .RST(n1), .CLK(CLK), .RBUF_FULL(RBUF_FULL), .CHK_ERROR(
        CHK_ERROR), .OE(OE) );
  uart_rcu_1 U_2 ( .CLK(CLK), .RST(n1), .START_BIT(START_BIT), .STOP_RCVING(
        STOP_RCVING), .SB_DETECT(SB_DETECT), .RBUF_LOAD(RBUF_LOAD), 
        .TIMER_TRIG(TIMER_TRIG), .CHK_ERROR(CHK_ERROR), .SET_RBUF_FULL(
        SET_RBUF_FULL), .SBC_EN(SBC_EN), .SBC_CLR(SBC_CLR) );
  uart_rcv_buf_1 U_3 ( .CLK(CLK), .RST(n1), .LOAD_RBUF(RBUF_LOAD), .LOAD_DATA(
        LOAD_DATA), .RCV_DATA(RCV_DATA) );
  uart_rcv_buf_full_1 U_4 ( .CLK(CLK), .RST(n1), .CLR_RBUF(CLR_RBUF), 
        .SET_RBUF_FULL(SET_RBUF_FULL), .RBUF_FULL(RBUF_FULL) );
  uart_sb_check_1 U_5 ( .RST(n1), .CLK(CLK), .SBC_CLR(SBC_CLR), .SBC_EN(SBC_EN), .STOP_DATA(STOP_DATA), .SB_DETECT(SB_DETECT), .SBE(SBE) );
  uart_sr_10bit_1 U_6 ( .CLK(CLK), .RST(n1), .SHIFT_STROBE(SHIFT_STROBE), 
        .SERIAL_IN(SERIAL_IN), .LOAD_DATA(LOAD_DATA), .STOP_DATA(STOP_DATA) );
  keyreg_1 U_8 ( .CLK(CLK), .RST(n1), .SBE(SBE), .OE(OE), .RBUF_FULL(RBUF_FULL), .RCV_DATA(RCV_DATA), .PLAINKEY(PLAINKEY), .KEY_ERROR(KEY_ERROR), 
        .PROG_ERROR(PROG_ERROR), .CLR_RBUFF(CLR_RBUF), .PARITY_ERROR(
        PARITY_ERROR) );
  uart_timer_1 U_7 ( .CLK(CLK), .RST(n1), .TIMER_TRIG(TIMER_TRIG), 
        .STOP_RCVING(STOP_RCVING), .SHIFT_STROBE(SHIFT_STROBE) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module EDBlock_1 ( BYTE, BYTE_READY, CLK, OPCODE, RST, SERIAL_IN, DATA_IN, 
        KEY_ERROR, PARITY_ERROR, PDATA_READY, PROCESSED_DATA, PROG_ERROR, 
        RBUF_FULL, W_ENABLE, R_ENABLE, DATA, ADDR );
  input [7:0] BYTE;
  input [1:0] OPCODE;
  input [7:0] DATA_IN;
  output [7:0] PROCESSED_DATA;
  output [7:0] DATA;
  output [7:0] ADDR;
  input BYTE_READY, CLK, RST, SERIAL_IN;
  output KEY_ERROR, PARITY_ERROR, PDATA_READY, PROG_ERROR, RBUF_FULL, W_ENABLE,
         R_ENABLE;

  wire   [63:0] PLAINKEY;

  KSA_1 U_0 ( .KEY(PLAINKEY), .CLK(CLK), .RST(RST), .KEY_ERROR(KEY_ERROR), 
        .BYTE_READY(BYTE_READY), .BYTE(BYTE), .OPCODE(OPCODE), .DATA_IN(
        DATA_IN), .PROCESSED_DATA(PROCESSED_DATA), .PDATA_READY(PDATA_READY), 
        .W_ENABLE(W_ENABLE), .R_ENABLE(R_ENABLE), .ADDR(ADDR), .DATA(DATA) );
  uart_rcv_block_1 U_1 ( .CLK(CLK), .RST(RST), .SERIAL_IN(SERIAL_IN), 
        .KEY_ERROR(KEY_ERROR), .PROG_ERROR(PROG_ERROR), .PLAINKEY(PLAINKEY), 
        .RBUF_FULL(RBUF_FULL), .PARITY_ERROR(PARITY_ERROR) );
endmodule


module RBUFFER_1 ( CLK, RST, NEXT_BYTE, DATA, OPCODE, BYTE_COUNT, EOP, B_READY, 
        R_ENABLE, PRGA_IN, PRGA_OPCODE );
  input [7:0] DATA;
  input [1:0] OPCODE;
  input [4:0] BYTE_COUNT;
  output [7:0] PRGA_IN;
  output [1:0] PRGA_OPCODE;
  input CLK, RST, NEXT_BYTE, EOP;
  output B_READY, R_ENABLE;
  wire   N39, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n97, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n86, n88;
  wire   [2:0] state;
  wire   [2:0] nextState;
  wire   [7:0] tempData;
  wire   [1:0] tempOpcode;
  assign N39 = BYTE_COUNT[4];

  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n1), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n1), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n1), .S(1'b1), .Q(
        state[1]) );
  DFFPOSX1 B_READY_reg ( .D(n97), .CLK(CLK), .Q(B_READY) );
  DFFPOSX1 \tempData_reg[7]  ( .D(n68), .CLK(CLK), .Q(tempData[7]) );
  DFFPOSX1 \tempData_reg[6]  ( .D(n69), .CLK(CLK), .Q(tempData[6]) );
  DFFPOSX1 \tempData_reg[5]  ( .D(n70), .CLK(CLK), .Q(tempData[5]) );
  DFFPOSX1 \tempData_reg[4]  ( .D(n71), .CLK(CLK), .Q(tempData[4]) );
  DFFPOSX1 \tempData_reg[3]  ( .D(n72), .CLK(CLK), .Q(tempData[3]) );
  DFFPOSX1 \tempData_reg[2]  ( .D(n73), .CLK(CLK), .Q(tempData[2]) );
  DFFPOSX1 \tempData_reg[1]  ( .D(n74), .CLK(CLK), .Q(tempData[1]) );
  DFFPOSX1 \tempData_reg[0]  ( .D(n75), .CLK(CLK), .Q(tempData[0]) );
  DFFPOSX1 \tempOpcode_reg[1]  ( .D(n86), .CLK(CLK), .Q(tempOpcode[1]) );
  DFFPOSX1 \PRGA_OPCODE_reg[1]  ( .D(n87), .CLK(CLK), .Q(PRGA_OPCODE[1]) );
  DFFPOSX1 \tempOpcode_reg[0]  ( .D(n88), .CLK(CLK), .Q(tempOpcode[0]) );
  DFFPOSX1 \PRGA_OPCODE_reg[0]  ( .D(n85), .CLK(CLK), .Q(PRGA_OPCODE[0]) );
  DFFPOSX1 R_ENABLE_reg ( .D(n84), .CLK(CLK), .Q(R_ENABLE) );
  DFFPOSX1 \PRGA_IN_reg[7]  ( .D(n83), .CLK(CLK), .Q(PRGA_IN[7]) );
  DFFPOSX1 \PRGA_IN_reg[6]  ( .D(n82), .CLK(CLK), .Q(PRGA_IN[6]) );
  DFFPOSX1 \PRGA_IN_reg[5]  ( .D(n81), .CLK(CLK), .Q(PRGA_IN[5]) );
  DFFPOSX1 \PRGA_IN_reg[4]  ( .D(n80), .CLK(CLK), .Q(PRGA_IN[4]) );
  DFFPOSX1 \PRGA_IN_reg[3]  ( .D(n79), .CLK(CLK), .Q(PRGA_IN[3]) );
  DFFPOSX1 \PRGA_IN_reg[2]  ( .D(n78), .CLK(CLK), .Q(PRGA_IN[2]) );
  DFFPOSX1 \PRGA_IN_reg[1]  ( .D(n77), .CLK(CLK), .Q(PRGA_IN[1]) );
  DFFPOSX1 \PRGA_IN_reg[0]  ( .D(n76), .CLK(CLK), .Q(PRGA_IN[0]) );
  INVX2 U3 ( .A(n41), .Y(n28) );
  INVX2 U4 ( .A(RST), .Y(n1) );
  OR2X2 U5 ( .A(n39), .B(RST), .Y(n29) );
  AND2X2 U6 ( .A(n39), .B(n1), .Y(n44) );
  OAI21X1 U7 ( .A(n2), .B(n3), .C(n4), .Y(nextState[2]) );
  MUX2X1 U8 ( .B(n5), .A(n6), .S(state[0]), .Y(n4) );
  NOR2X1 U9 ( .A(state[2]), .B(n7), .Y(n6) );
  AND2X1 U10 ( .A(state[2]), .B(n8), .Y(n5) );
  OAI21X1 U11 ( .A(NEXT_BYTE), .B(n9), .C(state[1]), .Y(n8) );
  AND2X1 U12 ( .A(n10), .B(NEXT_BYTE), .Y(n2) );
  OAI21X1 U13 ( .A(state[2]), .B(n11), .C(n12), .Y(nextState[1]) );
  OAI21X1 U14 ( .A(n13), .B(n14), .C(n15), .Y(n12) );
  INVX1 U15 ( .A(n3), .Y(n14) );
  OAI21X1 U16 ( .A(state[2]), .B(n16), .C(n17), .Y(nextState[0]) );
  AOI22X1 U17 ( .A(n18), .B(n19), .C(NEXT_BYTE), .D(n20), .Y(n17) );
  OAI21X1 U18 ( .A(n10), .B(n3), .C(n21), .Y(n20) );
  INVX1 U19 ( .A(n13), .Y(n21) );
  NOR2X1 U20 ( .A(n16), .B(n9), .Y(n13) );
  NOR2X1 U21 ( .A(n22), .B(N39), .Y(n9) );
  NAND3X1 U22 ( .A(state[0]), .B(n7), .C(state[2]), .Y(n3) );
  AND2X1 U23 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n10) );
  OAI21X1 U24 ( .A(n23), .B(n15), .C(n24), .Y(n19) );
  INVX1 U25 ( .A(NEXT_BYTE), .Y(n15) );
  AOI21X1 U26 ( .A(EOP), .B(n22), .C(N39), .Y(n23) );
  NAND2X1 U27 ( .A(n25), .B(n26), .Y(n22) );
  NOR2X1 U28 ( .A(BYTE_COUNT[3]), .B(BYTE_COUNT[2]), .Y(n26) );
  NOR2X1 U29 ( .A(BYTE_COUNT[1]), .B(BYTE_COUNT[0]), .Y(n25) );
  NOR2X1 U30 ( .A(state[1]), .B(state[0]), .Y(n18) );
  INVX1 U31 ( .A(n27), .Y(n68) );
  AOI22X1 U32 ( .A(n28), .B(DATA[7]), .C(n29), .D(tempData[7]), .Y(n27) );
  INVX1 U33 ( .A(n30), .Y(n69) );
  AOI22X1 U34 ( .A(n28), .B(DATA[6]), .C(n29), .D(tempData[6]), .Y(n30) );
  INVX1 U35 ( .A(n31), .Y(n70) );
  AOI22X1 U36 ( .A(n28), .B(DATA[5]), .C(n29), .D(tempData[5]), .Y(n31) );
  INVX1 U37 ( .A(n32), .Y(n71) );
  AOI22X1 U38 ( .A(n28), .B(DATA[4]), .C(n29), .D(tempData[4]), .Y(n32) );
  INVX1 U39 ( .A(n33), .Y(n72) );
  AOI22X1 U40 ( .A(n28), .B(DATA[3]), .C(n29), .D(tempData[3]), .Y(n33) );
  INVX1 U41 ( .A(n34), .Y(n73) );
  AOI22X1 U42 ( .A(n28), .B(DATA[2]), .C(n29), .D(tempData[2]), .Y(n34) );
  INVX1 U43 ( .A(n35), .Y(n74) );
  AOI22X1 U44 ( .A(n28), .B(DATA[1]), .C(n29), .D(tempData[1]), .Y(n35) );
  INVX1 U45 ( .A(n36), .Y(n75) );
  AOI22X1 U46 ( .A(n28), .B(DATA[0]), .C(n29), .D(tempData[0]), .Y(n36) );
  INVX1 U47 ( .A(n37), .Y(n86) );
  AOI22X1 U48 ( .A(OPCODE[1]), .B(n28), .C(n29), .D(tempOpcode[1]), .Y(n37) );
  INVX1 U49 ( .A(n38), .Y(n88) );
  AOI22X1 U50 ( .A(OPCODE[0]), .B(n28), .C(n29), .D(tempOpcode[0]), .Y(n38) );
  OAI21X1 U51 ( .A(n1), .B(n40), .C(n41), .Y(n97) );
  INVX1 U52 ( .A(B_READY), .Y(n40) );
  OAI21X1 U53 ( .A(n1), .B(n42), .C(n43), .Y(n87) );
  AOI22X1 U54 ( .A(n28), .B(OPCODE[1]), .C(n44), .D(tempOpcode[1]), .Y(n43) );
  INVX1 U55 ( .A(PRGA_OPCODE[1]), .Y(n42) );
  OAI21X1 U56 ( .A(n1), .B(n45), .C(n46), .Y(n85) );
  AOI22X1 U57 ( .A(n28), .B(OPCODE[0]), .C(n44), .D(tempOpcode[0]), .Y(n46) );
  INVX1 U58 ( .A(PRGA_OPCODE[0]), .Y(n45) );
  MUX2X1 U59 ( .B(n47), .A(n48), .S(RST), .Y(n84) );
  INVX1 U60 ( .A(R_ENABLE), .Y(n48) );
  NAND3X1 U61 ( .A(n7), .B(n24), .C(state[0]), .Y(n47) );
  OAI21X1 U62 ( .A(n1), .B(n49), .C(n50), .Y(n83) );
  AOI22X1 U63 ( .A(DATA[7]), .B(n28), .C(n44), .D(tempData[7]), .Y(n50) );
  INVX1 U64 ( .A(PRGA_IN[7]), .Y(n49) );
  OAI21X1 U65 ( .A(n1), .B(n51), .C(n52), .Y(n82) );
  AOI22X1 U66 ( .A(DATA[6]), .B(n28), .C(n44), .D(tempData[6]), .Y(n52) );
  INVX1 U67 ( .A(PRGA_IN[6]), .Y(n51) );
  OAI21X1 U68 ( .A(n1), .B(n53), .C(n54), .Y(n81) );
  AOI22X1 U69 ( .A(DATA[5]), .B(n28), .C(n44), .D(tempData[5]), .Y(n54) );
  INVX1 U70 ( .A(PRGA_IN[5]), .Y(n53) );
  OAI21X1 U71 ( .A(n1), .B(n55), .C(n56), .Y(n80) );
  AOI22X1 U72 ( .A(DATA[4]), .B(n28), .C(n44), .D(tempData[4]), .Y(n56) );
  INVX1 U73 ( .A(PRGA_IN[4]), .Y(n55) );
  OAI21X1 U74 ( .A(n1), .B(n57), .C(n58), .Y(n79) );
  AOI22X1 U75 ( .A(DATA[3]), .B(n28), .C(n44), .D(tempData[3]), .Y(n58) );
  INVX1 U76 ( .A(PRGA_IN[3]), .Y(n57) );
  OAI21X1 U77 ( .A(n1), .B(n59), .C(n60), .Y(n78) );
  AOI22X1 U78 ( .A(DATA[2]), .B(n28), .C(n44), .D(tempData[2]), .Y(n60) );
  INVX1 U79 ( .A(PRGA_IN[2]), .Y(n59) );
  OAI21X1 U80 ( .A(n1), .B(n61), .C(n62), .Y(n77) );
  AOI22X1 U81 ( .A(DATA[1]), .B(n28), .C(n44), .D(tempData[1]), .Y(n62) );
  INVX1 U82 ( .A(PRGA_IN[1]), .Y(n61) );
  OAI21X1 U83 ( .A(n1), .B(n63), .C(n64), .Y(n76) );
  AOI22X1 U84 ( .A(DATA[0]), .B(n28), .C(n44), .D(tempData[0]), .Y(n64) );
  NAND2X1 U85 ( .A(n11), .B(state[2]), .Y(n39) );
  INVX1 U86 ( .A(n65), .Y(n11) );
  OAI21X1 U87 ( .A(state[1]), .B(n66), .C(n16), .Y(n65) );
  NAND2X1 U88 ( .A(state[1]), .B(n66), .Y(n16) );
  NAND3X1 U89 ( .A(n66), .B(n7), .C(n67), .Y(n41) );
  NOR2X1 U90 ( .A(RST), .B(n24), .Y(n67) );
  INVX1 U91 ( .A(state[2]), .Y(n24) );
  INVX1 U92 ( .A(state[1]), .Y(n7) );
  INVX1 U93 ( .A(state[0]), .Y(n66) );
  INVX1 U94 ( .A(PRGA_IN[0]), .Y(n63) );
endmodule


module RFIFO_1 ( CLK, RST, W_ENABLE, R_ENABLE, RCV_DATA, RCV_OPCODE, DATA, 
        OUT_OPCODE, BYTE_COUNT, EMPTY, FULL );
  input [7:0] RCV_DATA;
  input [1:0] RCV_OPCODE;
  output [7:0] DATA;
  output [1:0] OUT_OPCODE;
  output [4:0] BYTE_COUNT;
  input CLK, RST, W_ENABLE, R_ENABLE;
  output EMPTY, FULL;
  wire   state, \opcode[0][1] , \opcode[0][0] , \opcode[1][1] , \opcode[1][0] ,
         \opcode[2][1] , \opcode[2][0] , \opcode[3][1] , \opcode[3][0] ,
         \opcode[4][1] , \opcode[4][0] , \opcode[5][1] , \opcode[5][0] ,
         \opcode[6][1] , \opcode[6][0] , \opcode[7][1] , \opcode[7][0] ,
         \opcode[8][1] , \opcode[8][0] , \opcode[9][1] , \opcode[9][0] ,
         \opcode[10][1] , \opcode[10][0] , \opcode[11][1] , \opcode[11][0] ,
         \opcode[12][1] , \opcode[12][0] , \opcode[13][1] , \opcode[13][0] ,
         \opcode[14][1] , \opcode[14][0] , \opcode[15][1] , \opcode[15][0] ,
         \opcode[16][1] , \opcode[16][0] , \opcode[17][1] , \opcode[17][0] ,
         \opcode[18][1] , \opcode[18][0] , \opcode[19][1] , \opcode[19][0] ,
         \opcode[20][1] , \opcode[20][0] , \opcode[21][1] , \opcode[21][0] ,
         \opcode[22][1] , \opcode[22][0] , \opcode[23][1] , \opcode[23][0] ,
         \opcode[24][1] , \opcode[24][0] , \opcode[25][1] , \opcode[25][0] ,
         \opcode[26][1] , \opcode[26][0] , \opcode[27][1] , \opcode[27][0] ,
         \opcode[28][1] , \opcode[28][0] , \opcode[29][1] , \opcode[29][0] ,
         \opcode[30][1] , \opcode[30][0] , \opcode[31][1] , \opcode[31][0] ,
         \memory[0][7] , \memory[0][6] , \memory[0][5] , \memory[0][4] ,
         \memory[0][3] , \memory[0][2] , \memory[0][1] , \memory[0][0] ,
         \memory[1][7] , \memory[1][6] , \memory[1][5] , \memory[1][4] ,
         \memory[1][3] , \memory[1][2] , \memory[1][1] , \memory[1][0] ,
         \memory[2][7] , \memory[2][6] , \memory[2][5] , \memory[2][4] ,
         \memory[2][3] , \memory[2][2] , \memory[2][1] , \memory[2][0] ,
         \memory[3][7] , \memory[3][6] , \memory[3][5] , \memory[3][4] ,
         \memory[3][3] , \memory[3][2] , \memory[3][1] , \memory[3][0] ,
         \memory[4][7] , \memory[4][6] , \memory[4][5] , \memory[4][4] ,
         \memory[4][3] , \memory[4][2] , \memory[4][1] , \memory[4][0] ,
         \memory[5][7] , \memory[5][6] , \memory[5][5] , \memory[5][4] ,
         \memory[5][3] , \memory[5][2] , \memory[5][1] , \memory[5][0] ,
         \memory[6][7] , \memory[6][6] , \memory[6][5] , \memory[6][4] ,
         \memory[6][3] , \memory[6][2] , \memory[6][1] , \memory[6][0] ,
         \memory[7][7] , \memory[7][6] , \memory[7][5] , \memory[7][4] ,
         \memory[7][3] , \memory[7][2] , \memory[7][1] , \memory[7][0] ,
         \memory[8][7] , \memory[8][6] , \memory[8][5] , \memory[8][4] ,
         \memory[8][3] , \memory[8][2] , \memory[8][1] , \memory[8][0] ,
         \memory[9][7] , \memory[9][6] , \memory[9][5] , \memory[9][4] ,
         \memory[9][3] , \memory[9][2] , \memory[9][1] , \memory[9][0] ,
         \memory[10][7] , \memory[10][6] , \memory[10][5] , \memory[10][4] ,
         \memory[10][3] , \memory[10][2] , \memory[10][1] , \memory[10][0] ,
         \memory[11][7] , \memory[11][6] , \memory[11][5] , \memory[11][4] ,
         \memory[11][3] , \memory[11][2] , \memory[11][1] , \memory[11][0] ,
         \memory[12][7] , \memory[12][6] , \memory[12][5] , \memory[12][4] ,
         \memory[12][3] , \memory[12][2] , \memory[12][1] , \memory[12][0] ,
         \memory[13][7] , \memory[13][6] , \memory[13][5] , \memory[13][4] ,
         \memory[13][3] , \memory[13][2] , \memory[13][1] , \memory[13][0] ,
         \memory[14][7] , \memory[14][6] , \memory[14][5] , \memory[14][4] ,
         \memory[14][3] , \memory[14][2] , \memory[14][1] , \memory[14][0] ,
         \memory[15][7] , \memory[15][6] , \memory[15][5] , \memory[15][4] ,
         \memory[15][3] , \memory[15][2] , \memory[15][1] , \memory[15][0] ,
         \memory[16][7] , \memory[16][6] , \memory[16][5] , \memory[16][4] ,
         \memory[16][3] , \memory[16][2] , \memory[16][1] , \memory[16][0] ,
         \memory[17][7] , \memory[17][6] , \memory[17][5] , \memory[17][4] ,
         \memory[17][3] , \memory[17][2] , \memory[17][1] , \memory[17][0] ,
         \memory[18][7] , \memory[18][6] , \memory[18][5] , \memory[18][4] ,
         \memory[18][3] , \memory[18][2] , \memory[18][1] , \memory[18][0] ,
         \memory[19][7] , \memory[19][6] , \memory[19][5] , \memory[19][4] ,
         \memory[19][3] , \memory[19][2] , \memory[19][1] , \memory[19][0] ,
         \memory[20][7] , \memory[20][6] , \memory[20][5] , \memory[20][4] ,
         \memory[20][3] , \memory[20][2] , \memory[20][1] , \memory[20][0] ,
         \memory[21][7] , \memory[21][6] , \memory[21][5] , \memory[21][4] ,
         \memory[21][3] , \memory[21][2] , \memory[21][1] , \memory[21][0] ,
         \memory[22][7] , \memory[22][6] , \memory[22][5] , \memory[22][4] ,
         \memory[22][3] , \memory[22][2] , \memory[22][1] , \memory[22][0] ,
         \memory[23][7] , \memory[23][6] , \memory[23][5] , \memory[23][4] ,
         \memory[23][3] , \memory[23][2] , \memory[23][1] , \memory[23][0] ,
         \memory[24][7] , \memory[24][6] , \memory[24][5] , \memory[24][4] ,
         \memory[24][3] , \memory[24][2] , \memory[24][1] , \memory[24][0] ,
         \memory[25][7] , \memory[25][6] , \memory[25][5] , \memory[25][4] ,
         \memory[25][3] , \memory[25][2] , \memory[25][1] , \memory[25][0] ,
         \memory[26][7] , \memory[26][6] , \memory[26][5] , \memory[26][4] ,
         \memory[26][3] , \memory[26][2] , \memory[26][1] , \memory[26][0] ,
         \memory[27][7] , \memory[27][6] , \memory[27][5] , \memory[27][4] ,
         \memory[27][3] , \memory[27][2] , \memory[27][1] , \memory[27][0] ,
         \memory[28][7] , \memory[28][6] , \memory[28][5] , \memory[28][4] ,
         \memory[28][3] , \memory[28][2] , \memory[28][1] , \memory[28][0] ,
         \memory[29][7] , \memory[29][6] , \memory[29][5] , \memory[29][4] ,
         \memory[29][3] , \memory[29][2] , \memory[29][1] , \memory[29][0] ,
         \memory[30][7] , \memory[30][6] , \memory[30][5] , \memory[30][4] ,
         \memory[30][3] , \memory[30][2] , \memory[30][1] , \memory[30][0] ,
         \memory[31][7] , \memory[31][6] , \memory[31][5] , \memory[31][4] ,
         \memory[31][3] , \memory[31][2] , \memory[31][1] , \memory[31][0] ,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, n854,
         n856, n858, n860, n862, n869, n870, n871, n872, n873, n874, n875,
         n876, n879, n880, n881, n882, n883, n884, n885, n886, n889, n890,
         n891, n892, n893, n894, n895, n896, n899, n900, n901, n902, n903,
         n904, n905, n906, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1056, n1057, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n852,
         n865, n877, n878, n887, n888, n897, n898, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415;
  wire   [4:0] readptr;
  wire   [4:0] writeptr;

  DFFSR state_reg ( .D(1'b1), .CLK(CLK), .R(n177), .S(1'b1), .Q(state) );
  DFFSR \readptr_reg[0]  ( .D(N343), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        readptr[0]) );
  DFFSR \readptr_reg[1]  ( .D(N344), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        readptr[1]) );
  DFFSR \readptr_reg[3]  ( .D(N346), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        readptr[3]) );
  DFFSR \readptr_reg[4]  ( .D(N347), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        readptr[4]) );
  DFFSR \writeptr_reg[4]  ( .D(n862), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        writeptr[4]) );
  DFFSR \writeptr_reg[3]  ( .D(n860), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        writeptr[3]) );
  DFFSR \writeptr_reg[0]  ( .D(n858), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        writeptr[0]) );
  DFFSR \writeptr_reg[1]  ( .D(n856), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        writeptr[1]) );
  DFFSR \writeptr_reg[2]  ( .D(n854), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        writeptr[2]) );
  DFFPOSX1 FULL_reg ( .D(n1414), .CLK(CLK), .Q(FULL) );
  DFFSR \BYTE_COUNT_reg[4]  ( .D(N342), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        BYTE_COUNT[4]) );
  DFFSR \BYTE_COUNT_reg[3]  ( .D(N341), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        BYTE_COUNT[3]) );
  DFFSR \BYTE_COUNT_reg[2]  ( .D(N340), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        BYTE_COUNT[2]) );
  DFFSR \BYTE_COUNT_reg[1]  ( .D(N339), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        BYTE_COUNT[1]) );
  DFFSR \BYTE_COUNT_reg[0]  ( .D(N338), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        BYTE_COUNT[0]) );
  DFFPOSX1 \memory_reg[0][7]  ( .D(n1389), .CLK(CLK), .Q(\memory[0][7] ) );
  DFFPOSX1 \memory_reg[0][6]  ( .D(n1388), .CLK(CLK), .Q(\memory[0][6] ) );
  DFFPOSX1 \memory_reg[0][5]  ( .D(n1387), .CLK(CLK), .Q(\memory[0][5] ) );
  DFFPOSX1 \memory_reg[0][4]  ( .D(n1386), .CLK(CLK), .Q(\memory[0][4] ) );
  DFFPOSX1 \memory_reg[0][3]  ( .D(n1385), .CLK(CLK), .Q(\memory[0][3] ) );
  DFFPOSX1 \memory_reg[0][2]  ( .D(n1384), .CLK(CLK), .Q(\memory[0][2] ) );
  DFFPOSX1 \memory_reg[0][1]  ( .D(n1383), .CLK(CLK), .Q(\memory[0][1] ) );
  DFFPOSX1 \memory_reg[0][0]  ( .D(n1382), .CLK(CLK), .Q(\memory[0][0] ) );
  DFFPOSX1 \memory_reg[1][7]  ( .D(n1397), .CLK(CLK), .Q(\memory[1][7] ) );
  DFFPOSX1 \memory_reg[1][6]  ( .D(n1396), .CLK(CLK), .Q(\memory[1][6] ) );
  DFFPOSX1 \memory_reg[1][5]  ( .D(n1395), .CLK(CLK), .Q(\memory[1][5] ) );
  DFFPOSX1 \memory_reg[1][4]  ( .D(n1394), .CLK(CLK), .Q(\memory[1][4] ) );
  DFFPOSX1 \memory_reg[1][3]  ( .D(n1393), .CLK(CLK), .Q(\memory[1][3] ) );
  DFFPOSX1 \memory_reg[1][2]  ( .D(n1392), .CLK(CLK), .Q(\memory[1][2] ) );
  DFFPOSX1 \memory_reg[1][1]  ( .D(n1391), .CLK(CLK), .Q(\memory[1][1] ) );
  DFFPOSX1 \memory_reg[1][0]  ( .D(n1390), .CLK(CLK), .Q(\memory[1][0] ) );
  DFFPOSX1 \memory_reg[2][7]  ( .D(n1405), .CLK(CLK), .Q(\memory[2][7] ) );
  DFFPOSX1 \memory_reg[2][6]  ( .D(n1404), .CLK(CLK), .Q(\memory[2][6] ) );
  DFFPOSX1 \memory_reg[2][5]  ( .D(n1403), .CLK(CLK), .Q(\memory[2][5] ) );
  DFFPOSX1 \memory_reg[2][4]  ( .D(n1402), .CLK(CLK), .Q(\memory[2][4] ) );
  DFFPOSX1 \memory_reg[2][3]  ( .D(n1401), .CLK(CLK), .Q(\memory[2][3] ) );
  DFFPOSX1 \memory_reg[2][2]  ( .D(n1400), .CLK(CLK), .Q(\memory[2][2] ) );
  DFFPOSX1 \memory_reg[2][1]  ( .D(n1399), .CLK(CLK), .Q(\memory[2][1] ) );
  DFFPOSX1 \memory_reg[2][0]  ( .D(n1398), .CLK(CLK), .Q(\memory[2][0] ) );
  DFFPOSX1 \memory_reg[3][7]  ( .D(n1413), .CLK(CLK), .Q(\memory[3][7] ) );
  DFFPOSX1 \memory_reg[3][6]  ( .D(n1412), .CLK(CLK), .Q(\memory[3][6] ) );
  DFFPOSX1 \memory_reg[3][5]  ( .D(n1411), .CLK(CLK), .Q(\memory[3][5] ) );
  DFFPOSX1 \memory_reg[3][4]  ( .D(n1410), .CLK(CLK), .Q(\memory[3][4] ) );
  DFFPOSX1 \memory_reg[3][3]  ( .D(n1409), .CLK(CLK), .Q(\memory[3][3] ) );
  DFFPOSX1 \memory_reg[3][2]  ( .D(n1408), .CLK(CLK), .Q(\memory[3][2] ) );
  DFFPOSX1 \memory_reg[3][1]  ( .D(n1407), .CLK(CLK), .Q(\memory[3][1] ) );
  DFFPOSX1 \memory_reg[3][0]  ( .D(n1406), .CLK(CLK), .Q(\memory[3][0] ) );
  DFFPOSX1 \memory_reg[4][7]  ( .D(n869), .CLK(CLK), .Q(\memory[4][7] ) );
  DFFPOSX1 \memory_reg[4][6]  ( .D(n870), .CLK(CLK), .Q(\memory[4][6] ) );
  DFFPOSX1 \memory_reg[4][5]  ( .D(n871), .CLK(CLK), .Q(\memory[4][5] ) );
  DFFPOSX1 \memory_reg[4][4]  ( .D(n872), .CLK(CLK), .Q(\memory[4][4] ) );
  DFFPOSX1 \memory_reg[4][3]  ( .D(n873), .CLK(CLK), .Q(\memory[4][3] ) );
  DFFPOSX1 \memory_reg[4][2]  ( .D(n874), .CLK(CLK), .Q(\memory[4][2] ) );
  DFFPOSX1 \memory_reg[4][1]  ( .D(n875), .CLK(CLK), .Q(\memory[4][1] ) );
  DFFPOSX1 \memory_reg[4][0]  ( .D(n876), .CLK(CLK), .Q(\memory[4][0] ) );
  DFFPOSX1 \memory_reg[5][7]  ( .D(n879), .CLK(CLK), .Q(\memory[5][7] ) );
  DFFPOSX1 \memory_reg[5][6]  ( .D(n880), .CLK(CLK), .Q(\memory[5][6] ) );
  DFFPOSX1 \memory_reg[5][5]  ( .D(n881), .CLK(CLK), .Q(\memory[5][5] ) );
  DFFPOSX1 \memory_reg[5][4]  ( .D(n882), .CLK(CLK), .Q(\memory[5][4] ) );
  DFFPOSX1 \memory_reg[5][3]  ( .D(n883), .CLK(CLK), .Q(\memory[5][3] ) );
  DFFPOSX1 \memory_reg[5][2]  ( .D(n884), .CLK(CLK), .Q(\memory[5][2] ) );
  DFFPOSX1 \memory_reg[5][1]  ( .D(n885), .CLK(CLK), .Q(\memory[5][1] ) );
  DFFPOSX1 \memory_reg[5][0]  ( .D(n886), .CLK(CLK), .Q(\memory[5][0] ) );
  DFFPOSX1 \memory_reg[6][7]  ( .D(n889), .CLK(CLK), .Q(\memory[6][7] ) );
  DFFPOSX1 \memory_reg[6][6]  ( .D(n890), .CLK(CLK), .Q(\memory[6][6] ) );
  DFFPOSX1 \memory_reg[6][5]  ( .D(n891), .CLK(CLK), .Q(\memory[6][5] ) );
  DFFPOSX1 \memory_reg[6][4]  ( .D(n892), .CLK(CLK), .Q(\memory[6][4] ) );
  DFFPOSX1 \memory_reg[6][3]  ( .D(n893), .CLK(CLK), .Q(\memory[6][3] ) );
  DFFPOSX1 \memory_reg[6][2]  ( .D(n894), .CLK(CLK), .Q(\memory[6][2] ) );
  DFFPOSX1 \memory_reg[6][1]  ( .D(n895), .CLK(CLK), .Q(\memory[6][1] ) );
  DFFPOSX1 \memory_reg[6][0]  ( .D(n896), .CLK(CLK), .Q(\memory[6][0] ) );
  DFFPOSX1 \memory_reg[7][7]  ( .D(n899), .CLK(CLK), .Q(\memory[7][7] ) );
  DFFPOSX1 \memory_reg[7][6]  ( .D(n900), .CLK(CLK), .Q(\memory[7][6] ) );
  DFFPOSX1 \memory_reg[7][5]  ( .D(n901), .CLK(CLK), .Q(\memory[7][5] ) );
  DFFPOSX1 \memory_reg[7][4]  ( .D(n902), .CLK(CLK), .Q(\memory[7][4] ) );
  DFFPOSX1 \memory_reg[7][3]  ( .D(n903), .CLK(CLK), .Q(\memory[7][3] ) );
  DFFPOSX1 \memory_reg[7][2]  ( .D(n904), .CLK(CLK), .Q(\memory[7][2] ) );
  DFFPOSX1 \memory_reg[7][1]  ( .D(n905), .CLK(CLK), .Q(\memory[7][1] ) );
  DFFPOSX1 \memory_reg[7][0]  ( .D(n906), .CLK(CLK), .Q(\memory[7][0] ) );
  DFFPOSX1 \memory_reg[8][7]  ( .D(n1167), .CLK(CLK), .Q(\memory[8][7] ) );
  DFFPOSX1 \memory_reg[8][6]  ( .D(n1166), .CLK(CLK), .Q(\memory[8][6] ) );
  DFFPOSX1 \memory_reg[8][5]  ( .D(n1165), .CLK(CLK), .Q(\memory[8][5] ) );
  DFFPOSX1 \memory_reg[8][4]  ( .D(n1164), .CLK(CLK), .Q(\memory[8][4] ) );
  DFFPOSX1 \memory_reg[8][3]  ( .D(n1163), .CLK(CLK), .Q(\memory[8][3] ) );
  DFFPOSX1 \memory_reg[8][2]  ( .D(n1162), .CLK(CLK), .Q(\memory[8][2] ) );
  DFFPOSX1 \memory_reg[8][1]  ( .D(n1161), .CLK(CLK), .Q(\memory[8][1] ) );
  DFFPOSX1 \memory_reg[8][0]  ( .D(n1160), .CLK(CLK), .Q(\memory[8][0] ) );
  DFFPOSX1 \memory_reg[9][7]  ( .D(n1159), .CLK(CLK), .Q(\memory[9][7] ) );
  DFFPOSX1 \memory_reg[9][6]  ( .D(n1158), .CLK(CLK), .Q(\memory[9][6] ) );
  DFFPOSX1 \memory_reg[9][5]  ( .D(n1157), .CLK(CLK), .Q(\memory[9][5] ) );
  DFFPOSX1 \memory_reg[9][4]  ( .D(n1156), .CLK(CLK), .Q(\memory[9][4] ) );
  DFFPOSX1 \memory_reg[9][3]  ( .D(n1155), .CLK(CLK), .Q(\memory[9][3] ) );
  DFFPOSX1 \memory_reg[9][2]  ( .D(n1154), .CLK(CLK), .Q(\memory[9][2] ) );
  DFFPOSX1 \memory_reg[9][1]  ( .D(n1153), .CLK(CLK), .Q(\memory[9][1] ) );
  DFFPOSX1 \memory_reg[9][0]  ( .D(n1152), .CLK(CLK), .Q(\memory[9][0] ) );
  DFFPOSX1 \memory_reg[10][7]  ( .D(n1151), .CLK(CLK), .Q(\memory[10][7] ) );
  DFFPOSX1 \memory_reg[10][6]  ( .D(n1150), .CLK(CLK), .Q(\memory[10][6] ) );
  DFFPOSX1 \memory_reg[10][5]  ( .D(n1149), .CLK(CLK), .Q(\memory[10][5] ) );
  DFFPOSX1 \memory_reg[10][4]  ( .D(n1148), .CLK(CLK), .Q(\memory[10][4] ) );
  DFFPOSX1 \memory_reg[10][3]  ( .D(n1147), .CLK(CLK), .Q(\memory[10][3] ) );
  DFFPOSX1 \memory_reg[10][2]  ( .D(n1146), .CLK(CLK), .Q(\memory[10][2] ) );
  DFFPOSX1 \memory_reg[10][1]  ( .D(n1145), .CLK(CLK), .Q(\memory[10][1] ) );
  DFFPOSX1 \memory_reg[10][0]  ( .D(n1144), .CLK(CLK), .Q(\memory[10][0] ) );
  DFFPOSX1 \memory_reg[11][7]  ( .D(n1143), .CLK(CLK), .Q(\memory[11][7] ) );
  DFFPOSX1 \memory_reg[11][6]  ( .D(n1142), .CLK(CLK), .Q(\memory[11][6] ) );
  DFFPOSX1 \memory_reg[11][5]  ( .D(n1141), .CLK(CLK), .Q(\memory[11][5] ) );
  DFFPOSX1 \memory_reg[11][4]  ( .D(n1140), .CLK(CLK), .Q(\memory[11][4] ) );
  DFFPOSX1 \memory_reg[11][3]  ( .D(n1139), .CLK(CLK), .Q(\memory[11][3] ) );
  DFFPOSX1 \memory_reg[11][2]  ( .D(n1138), .CLK(CLK), .Q(\memory[11][2] ) );
  DFFPOSX1 \memory_reg[11][1]  ( .D(n1137), .CLK(CLK), .Q(\memory[11][1] ) );
  DFFPOSX1 \memory_reg[11][0]  ( .D(n1136), .CLK(CLK), .Q(\memory[11][0] ) );
  DFFPOSX1 \memory_reg[12][7]  ( .D(n1374), .CLK(CLK), .Q(\memory[12][7] ) );
  DFFPOSX1 \memory_reg[12][6]  ( .D(n1375), .CLK(CLK), .Q(\memory[12][6] ) );
  DFFPOSX1 \memory_reg[12][5]  ( .D(n1376), .CLK(CLK), .Q(\memory[12][5] ) );
  DFFPOSX1 \memory_reg[12][4]  ( .D(n1377), .CLK(CLK), .Q(\memory[12][4] ) );
  DFFPOSX1 \memory_reg[12][3]  ( .D(n1378), .CLK(CLK), .Q(\memory[12][3] ) );
  DFFPOSX1 \memory_reg[12][2]  ( .D(n1379), .CLK(CLK), .Q(\memory[12][2] ) );
  DFFPOSX1 \memory_reg[12][1]  ( .D(n1380), .CLK(CLK), .Q(\memory[12][1] ) );
  DFFPOSX1 \memory_reg[12][0]  ( .D(n1381), .CLK(CLK), .Q(\memory[12][0] ) );
  DFFPOSX1 \memory_reg[13][7]  ( .D(n1366), .CLK(CLK), .Q(\memory[13][7] ) );
  DFFPOSX1 \memory_reg[13][6]  ( .D(n1367), .CLK(CLK), .Q(\memory[13][6] ) );
  DFFPOSX1 \memory_reg[13][5]  ( .D(n1368), .CLK(CLK), .Q(\memory[13][5] ) );
  DFFPOSX1 \memory_reg[13][4]  ( .D(n1369), .CLK(CLK), .Q(\memory[13][4] ) );
  DFFPOSX1 \memory_reg[13][3]  ( .D(n1370), .CLK(CLK), .Q(\memory[13][3] ) );
  DFFPOSX1 \memory_reg[13][2]  ( .D(n1371), .CLK(CLK), .Q(\memory[13][2] ) );
  DFFPOSX1 \memory_reg[13][1]  ( .D(n1372), .CLK(CLK), .Q(\memory[13][1] ) );
  DFFPOSX1 \memory_reg[13][0]  ( .D(n1373), .CLK(CLK), .Q(\memory[13][0] ) );
  DFFPOSX1 \memory_reg[14][7]  ( .D(n1358), .CLK(CLK), .Q(\memory[14][7] ) );
  DFFPOSX1 \memory_reg[14][6]  ( .D(n1359), .CLK(CLK), .Q(\memory[14][6] ) );
  DFFPOSX1 \memory_reg[14][5]  ( .D(n1360), .CLK(CLK), .Q(\memory[14][5] ) );
  DFFPOSX1 \memory_reg[14][4]  ( .D(n1361), .CLK(CLK), .Q(\memory[14][4] ) );
  DFFPOSX1 \memory_reg[14][3]  ( .D(n1362), .CLK(CLK), .Q(\memory[14][3] ) );
  DFFPOSX1 \memory_reg[14][2]  ( .D(n1363), .CLK(CLK), .Q(\memory[14][2] ) );
  DFFPOSX1 \memory_reg[14][1]  ( .D(n1364), .CLK(CLK), .Q(\memory[14][1] ) );
  DFFPOSX1 \memory_reg[14][0]  ( .D(n1365), .CLK(CLK), .Q(\memory[14][0] ) );
  DFFPOSX1 \memory_reg[15][7]  ( .D(n1350), .CLK(CLK), .Q(\memory[15][7] ) );
  DFFPOSX1 \memory_reg[15][6]  ( .D(n1351), .CLK(CLK), .Q(\memory[15][6] ) );
  DFFPOSX1 \memory_reg[15][5]  ( .D(n1352), .CLK(CLK), .Q(\memory[15][5] ) );
  DFFPOSX1 \memory_reg[15][4]  ( .D(n1353), .CLK(CLK), .Q(\memory[15][4] ) );
  DFFPOSX1 \memory_reg[15][3]  ( .D(n1354), .CLK(CLK), .Q(\memory[15][3] ) );
  DFFPOSX1 \memory_reg[15][2]  ( .D(n1355), .CLK(CLK), .Q(\memory[15][2] ) );
  DFFPOSX1 \memory_reg[15][1]  ( .D(n1356), .CLK(CLK), .Q(\memory[15][1] ) );
  DFFPOSX1 \memory_reg[15][0]  ( .D(n1357), .CLK(CLK), .Q(\memory[15][0] ) );
  DFFPOSX1 \memory_reg[16][7]  ( .D(n1135), .CLK(CLK), .Q(\memory[16][7] ) );
  DFFPOSX1 \memory_reg[16][6]  ( .D(n1134), .CLK(CLK), .Q(\memory[16][6] ) );
  DFFPOSX1 \memory_reg[16][5]  ( .D(n1133), .CLK(CLK), .Q(\memory[16][5] ) );
  DFFPOSX1 \memory_reg[16][4]  ( .D(n1132), .CLK(CLK), .Q(\memory[16][4] ) );
  DFFPOSX1 \memory_reg[16][3]  ( .D(n1131), .CLK(CLK), .Q(\memory[16][3] ) );
  DFFPOSX1 \memory_reg[16][2]  ( .D(n1130), .CLK(CLK), .Q(\memory[16][2] ) );
  DFFPOSX1 \memory_reg[16][1]  ( .D(n1129), .CLK(CLK), .Q(\memory[16][1] ) );
  DFFPOSX1 \memory_reg[16][0]  ( .D(n1128), .CLK(CLK), .Q(\memory[16][0] ) );
  DFFPOSX1 \memory_reg[17][7]  ( .D(n1127), .CLK(CLK), .Q(\memory[17][7] ) );
  DFFPOSX1 \memory_reg[17][6]  ( .D(n1126), .CLK(CLK), .Q(\memory[17][6] ) );
  DFFPOSX1 \memory_reg[17][5]  ( .D(n1125), .CLK(CLK), .Q(\memory[17][5] ) );
  DFFPOSX1 \memory_reg[17][4]  ( .D(n1124), .CLK(CLK), .Q(\memory[17][4] ) );
  DFFPOSX1 \memory_reg[17][3]  ( .D(n1123), .CLK(CLK), .Q(\memory[17][3] ) );
  DFFPOSX1 \memory_reg[17][2]  ( .D(n1122), .CLK(CLK), .Q(\memory[17][2] ) );
  DFFPOSX1 \memory_reg[17][1]  ( .D(n1121), .CLK(CLK), .Q(\memory[17][1] ) );
  DFFPOSX1 \memory_reg[17][0]  ( .D(n1120), .CLK(CLK), .Q(\memory[17][0] ) );
  DFFPOSX1 \memory_reg[18][7]  ( .D(n1119), .CLK(CLK), .Q(\memory[18][7] ) );
  DFFPOSX1 \memory_reg[18][6]  ( .D(n1118), .CLK(CLK), .Q(\memory[18][6] ) );
  DFFPOSX1 \memory_reg[18][5]  ( .D(n1117), .CLK(CLK), .Q(\memory[18][5] ) );
  DFFPOSX1 \memory_reg[18][4]  ( .D(n1116), .CLK(CLK), .Q(\memory[18][4] ) );
  DFFPOSX1 \memory_reg[18][3]  ( .D(n1115), .CLK(CLK), .Q(\memory[18][3] ) );
  DFFPOSX1 \memory_reg[18][2]  ( .D(n1114), .CLK(CLK), .Q(\memory[18][2] ) );
  DFFPOSX1 \memory_reg[18][1]  ( .D(n1113), .CLK(CLK), .Q(\memory[18][1] ) );
  DFFPOSX1 \memory_reg[18][0]  ( .D(n1112), .CLK(CLK), .Q(\memory[18][0] ) );
  DFFPOSX1 \memory_reg[19][7]  ( .D(n1111), .CLK(CLK), .Q(\memory[19][7] ) );
  DFFPOSX1 \memory_reg[19][6]  ( .D(n1110), .CLK(CLK), .Q(\memory[19][6] ) );
  DFFPOSX1 \memory_reg[19][5]  ( .D(n1109), .CLK(CLK), .Q(\memory[19][5] ) );
  DFFPOSX1 \memory_reg[19][4]  ( .D(n1108), .CLK(CLK), .Q(\memory[19][4] ) );
  DFFPOSX1 \memory_reg[19][3]  ( .D(n1107), .CLK(CLK), .Q(\memory[19][3] ) );
  DFFPOSX1 \memory_reg[19][2]  ( .D(n1106), .CLK(CLK), .Q(\memory[19][2] ) );
  DFFPOSX1 \memory_reg[19][1]  ( .D(n1105), .CLK(CLK), .Q(\memory[19][1] ) );
  DFFPOSX1 \memory_reg[19][0]  ( .D(n1104), .CLK(CLK), .Q(\memory[19][0] ) );
  DFFPOSX1 \memory_reg[20][7]  ( .D(n1342), .CLK(CLK), .Q(\memory[20][7] ) );
  DFFPOSX1 \memory_reg[20][6]  ( .D(n1343), .CLK(CLK), .Q(\memory[20][6] ) );
  DFFPOSX1 \memory_reg[20][5]  ( .D(n1344), .CLK(CLK), .Q(\memory[20][5] ) );
  DFFPOSX1 \memory_reg[20][4]  ( .D(n1345), .CLK(CLK), .Q(\memory[20][4] ) );
  DFFPOSX1 \memory_reg[20][3]  ( .D(n1346), .CLK(CLK), .Q(\memory[20][3] ) );
  DFFPOSX1 \memory_reg[20][2]  ( .D(n1347), .CLK(CLK), .Q(\memory[20][2] ) );
  DFFPOSX1 \memory_reg[20][1]  ( .D(n1348), .CLK(CLK), .Q(\memory[20][1] ) );
  DFFPOSX1 \memory_reg[20][0]  ( .D(n1349), .CLK(CLK), .Q(\memory[20][0] ) );
  DFFPOSX1 \memory_reg[21][7]  ( .D(n1334), .CLK(CLK), .Q(\memory[21][7] ) );
  DFFPOSX1 \memory_reg[21][6]  ( .D(n1335), .CLK(CLK), .Q(\memory[21][6] ) );
  DFFPOSX1 \memory_reg[21][5]  ( .D(n1336), .CLK(CLK), .Q(\memory[21][5] ) );
  DFFPOSX1 \memory_reg[21][4]  ( .D(n1337), .CLK(CLK), .Q(\memory[21][4] ) );
  DFFPOSX1 \memory_reg[21][3]  ( .D(n1338), .CLK(CLK), .Q(\memory[21][3] ) );
  DFFPOSX1 \memory_reg[21][2]  ( .D(n1339), .CLK(CLK), .Q(\memory[21][2] ) );
  DFFPOSX1 \memory_reg[21][1]  ( .D(n1340), .CLK(CLK), .Q(\memory[21][1] ) );
  DFFPOSX1 \memory_reg[21][0]  ( .D(n1341), .CLK(CLK), .Q(\memory[21][0] ) );
  DFFPOSX1 \memory_reg[22][7]  ( .D(n1326), .CLK(CLK), .Q(\memory[22][7] ) );
  DFFPOSX1 \memory_reg[22][6]  ( .D(n1327), .CLK(CLK), .Q(\memory[22][6] ) );
  DFFPOSX1 \memory_reg[22][5]  ( .D(n1328), .CLK(CLK), .Q(\memory[22][5] ) );
  DFFPOSX1 \memory_reg[22][4]  ( .D(n1329), .CLK(CLK), .Q(\memory[22][4] ) );
  DFFPOSX1 \memory_reg[22][3]  ( .D(n1330), .CLK(CLK), .Q(\memory[22][3] ) );
  DFFPOSX1 \memory_reg[22][2]  ( .D(n1331), .CLK(CLK), .Q(\memory[22][2] ) );
  DFFPOSX1 \memory_reg[22][1]  ( .D(n1332), .CLK(CLK), .Q(\memory[22][1] ) );
  DFFPOSX1 \memory_reg[22][0]  ( .D(n1333), .CLK(CLK), .Q(\memory[22][0] ) );
  DFFPOSX1 \memory_reg[23][7]  ( .D(n1318), .CLK(CLK), .Q(\memory[23][7] ) );
  DFFPOSX1 \memory_reg[23][6]  ( .D(n1319), .CLK(CLK), .Q(\memory[23][6] ) );
  DFFPOSX1 \memory_reg[23][5]  ( .D(n1320), .CLK(CLK), .Q(\memory[23][5] ) );
  DFFPOSX1 \memory_reg[23][4]  ( .D(n1321), .CLK(CLK), .Q(\memory[23][4] ) );
  DFFPOSX1 \memory_reg[23][3]  ( .D(n1322), .CLK(CLK), .Q(\memory[23][3] ) );
  DFFPOSX1 \memory_reg[23][2]  ( .D(n1323), .CLK(CLK), .Q(\memory[23][2] ) );
  DFFPOSX1 \memory_reg[23][1]  ( .D(n1324), .CLK(CLK), .Q(\memory[23][1] ) );
  DFFPOSX1 \memory_reg[23][0]  ( .D(n1325), .CLK(CLK), .Q(\memory[23][0] ) );
  DFFPOSX1 \memory_reg[24][7]  ( .D(n1310), .CLK(CLK), .Q(\memory[24][7] ) );
  DFFPOSX1 \memory_reg[24][6]  ( .D(n1311), .CLK(CLK), .Q(\memory[24][6] ) );
  DFFPOSX1 \memory_reg[24][5]  ( .D(n1312), .CLK(CLK), .Q(\memory[24][5] ) );
  DFFPOSX1 \memory_reg[24][4]  ( .D(n1313), .CLK(CLK), .Q(\memory[24][4] ) );
  DFFPOSX1 \memory_reg[24][3]  ( .D(n1314), .CLK(CLK), .Q(\memory[24][3] ) );
  DFFPOSX1 \memory_reg[24][2]  ( .D(n1315), .CLK(CLK), .Q(\memory[24][2] ) );
  DFFPOSX1 \memory_reg[24][1]  ( .D(n1316), .CLK(CLK), .Q(\memory[24][1] ) );
  DFFPOSX1 \memory_reg[24][0]  ( .D(n1317), .CLK(CLK), .Q(\memory[24][0] ) );
  DFFPOSX1 \memory_reg[25][7]  ( .D(n1302), .CLK(CLK), .Q(\memory[25][7] ) );
  DFFPOSX1 \memory_reg[25][6]  ( .D(n1303), .CLK(CLK), .Q(\memory[25][6] ) );
  DFFPOSX1 \memory_reg[25][5]  ( .D(n1304), .CLK(CLK), .Q(\memory[25][5] ) );
  DFFPOSX1 \memory_reg[25][4]  ( .D(n1305), .CLK(CLK), .Q(\memory[25][4] ) );
  DFFPOSX1 \memory_reg[25][3]  ( .D(n1306), .CLK(CLK), .Q(\memory[25][3] ) );
  DFFPOSX1 \memory_reg[25][2]  ( .D(n1307), .CLK(CLK), .Q(\memory[25][2] ) );
  DFFPOSX1 \memory_reg[25][1]  ( .D(n1308), .CLK(CLK), .Q(\memory[25][1] ) );
  DFFPOSX1 \memory_reg[25][0]  ( .D(n1309), .CLK(CLK), .Q(\memory[25][0] ) );
  DFFPOSX1 \memory_reg[26][7]  ( .D(n1294), .CLK(CLK), .Q(\memory[26][7] ) );
  DFFPOSX1 \memory_reg[26][6]  ( .D(n1295), .CLK(CLK), .Q(\memory[26][6] ) );
  DFFPOSX1 \memory_reg[26][5]  ( .D(n1296), .CLK(CLK), .Q(\memory[26][5] ) );
  DFFPOSX1 \memory_reg[26][4]  ( .D(n1297), .CLK(CLK), .Q(\memory[26][4] ) );
  DFFPOSX1 \memory_reg[26][3]  ( .D(n1298), .CLK(CLK), .Q(\memory[26][3] ) );
  DFFPOSX1 \memory_reg[26][2]  ( .D(n1299), .CLK(CLK), .Q(\memory[26][2] ) );
  DFFPOSX1 \memory_reg[26][1]  ( .D(n1300), .CLK(CLK), .Q(\memory[26][1] ) );
  DFFPOSX1 \memory_reg[26][0]  ( .D(n1301), .CLK(CLK), .Q(\memory[26][0] ) );
  DFFPOSX1 \memory_reg[27][7]  ( .D(n1286), .CLK(CLK), .Q(\memory[27][7] ) );
  DFFPOSX1 \memory_reg[27][6]  ( .D(n1287), .CLK(CLK), .Q(\memory[27][6] ) );
  DFFPOSX1 \memory_reg[27][5]  ( .D(n1288), .CLK(CLK), .Q(\memory[27][5] ) );
  DFFPOSX1 \memory_reg[27][4]  ( .D(n1289), .CLK(CLK), .Q(\memory[27][4] ) );
  DFFPOSX1 \memory_reg[27][3]  ( .D(n1290), .CLK(CLK), .Q(\memory[27][3] ) );
  DFFPOSX1 \memory_reg[27][2]  ( .D(n1291), .CLK(CLK), .Q(\memory[27][2] ) );
  DFFPOSX1 \memory_reg[27][1]  ( .D(n1292), .CLK(CLK), .Q(\memory[27][1] ) );
  DFFPOSX1 \memory_reg[27][0]  ( .D(n1293), .CLK(CLK), .Q(\memory[27][0] ) );
  DFFPOSX1 \memory_reg[28][7]  ( .D(n1103), .CLK(CLK), .Q(\memory[28][7] ) );
  DFFPOSX1 \memory_reg[28][6]  ( .D(n1102), .CLK(CLK), .Q(\memory[28][6] ) );
  DFFPOSX1 \memory_reg[28][5]  ( .D(n1101), .CLK(CLK), .Q(\memory[28][5] ) );
  DFFPOSX1 \memory_reg[28][4]  ( .D(n1100), .CLK(CLK), .Q(\memory[28][4] ) );
  DFFPOSX1 \memory_reg[28][3]  ( .D(n1099), .CLK(CLK), .Q(\memory[28][3] ) );
  DFFPOSX1 \memory_reg[28][2]  ( .D(n1098), .CLK(CLK), .Q(\memory[28][2] ) );
  DFFPOSX1 \memory_reg[28][1]  ( .D(n1097), .CLK(CLK), .Q(\memory[28][1] ) );
  DFFPOSX1 \memory_reg[28][0]  ( .D(n1096), .CLK(CLK), .Q(\memory[28][0] ) );
  DFFPOSX1 \memory_reg[29][7]  ( .D(n1095), .CLK(CLK), .Q(\memory[29][7] ) );
  DFFPOSX1 \memory_reg[29][6]  ( .D(n1094), .CLK(CLK), .Q(\memory[29][6] ) );
  DFFPOSX1 \memory_reg[29][5]  ( .D(n1093), .CLK(CLK), .Q(\memory[29][5] ) );
  DFFPOSX1 \memory_reg[29][4]  ( .D(n1092), .CLK(CLK), .Q(\memory[29][4] ) );
  DFFPOSX1 \memory_reg[29][3]  ( .D(n1091), .CLK(CLK), .Q(\memory[29][3] ) );
  DFFPOSX1 \memory_reg[29][2]  ( .D(n1090), .CLK(CLK), .Q(\memory[29][2] ) );
  DFFPOSX1 \memory_reg[29][1]  ( .D(n1089), .CLK(CLK), .Q(\memory[29][1] ) );
  DFFPOSX1 \memory_reg[29][0]  ( .D(n1088), .CLK(CLK), .Q(\memory[29][0] ) );
  DFFPOSX1 \memory_reg[30][7]  ( .D(n1087), .CLK(CLK), .Q(\memory[30][7] ) );
  DFFPOSX1 \memory_reg[30][6]  ( .D(n1086), .CLK(CLK), .Q(\memory[30][6] ) );
  DFFPOSX1 \memory_reg[30][5]  ( .D(n1085), .CLK(CLK), .Q(\memory[30][5] ) );
  DFFPOSX1 \memory_reg[30][4]  ( .D(n1084), .CLK(CLK), .Q(\memory[30][4] ) );
  DFFPOSX1 \memory_reg[30][3]  ( .D(n1083), .CLK(CLK), .Q(\memory[30][3] ) );
  DFFPOSX1 \memory_reg[30][2]  ( .D(n1082), .CLK(CLK), .Q(\memory[30][2] ) );
  DFFPOSX1 \memory_reg[30][1]  ( .D(n1081), .CLK(CLK), .Q(\memory[30][1] ) );
  DFFPOSX1 \memory_reg[30][0]  ( .D(n1080), .CLK(CLK), .Q(\memory[30][0] ) );
  DFFPOSX1 \memory_reg[31][7]  ( .D(n1079), .CLK(CLK), .Q(\memory[31][7] ) );
  DFFPOSX1 \memory_reg[31][6]  ( .D(n1078), .CLK(CLK), .Q(\memory[31][6] ) );
  DFFPOSX1 \memory_reg[31][5]  ( .D(n1077), .CLK(CLK), .Q(\memory[31][5] ) );
  DFFPOSX1 \memory_reg[31][4]  ( .D(n1076), .CLK(CLK), .Q(\memory[31][4] ) );
  DFFPOSX1 \memory_reg[31][3]  ( .D(n1075), .CLK(CLK), .Q(\memory[31][3] ) );
  DFFPOSX1 \memory_reg[31][2]  ( .D(n1074), .CLK(CLK), .Q(\memory[31][2] ) );
  DFFPOSX1 \memory_reg[31][1]  ( .D(n1073), .CLK(CLK), .Q(\memory[31][1] ) );
  DFFPOSX1 \memory_reg[31][0]  ( .D(n1072), .CLK(CLK), .Q(\memory[31][0] ) );
  DFFPOSX1 \opcode_reg[0][1]  ( .D(n610), .CLK(CLK), .Q(\opcode[0][1] ) );
  DFFPOSX1 \opcode_reg[0][0]  ( .D(n611), .CLK(CLK), .Q(\opcode[0][0] ) );
  DFFPOSX1 \opcode_reg[1][1]  ( .D(n652), .CLK(CLK), .Q(\opcode[1][1] ) );
  DFFPOSX1 \opcode_reg[1][0]  ( .D(n653), .CLK(CLK), .Q(\opcode[1][0] ) );
  DFFPOSX1 \opcode_reg[2][1]  ( .D(n654), .CLK(CLK), .Q(\opcode[2][1] ) );
  DFFPOSX1 \opcode_reg[2][0]  ( .D(n655), .CLK(CLK), .Q(\opcode[2][0] ) );
  DFFPOSX1 \opcode_reg[3][1]  ( .D(n624), .CLK(CLK), .Q(\opcode[3][1] ) );
  DFFPOSX1 \opcode_reg[3][0]  ( .D(n625), .CLK(CLK), .Q(\opcode[3][0] ) );
  DFFPOSX1 \opcode_reg[4][1]  ( .D(n640), .CLK(CLK), .Q(\opcode[4][1] ) );
  DFFPOSX1 \opcode_reg[4][0]  ( .D(n641), .CLK(CLK), .Q(\opcode[4][0] ) );
  DFFPOSX1 \opcode_reg[5][1]  ( .D(n614), .CLK(CLK), .Q(\opcode[5][1] ) );
  DFFPOSX1 \opcode_reg[5][0]  ( .D(n615), .CLK(CLK), .Q(\opcode[5][0] ) );
  DFFPOSX1 \opcode_reg[6][1]  ( .D(n600), .CLK(CLK), .Q(\opcode[6][1] ) );
  DFFPOSX1 \opcode_reg[6][0]  ( .D(n601), .CLK(CLK), .Q(\opcode[6][0] ) );
  DFFPOSX1 \opcode_reg[7][1]  ( .D(n608), .CLK(CLK), .Q(\opcode[7][1] ) );
  DFFPOSX1 \opcode_reg[7][0]  ( .D(n609), .CLK(CLK), .Q(\opcode[7][0] ) );
  DFFPOSX1 \opcode_reg[8][1]  ( .D(n634), .CLK(CLK), .Q(\opcode[8][1] ) );
  DFFPOSX1 \opcode_reg[8][0]  ( .D(n635), .CLK(CLK), .Q(\opcode[8][0] ) );
  DFFPOSX1 \opcode_reg[9][1]  ( .D(n622), .CLK(CLK), .Q(\opcode[9][1] ) );
  DFFPOSX1 \opcode_reg[9][0]  ( .D(n623), .CLK(CLK), .Q(\opcode[9][0] ) );
  DFFPOSX1 \opcode_reg[10][1]  ( .D(n646), .CLK(CLK), .Q(\opcode[10][1] ) );
  DFFPOSX1 \opcode_reg[10][0]  ( .D(n647), .CLK(CLK), .Q(\opcode[10][0] ) );
  DFFPOSX1 \opcode_reg[11][1]  ( .D(n1057), .CLK(CLK), .Q(\opcode[11][1] ) );
  DFFPOSX1 \opcode_reg[11][0]  ( .D(n1056), .CLK(CLK), .Q(\opcode[11][0] ) );
  DFFPOSX1 \opcode_reg[12][1]  ( .D(n642), .CLK(CLK), .Q(\opcode[12][1] ) );
  DFFPOSX1 \opcode_reg[12][0]  ( .D(n643), .CLK(CLK), .Q(\opcode[12][0] ) );
  DFFPOSX1 \opcode_reg[13][1]  ( .D(n638), .CLK(CLK), .Q(\opcode[13][1] ) );
  DFFPOSX1 \opcode_reg[13][0]  ( .D(n639), .CLK(CLK), .Q(\opcode[13][0] ) );
  DFFPOSX1 \opcode_reg[14][1]  ( .D(n636), .CLK(CLK), .Q(\opcode[14][1] ) );
  DFFPOSX1 \opcode_reg[14][0]  ( .D(n637), .CLK(CLK), .Q(\opcode[14][0] ) );
  DFFPOSX1 \opcode_reg[15][1]  ( .D(n648), .CLK(CLK), .Q(\opcode[15][1] ) );
  DFFPOSX1 \opcode_reg[15][0]  ( .D(n649), .CLK(CLK), .Q(\opcode[15][0] ) );
  DFFPOSX1 \opcode_reg[16][1]  ( .D(n626), .CLK(CLK), .Q(\opcode[16][1] ) );
  DFFPOSX1 \opcode_reg[16][0]  ( .D(n627), .CLK(CLK), .Q(\opcode[16][0] ) );
  DFFPOSX1 \opcode_reg[17][1]  ( .D(n612), .CLK(CLK), .Q(\opcode[17][1] ) );
  DFFPOSX1 \opcode_reg[17][0]  ( .D(n613), .CLK(CLK), .Q(\opcode[17][0] ) );
  DFFPOSX1 \opcode_reg[18][1]  ( .D(n602), .CLK(CLK), .Q(\opcode[18][1] ) );
  DFFPOSX1 \opcode_reg[18][0]  ( .D(n603), .CLK(CLK), .Q(\opcode[18][0] ) );
  DFFPOSX1 \opcode_reg[19][1]  ( .D(n628), .CLK(CLK), .Q(\opcode[19][1] ) );
  DFFPOSX1 \opcode_reg[19][0]  ( .D(n629), .CLK(CLK), .Q(\opcode[19][0] ) );
  DFFPOSX1 \opcode_reg[20][1]  ( .D(n658), .CLK(CLK), .Q(\opcode[20][1] ) );
  DFFPOSX1 \opcode_reg[20][0]  ( .D(n659), .CLK(CLK), .Q(\opcode[20][0] ) );
  DFFPOSX1 \opcode_reg[21][1]  ( .D(n660), .CLK(CLK), .Q(\opcode[21][1] ) );
  DFFPOSX1 \opcode_reg[21][0]  ( .D(n661), .CLK(CLK), .Q(\opcode[21][0] ) );
  DFFPOSX1 \opcode_reg[22][1]  ( .D(n620), .CLK(CLK), .Q(\opcode[22][1] ) );
  DFFPOSX1 \opcode_reg[22][0]  ( .D(n621), .CLK(CLK), .Q(\opcode[22][0] ) );
  DFFPOSX1 \opcode_reg[23][1]  ( .D(n618), .CLK(CLK), .Q(\opcode[23][1] ) );
  DFFPOSX1 \opcode_reg[23][0]  ( .D(n619), .CLK(CLK), .Q(\opcode[23][0] ) );
  DFFPOSX1 \opcode_reg[24][1]  ( .D(n606), .CLK(CLK), .Q(\opcode[24][1] ) );
  DFFPOSX1 \opcode_reg[24][0]  ( .D(n607), .CLK(CLK), .Q(\opcode[24][0] ) );
  DFFPOSX1 \opcode_reg[25][1]  ( .D(n656), .CLK(CLK), .Q(\opcode[25][1] ) );
  DFFPOSX1 \opcode_reg[25][0]  ( .D(n657), .CLK(CLK), .Q(\opcode[25][0] ) );
  DFFPOSX1 \opcode_reg[26][1]  ( .D(n630), .CLK(CLK), .Q(\opcode[26][1] ) );
  DFFPOSX1 \opcode_reg[26][0]  ( .D(n631), .CLK(CLK), .Q(\opcode[26][0] ) );
  DFFPOSX1 \opcode_reg[27][1]  ( .D(n650), .CLK(CLK), .Q(\opcode[27][1] ) );
  DFFPOSX1 \opcode_reg[27][0]  ( .D(n651), .CLK(CLK), .Q(\opcode[27][0] ) );
  DFFPOSX1 \opcode_reg[28][1]  ( .D(n644), .CLK(CLK), .Q(\opcode[28][1] ) );
  DFFPOSX1 \opcode_reg[28][0]  ( .D(n645), .CLK(CLK), .Q(\opcode[28][0] ) );
  DFFPOSX1 \opcode_reg[29][1]  ( .D(n632), .CLK(CLK), .Q(\opcode[29][1] ) );
  DFFPOSX1 \opcode_reg[29][0]  ( .D(n633), .CLK(CLK), .Q(\opcode[29][0] ) );
  DFFPOSX1 \opcode_reg[30][1]  ( .D(n616), .CLK(CLK), .Q(\opcode[30][1] ) );
  DFFPOSX1 \opcode_reg[30][0]  ( .D(n617), .CLK(CLK), .Q(\opcode[30][0] ) );
  DFFPOSX1 \opcode_reg[31][1]  ( .D(n604), .CLK(CLK), .Q(\opcode[31][1] ) );
  DFFPOSX1 \opcode_reg[31][0]  ( .D(n605), .CLK(CLK), .Q(\opcode[31][0] ) );
  DFFPOSX1 \DATA_reg[7]  ( .D(n1039), .CLK(CLK), .Q(DATA[7]) );
  DFFPOSX1 \DATA_reg[6]  ( .D(n1038), .CLK(CLK), .Q(DATA[6]) );
  DFFPOSX1 \DATA_reg[5]  ( .D(n1037), .CLK(CLK), .Q(DATA[5]) );
  DFFPOSX1 \DATA_reg[4]  ( .D(n1036), .CLK(CLK), .Q(DATA[4]) );
  DFFPOSX1 \DATA_reg[3]  ( .D(n1035), .CLK(CLK), .Q(DATA[3]) );
  DFFPOSX1 \DATA_reg[2]  ( .D(n1034), .CLK(CLK), .Q(DATA[2]) );
  DFFPOSX1 \DATA_reg[1]  ( .D(n1033), .CLK(CLK), .Q(DATA[1]) );
  DFFPOSX1 \DATA_reg[0]  ( .D(n1032), .CLK(CLK), .Q(DATA[0]) );
  DFFPOSX1 \OUT_OPCODE_reg[1]  ( .D(n1031), .CLK(CLK), .Q(OUT_OPCODE[1]) );
  DFFPOSX1 \OUT_OPCODE_reg[0]  ( .D(n1030), .CLK(CLK), .Q(OUT_OPCODE[0]) );
  DFFPOSX1 EMPTY_reg ( .D(n1415), .CLK(CLK), .Q(EMPTY) );
  DFFSR \readptr_reg[2]  ( .D(N345), .CLK(CLK), .R(n177), .S(1'b1), .Q(
        readptr[2]) );
  INVX1 U3 ( .A(n94), .Y(n568) );
  INVX4 U4 ( .A(n50), .Y(n51) );
  INVX2 U5 ( .A(n338), .Y(n512) );
  INVX2 U6 ( .A(n348), .Y(n514) );
  INVX2 U7 ( .A(n248), .Y(n1) );
  INVX2 U8 ( .A(n248), .Y(n33) );
  AND2X1 U9 ( .A(n2), .B(writeptr[1]), .Y(n86) );
  BUFX2 U10 ( .A(writeptr[0]), .Y(n2) );
  INVX1 U11 ( .A(writeptr[0]), .Y(n230) );
  INVX4 U12 ( .A(n338), .Y(n3) );
  INVX4 U13 ( .A(n348), .Y(n4) );
  INVX1 U14 ( .A(n542), .Y(n5) );
  INVX2 U15 ( .A(n5), .Y(n6) );
  INVX1 U16 ( .A(n573), .Y(n7) );
  INVX2 U17 ( .A(n7), .Y(n8) );
  BUFX4 U18 ( .A(n106), .Y(n92) );
  MUX2X1 U19 ( .B(n170), .A(\opcode[6][0] ), .S(n323), .Y(n324) );
  INVX2 U20 ( .A(n323), .Y(n492) );
  MUX2X1 U21 ( .B(n170), .A(\opcode[2][0] ), .S(n343), .Y(n344) );
  INVX2 U22 ( .A(n29), .Y(n555) );
  INVX2 U23 ( .A(n348), .Y(n48) );
  INVX2 U24 ( .A(n338), .Y(n47) );
  AND2X2 U25 ( .A(n1262), .B(n120), .Y(n9) );
  AND2X1 U26 ( .A(n1273), .B(n120), .Y(n10) );
  AND2X2 U27 ( .A(n1283), .B(n120), .Y(n11) );
  AND2X2 U28 ( .A(n1252), .B(n1262), .Y(n12) );
  AND2X2 U29 ( .A(n1282), .B(n1252), .Y(n13) );
  AND2X1 U30 ( .A(n1273), .B(n1252), .Y(n14) );
  AND2X1 U31 ( .A(n1253), .B(n1252), .Y(n15) );
  AND2X2 U32 ( .A(n1274), .B(n1252), .Y(n16) );
  AND2X2 U33 ( .A(n1283), .B(n1252), .Y(n17) );
  AND2X1 U34 ( .A(n1252), .B(n1263), .Y(n18) );
  AND2X1 U35 ( .A(n1253), .B(n120), .Y(n19) );
  AND2X1 U36 ( .A(n1274), .B(n120), .Y(n20) );
  AND2X1 U37 ( .A(n1263), .B(n120), .Y(n21) );
  AND2X2 U38 ( .A(n1282), .B(n120), .Y(n22) );
  INVX1 U39 ( .A(RCV_DATA[0]), .Y(n515) );
  INVX1 U40 ( .A(RCV_DATA[1]), .Y(n516) );
  INVX1 U41 ( .A(RCV_DATA[3]), .Y(n517) );
  INVX1 U42 ( .A(RCV_DATA[5]), .Y(n519) );
  INVX1 U44 ( .A(n553), .Y(n554) );
  INVX1 U45 ( .A(RCV_DATA[4]), .Y(n518) );
  INVX2 U46 ( .A(n225), .Y(n24) );
  INVX2 U47 ( .A(n225), .Y(n394) );
  INVX1 U48 ( .A(n230), .Y(n25) );
  INVX1 U49 ( .A(n547), .Y(n26) );
  INVX2 U50 ( .A(n26), .Y(n27) );
  BUFX2 U51 ( .A(n537), .Y(n28) );
  INVX1 U52 ( .A(RCV_DATA[6]), .Y(n520) );
  AND2X2 U53 ( .A(n2), .B(writeptr[1]), .Y(n29) );
  INVX1 U54 ( .A(RCV_DATA[7]), .Y(n521) );
  INVX1 U55 ( .A(n149), .Y(n229) );
  BUFX2 U56 ( .A(n107), .Y(n30) );
  INVX2 U57 ( .A(n272), .Y(n31) );
  INVX2 U58 ( .A(n272), .Y(n434) );
  AND2X2 U59 ( .A(n271), .B(n308), .Y(n32) );
  INVX2 U60 ( .A(n244), .Y(n34) );
  INVX2 U61 ( .A(n244), .Y(n404) );
  NOR2X1 U62 ( .A(n87), .B(n85), .Y(n35) );
  INVX4 U63 ( .A(n663), .Y(n36) );
  INVX1 U64 ( .A(n82), .Y(n37) );
  XNOR2X1 U65 ( .A(n547), .B(n36), .Y(n90) );
  INVX1 U66 ( .A(n566), .Y(n38) );
  INVX4 U67 ( .A(n41), .Y(n73) );
  INVX2 U68 ( .A(n333), .Y(n39) );
  INVX2 U69 ( .A(n343), .Y(n40) );
  NAND2X1 U70 ( .A(n271), .B(n308), .Y(n41) );
  INVX2 U71 ( .A(n264), .Y(n42) );
  INVX2 U72 ( .A(n264), .Y(n43) );
  INVX2 U73 ( .A(n264), .Y(n433) );
  INVX2 U74 ( .A(n256), .Y(n44) );
  INVX2 U75 ( .A(n256), .Y(n430) );
  INVX2 U76 ( .A(n252), .Y(n45) );
  INVX2 U77 ( .A(n252), .Y(n46) );
  INVX2 U78 ( .A(n252), .Y(n421) );
  INVX1 U79 ( .A(n574), .Y(n49) );
  INVX1 U80 ( .A(writeptr[4]), .Y(n574) );
  INVX2 U81 ( .A(readptr[1]), .Y(n50) );
  BUFX2 U82 ( .A(n37), .Y(n52) );
  NAND2X1 U83 ( .A(RCV_OPCODE[1]), .B(RCV_OPCODE[0]), .Y(n53) );
  NAND2X1 U84 ( .A(RCV_OPCODE[0]), .B(RCV_OPCODE[1]), .Y(n54) );
  INVX2 U85 ( .A(n243), .Y(n55) );
  INVX2 U86 ( .A(n243), .Y(n271) );
  INVX2 U87 ( .A(n260), .Y(n56) );
  INVX2 U88 ( .A(n260), .Y(n432) );
  INVX2 U89 ( .A(n323), .Y(n57) );
  INVX2 U90 ( .A(n323), .Y(n58) );
  INVX1 U91 ( .A(n235), .Y(n59) );
  INVX1 U92 ( .A(n231), .Y(n60) );
  INVX1 U93 ( .A(n221), .Y(n61) );
  INVX1 U94 ( .A(n216), .Y(n62) );
  INVX1 U95 ( .A(n211), .Y(n63) );
  INVX2 U96 ( .A(n207), .Y(n64) );
  INVX2 U97 ( .A(n207), .Y(n365) );
  INVX4 U98 ( .A(n284), .Y(n65) );
  INVX2 U99 ( .A(n284), .Y(n451) );
  INVX4 U100 ( .A(n328), .Y(n66) );
  INVX2 U101 ( .A(n328), .Y(n501) );
  INVX2 U102 ( .A(n279), .Y(n67) );
  INVX2 U103 ( .A(n279), .Y(n442) );
  AND2X2 U104 ( .A(n239), .B(n353), .Y(n106) );
  NAND2X1 U105 ( .A(n578), .B(n68), .Y(n577) );
  NOR2X1 U106 ( .A(n565), .B(n94), .Y(n68) );
  AND2X2 U107 ( .A(n353), .B(n354), .Y(n69) );
  AND2X2 U108 ( .A(n353), .B(n354), .Y(n70) );
  INVX2 U109 ( .A(n333), .Y(n71) );
  INVX4 U110 ( .A(n333), .Y(n510) );
  INVX4 U111 ( .A(n343), .Y(n513) );
  INVX2 U112 ( .A(n577), .Y(n583) );
  BUFX2 U113 ( .A(n555), .Y(n72) );
  INVX2 U114 ( .A(readptr[0]), .Y(n74) );
  INVX2 U115 ( .A(n74), .Y(n75) );
  INVX1 U116 ( .A(n74), .Y(n76) );
  INVX4 U117 ( .A(n51), .Y(n594) );
  AND2X2 U118 ( .A(n51), .B(n663), .Y(n120) );
  AND2X2 U119 ( .A(n51), .B(n36), .Y(n121) );
  INVX1 U120 ( .A(n150), .Y(n77) );
  INVX2 U121 ( .A(n569), .Y(n78) );
  INVX4 U122 ( .A(n150), .Y(n151) );
  AND2X1 U123 ( .A(n563), .B(n562), .Y(n564) );
  INVX1 U124 ( .A(n558), .Y(n89) );
  INVX4 U125 ( .A(n278), .Y(n472) );
  INVX4 U126 ( .A(n206), .Y(n239) );
  AND2X2 U127 ( .A(n353), .B(n354), .Y(n79) );
  AND2X2 U128 ( .A(n353), .B(n354), .Y(n80) );
  AND2X2 U129 ( .A(R_ENABLE), .B(n181), .Y(n81) );
  INVX2 U130 ( .A(n81), .Y(n597) );
  BUFX2 U131 ( .A(n230), .Y(n82) );
  INVX2 U132 ( .A(n471), .Y(n83) );
  BUFX4 U133 ( .A(readptr[4]), .Y(n84) );
  AND2X2 U134 ( .A(n524), .B(n178), .Y(n85) );
  INVX1 U135 ( .A(n85), .Y(n522) );
  XOR2X1 U136 ( .A(n317), .B(n88), .Y(n87) );
  INVX1 U137 ( .A(n87), .Y(n541) );
  XNOR2X1 U138 ( .A(n94), .B(n153), .Y(n88) );
  INVX1 U139 ( .A(n558), .Y(n581) );
  INVX1 U140 ( .A(n90), .Y(n540) );
  INVX1 U141 ( .A(n77), .Y(n215) );
  INVX8 U142 ( .A(n148), .Y(n149) );
  NAND3X1 U143 ( .A(n90), .B(n35), .C(n204), .Y(n91) );
  BUFX4 U144 ( .A(n106), .Y(n93) );
  BUFX4 U145 ( .A(writeptr[3]), .Y(n94) );
  INVX2 U146 ( .A(n21), .Y(n131) );
  INVX2 U147 ( .A(n18), .Y(n143) );
  INVX2 U148 ( .A(n14), .Y(n144) );
  INVX2 U149 ( .A(n19), .Y(n128) );
  INVX2 U150 ( .A(n20), .Y(n133) );
  AND2X1 U151 ( .A(writeptr[4]), .B(n124), .Y(n122) );
  AND2X2 U152 ( .A(n578), .B(n353), .Y(n95) );
  INVX2 U153 ( .A(n172), .Y(n170) );
  INVX2 U154 ( .A(n176), .Y(n174) );
  INVX2 U155 ( .A(n176), .Y(n173) );
  AND2X2 U156 ( .A(n308), .B(n578), .Y(n96) );
  AND2X2 U157 ( .A(n472), .B(n471), .Y(n97) );
  AND2X2 U158 ( .A(n569), .B(n578), .Y(n98) );
  AND2X2 U159 ( .A(n471), .B(n578), .Y(n99) );
  AND2X2 U160 ( .A(n293), .B(n578), .Y(n100) );
  AND2X2 U161 ( .A(n283), .B(n578), .Y(n101) );
  AND2X2 U162 ( .A(n303), .B(n578), .Y(n102) );
  INVX2 U163 ( .A(RCV_OPCODE[0]), .Y(n172) );
  INVX1 U164 ( .A(RCV_OPCODE[1]), .Y(n176) );
  AND2X2 U165 ( .A(n277), .B(W_ENABLE), .Y(n103) );
  AND2X2 U166 ( .A(W_ENABLE), .B(n91), .Y(n104) );
  AND2X2 U167 ( .A(n288), .B(n578), .Y(n105) );
  AND2X2 U168 ( .A(n148), .B(n2), .Y(n107) );
  INVX2 U169 ( .A(RST), .Y(n177) );
  AND2X2 U170 ( .A(n276), .B(n574), .Y(n108) );
  AND2X2 U171 ( .A(n1283), .B(n121), .Y(n109) );
  AND2X2 U172 ( .A(n1253), .B(n121), .Y(n110) );
  AND2X2 U173 ( .A(n1274), .B(n121), .Y(n111) );
  AND2X2 U174 ( .A(n1263), .B(n121), .Y(n112) );
  AND2X2 U175 ( .A(n1282), .B(n121), .Y(n113) );
  AND2X2 U176 ( .A(n1251), .B(n121), .Y(n114) );
  AND2X2 U177 ( .A(n1262), .B(n121), .Y(n115) );
  AND2X2 U178 ( .A(n1273), .B(n121), .Y(n116) );
  XNOR2X1 U179 ( .A(n573), .B(n537), .Y(n542) );
  AND2X2 U180 ( .A(n124), .B(n574), .Y(n117) );
  INVX2 U181 ( .A(n12), .Y(n142) );
  INVX4 U182 ( .A(n13), .Y(n146) );
  INVX2 U183 ( .A(n139), .Y(n140) );
  INVX1 U184 ( .A(n838), .Y(n139) );
  INVX4 U185 ( .A(n16), .Y(n145) );
  INVX4 U186 ( .A(n17), .Y(n147) );
  INVX2 U187 ( .A(n15), .Y(n141) );
  INVX4 U188 ( .A(n22), .Y(n136) );
  INVX2 U189 ( .A(n129), .Y(n130) );
  INVX1 U190 ( .A(n839), .Y(n129) );
  INVX2 U191 ( .A(n9), .Y(n132) );
  INVX2 U192 ( .A(n10), .Y(n134) );
  INVX4 U193 ( .A(n11), .Y(n135) );
  INVX2 U194 ( .A(n119), .Y(n137) );
  INVX2 U195 ( .A(n119), .Y(n138) );
  INVX2 U196 ( .A(n155), .Y(n154) );
  INVX2 U197 ( .A(n157), .Y(n156) );
  INVX2 U198 ( .A(RCV_DATA[2]), .Y(n158) );
  INVX2 U199 ( .A(RCV_DATA[2]), .Y(n159) );
  INVX2 U200 ( .A(n161), .Y(n160) );
  INVX2 U201 ( .A(n165), .Y(n164) );
  INVX2 U202 ( .A(n163), .Y(n162) );
  INVX2 U203 ( .A(n167), .Y(n166) );
  INVX2 U204 ( .A(n169), .Y(n168) );
  AND2X2 U205 ( .A(writeptr[4]), .B(n276), .Y(n118) );
  OR2X2 U206 ( .A(n597), .B(n182), .Y(n119) );
  XOR2X1 U207 ( .A(n151), .B(n51), .Y(n123) );
  INVX2 U208 ( .A(writeptr[1]), .Y(n150) );
  INVX2 U209 ( .A(readptr[3]), .Y(n152) );
  NOR2X1 U210 ( .A(RST), .B(n94), .Y(n124) );
  INVX2 U211 ( .A(n517), .Y(n161) );
  INVX2 U212 ( .A(n519), .Y(n165) );
  INVX2 U213 ( .A(n515), .Y(n155) );
  INVX2 U214 ( .A(n516), .Y(n157) );
  INVX2 U215 ( .A(n518), .Y(n163) );
  INVX2 U216 ( .A(n520), .Y(n167) );
  INVX2 U217 ( .A(n521), .Y(n169) );
  BUFX2 U218 ( .A(n352), .Y(n125) );
  BUFX4 U219 ( .A(n352), .Y(n126) );
  INVX2 U220 ( .A(writeptr[2]), .Y(n148) );
  INVX1 U221 ( .A(n337), .Y(n471) );
  INVX1 U222 ( .A(n317), .Y(n569) );
  INVX1 U223 ( .A(n172), .Y(n171) );
  INVX1 U224 ( .A(n176), .Y(n175) );
  INVX4 U225 ( .A(n318), .Y(n127) );
  INVX2 U226 ( .A(n318), .Y(n483) );
  INVX4 U227 ( .A(n563), .Y(n578) );
  INVX4 U228 ( .A(n211), .Y(n374) );
  INVX4 U229 ( .A(n216), .Y(n383) );
  INVX4 U230 ( .A(n221), .Y(n392) );
  INVX4 U231 ( .A(n231), .Y(n395) );
  INVX4 U232 ( .A(n235), .Y(n396) );
  INVX4 U233 ( .A(n289), .Y(n460) );
  INVX4 U234 ( .A(n294), .Y(n469) );
  INVX4 U235 ( .A(n304), .Y(n473) );
  INVX4 U236 ( .A(n309), .Y(n474) );
  INVX4 U237 ( .A(n313), .Y(n475) );
  AND2X2 U238 ( .A(n1253), .B(n1254), .Y(n841) );
  AND2X2 U239 ( .A(n1251), .B(n1254), .Y(n840) );
  AND2X2 U240 ( .A(n1254), .B(n1263), .Y(n865) );
  AND2X2 U241 ( .A(n1254), .B(n1262), .Y(n852) );
  AND2X2 U242 ( .A(n1274), .B(n1254), .Y(n909) );
  AND2X2 U243 ( .A(n1273), .B(n1254), .Y(n908) );
  AND2X2 U244 ( .A(n1283), .B(n1254), .Y(n916) );
  AND2X2 U245 ( .A(n1282), .B(n1254), .Y(n915) );
  INVX8 U246 ( .A(n152), .Y(n153) );
  INVX2 U247 ( .A(\memory[16][7] ), .Y(n780) );
  INVX2 U248 ( .A(\memory[17][7] ), .Y(n788) );
  INVX2 U249 ( .A(\memory[18][7] ), .Y(n796) );
  INVX2 U250 ( .A(readptr[2]), .Y(n663) );
  INVX2 U251 ( .A(\memory[19][7] ), .Y(n804) );
  NAND2X1 U252 ( .A(n1251), .B(n120), .Y(n839) );
  INVX2 U253 ( .A(\memory[24][7] ), .Y(n706) );
  INVX2 U254 ( .A(\memory[25][7] ), .Y(n698) );
  INVX2 U255 ( .A(\memory[26][7] ), .Y(n690) );
  INVX2 U256 ( .A(\memory[27][7] ), .Y(n682) );
  INVX2 U257 ( .A(\memory[3][7] ), .Y(n745) );
  INVX2 U258 ( .A(\memory[2][7] ), .Y(n737) );
  INVX2 U259 ( .A(\memory[1][7] ), .Y(n729) );
  INVX2 U260 ( .A(\memory[0][7] ), .Y(n721) );
  INVX2 U261 ( .A(\memory[8][7] ), .Y(n748) );
  INVX2 U262 ( .A(\memory[9][7] ), .Y(n756) );
  INVX2 U263 ( .A(\memory[10][7] ), .Y(n764) );
  INVX2 U264 ( .A(\memory[11][7] ), .Y(n772) );
  INVX2 U265 ( .A(\memory[16][6] ), .Y(n781) );
  INVX2 U266 ( .A(\memory[17][6] ), .Y(n789) );
  INVX2 U267 ( .A(\memory[18][6] ), .Y(n797) );
  INVX2 U268 ( .A(\memory[19][6] ), .Y(n805) );
  INVX2 U269 ( .A(\memory[24][6] ), .Y(n707) );
  INVX2 U270 ( .A(\memory[25][6] ), .Y(n699) );
  INVX2 U271 ( .A(\memory[26][6] ), .Y(n691) );
  INVX2 U272 ( .A(\memory[27][6] ), .Y(n683) );
  INVX2 U273 ( .A(\memory[3][6] ), .Y(n744) );
  INVX2 U274 ( .A(\memory[2][6] ), .Y(n736) );
  INVX2 U275 ( .A(\memory[1][6] ), .Y(n728) );
  INVX2 U276 ( .A(\memory[0][6] ), .Y(n720) );
  INVX2 U277 ( .A(\memory[8][6] ), .Y(n749) );
  INVX2 U278 ( .A(\memory[9][6] ), .Y(n757) );
  INVX2 U279 ( .A(\memory[10][6] ), .Y(n765) );
  INVX2 U280 ( .A(\memory[11][6] ), .Y(n773) );
  INVX2 U281 ( .A(\memory[16][5] ), .Y(n782) );
  INVX2 U282 ( .A(\memory[17][5] ), .Y(n790) );
  INVX2 U283 ( .A(\memory[18][5] ), .Y(n798) );
  INVX2 U284 ( .A(\memory[19][5] ), .Y(n806) );
  INVX2 U285 ( .A(\memory[24][5] ), .Y(n708) );
  INVX2 U286 ( .A(\memory[25][5] ), .Y(n700) );
  INVX2 U287 ( .A(\memory[26][5] ), .Y(n692) );
  INVX2 U288 ( .A(\memory[27][5] ), .Y(n684) );
  INVX2 U289 ( .A(\memory[3][5] ), .Y(n743) );
  INVX2 U290 ( .A(\memory[2][5] ), .Y(n735) );
  INVX2 U291 ( .A(\memory[1][5] ), .Y(n727) );
  INVX2 U292 ( .A(\memory[0][5] ), .Y(n719) );
  INVX2 U293 ( .A(\memory[8][5] ), .Y(n750) );
  INVX2 U294 ( .A(\memory[9][5] ), .Y(n758) );
  INVX2 U295 ( .A(\memory[10][5] ), .Y(n766) );
  INVX2 U296 ( .A(\memory[11][5] ), .Y(n774) );
  INVX2 U297 ( .A(\memory[16][4] ), .Y(n783) );
  INVX2 U298 ( .A(\memory[17][4] ), .Y(n791) );
  INVX2 U299 ( .A(\memory[18][4] ), .Y(n799) );
  INVX2 U300 ( .A(\memory[19][4] ), .Y(n807) );
  INVX2 U301 ( .A(\memory[24][4] ), .Y(n709) );
  INVX2 U302 ( .A(\memory[25][4] ), .Y(n701) );
  INVX2 U303 ( .A(\memory[26][4] ), .Y(n693) );
  INVX2 U304 ( .A(\memory[27][4] ), .Y(n685) );
  INVX2 U305 ( .A(\memory[3][4] ), .Y(n742) );
  INVX2 U306 ( .A(\memory[2][4] ), .Y(n734) );
  INVX2 U307 ( .A(\memory[1][4] ), .Y(n726) );
  INVX2 U308 ( .A(\memory[0][4] ), .Y(n718) );
  INVX2 U309 ( .A(\memory[8][4] ), .Y(n751) );
  INVX2 U310 ( .A(\memory[9][4] ), .Y(n759) );
  INVX2 U311 ( .A(\memory[10][4] ), .Y(n767) );
  INVX2 U312 ( .A(\memory[11][4] ), .Y(n775) );
  INVX2 U313 ( .A(\memory[16][3] ), .Y(n784) );
  INVX2 U314 ( .A(\memory[17][3] ), .Y(n792) );
  INVX2 U315 ( .A(\memory[18][3] ), .Y(n800) );
  INVX2 U316 ( .A(\memory[19][3] ), .Y(n808) );
  INVX2 U317 ( .A(\memory[24][3] ), .Y(n710) );
  INVX2 U318 ( .A(\memory[25][3] ), .Y(n702) );
  INVX2 U319 ( .A(\memory[26][3] ), .Y(n694) );
  INVX2 U320 ( .A(\memory[27][3] ), .Y(n686) );
  INVX2 U321 ( .A(\memory[3][3] ), .Y(n741) );
  INVX2 U322 ( .A(\memory[2][3] ), .Y(n733) );
  INVX2 U323 ( .A(\memory[1][3] ), .Y(n725) );
  INVX2 U324 ( .A(\memory[0][3] ), .Y(n717) );
  INVX2 U325 ( .A(\memory[8][3] ), .Y(n752) );
  INVX2 U326 ( .A(\memory[9][3] ), .Y(n760) );
  INVX2 U327 ( .A(\memory[10][3] ), .Y(n768) );
  INVX2 U328 ( .A(\memory[11][3] ), .Y(n776) );
  INVX2 U329 ( .A(\memory[16][2] ), .Y(n785) );
  INVX2 U330 ( .A(\memory[17][2] ), .Y(n793) );
  INVX2 U331 ( .A(\memory[18][2] ), .Y(n801) );
  INVX2 U332 ( .A(\memory[19][2] ), .Y(n809) );
  INVX2 U333 ( .A(\memory[24][2] ), .Y(n711) );
  INVX2 U334 ( .A(\memory[25][2] ), .Y(n703) );
  INVX2 U335 ( .A(\memory[26][2] ), .Y(n695) );
  INVX2 U336 ( .A(\memory[27][2] ), .Y(n687) );
  INVX2 U337 ( .A(\memory[3][2] ), .Y(n740) );
  INVX2 U338 ( .A(\memory[2][2] ), .Y(n732) );
  INVX2 U339 ( .A(\memory[1][2] ), .Y(n724) );
  INVX2 U340 ( .A(\memory[0][2] ), .Y(n716) );
  INVX2 U341 ( .A(\memory[8][2] ), .Y(n753) );
  INVX2 U342 ( .A(\memory[9][2] ), .Y(n761) );
  INVX2 U343 ( .A(\memory[10][2] ), .Y(n769) );
  INVX2 U344 ( .A(\memory[11][2] ), .Y(n777) );
  INVX2 U345 ( .A(\memory[16][1] ), .Y(n786) );
  INVX2 U346 ( .A(\memory[17][1] ), .Y(n794) );
  INVX2 U347 ( .A(\memory[18][1] ), .Y(n802) );
  INVX2 U348 ( .A(\memory[19][1] ), .Y(n810) );
  INVX2 U349 ( .A(\memory[24][1] ), .Y(n712) );
  INVX2 U350 ( .A(\memory[25][1] ), .Y(n704) );
  INVX2 U351 ( .A(\memory[26][1] ), .Y(n696) );
  INVX2 U352 ( .A(\memory[27][1] ), .Y(n688) );
  INVX2 U353 ( .A(\memory[3][1] ), .Y(n739) );
  INVX2 U354 ( .A(\memory[2][1] ), .Y(n731) );
  INVX2 U355 ( .A(\memory[1][1] ), .Y(n723) );
  INVX2 U356 ( .A(\memory[0][1] ), .Y(n715) );
  INVX2 U357 ( .A(\memory[8][1] ), .Y(n754) );
  INVX2 U358 ( .A(\memory[9][1] ), .Y(n762) );
  INVX2 U359 ( .A(\memory[10][1] ), .Y(n770) );
  INVX2 U360 ( .A(\memory[11][1] ), .Y(n778) );
  INVX2 U361 ( .A(\memory[16][0] ), .Y(n787) );
  INVX2 U362 ( .A(\memory[17][0] ), .Y(n795) );
  INVX2 U363 ( .A(\memory[18][0] ), .Y(n803) );
  INVX2 U364 ( .A(\memory[19][0] ), .Y(n811) );
  INVX2 U365 ( .A(\memory[24][0] ), .Y(n713) );
  INVX2 U366 ( .A(\memory[25][0] ), .Y(n705) );
  INVX2 U367 ( .A(\memory[26][0] ), .Y(n697) );
  INVX2 U368 ( .A(\memory[27][0] ), .Y(n689) );
  INVX2 U369 ( .A(\memory[3][0] ), .Y(n738) );
  INVX2 U370 ( .A(\memory[2][0] ), .Y(n730) );
  INVX2 U371 ( .A(\memory[1][0] ), .Y(n722) );
  INVX2 U372 ( .A(\memory[0][0] ), .Y(n714) );
  INVX2 U373 ( .A(\memory[8][0] ), .Y(n755) );
  INVX2 U374 ( .A(\memory[9][0] ), .Y(n763) );
  INVX2 U375 ( .A(\memory[10][0] ), .Y(n771) );
  INVX2 U376 ( .A(\memory[11][0] ), .Y(n779) );
  INVX2 U377 ( .A(\opcode[16][1] ), .Y(n820) );
  INVX2 U378 ( .A(\opcode[17][1] ), .Y(n822) );
  INVX2 U379 ( .A(\opcode[18][1] ), .Y(n824) );
  INVX2 U380 ( .A(\opcode[19][1] ), .Y(n826) );
  INVX2 U381 ( .A(\opcode[24][1] ), .Y(n672) );
  INVX2 U382 ( .A(\opcode[25][1] ), .Y(n670) );
  INVX2 U383 ( .A(\opcode[26][1] ), .Y(n668) );
  INVX2 U384 ( .A(\opcode[27][1] ), .Y(n666) );
  INVX2 U385 ( .A(\opcode[3][1] ), .Y(n681) );
  INVX2 U386 ( .A(\opcode[2][1] ), .Y(n679) );
  INVX2 U387 ( .A(\opcode[1][1] ), .Y(n677) );
  INVX2 U388 ( .A(\opcode[0][1] ), .Y(n675) );
  INVX2 U389 ( .A(\opcode[8][1] ), .Y(n812) );
  INVX2 U390 ( .A(\opcode[9][1] ), .Y(n814) );
  INVX2 U391 ( .A(\opcode[10][1] ), .Y(n816) );
  INVX2 U392 ( .A(\opcode[11][1] ), .Y(n818) );
  INVX2 U393 ( .A(\opcode[16][0] ), .Y(n821) );
  INVX2 U394 ( .A(\opcode[17][0] ), .Y(n823) );
  INVX2 U395 ( .A(\opcode[18][0] ), .Y(n825) );
  INVX2 U396 ( .A(\opcode[19][0] ), .Y(n827) );
  INVX2 U397 ( .A(n75), .Y(n662) );
  INVX2 U398 ( .A(n153), .Y(n664) );
  INVX2 U399 ( .A(\opcode[24][0] ), .Y(n673) );
  INVX2 U400 ( .A(\opcode[25][0] ), .Y(n671) );
  INVX2 U401 ( .A(\opcode[26][0] ), .Y(n669) );
  INVX2 U402 ( .A(\opcode[27][0] ), .Y(n667) );
  INVX2 U403 ( .A(\opcode[3][0] ), .Y(n680) );
  INVX2 U404 ( .A(\opcode[2][0] ), .Y(n678) );
  INVX2 U405 ( .A(\opcode[1][0] ), .Y(n676) );
  INVX2 U406 ( .A(\opcode[0][0] ), .Y(n674) );
  INVX2 U407 ( .A(n84), .Y(n665) );
  INVX2 U408 ( .A(\opcode[8][0] ), .Y(n813) );
  INVX2 U409 ( .A(\opcode[9][0] ), .Y(n815) );
  INVX2 U410 ( .A(\opcode[10][0] ), .Y(n817) );
  INVX2 U411 ( .A(\opcode[11][0] ), .Y(n819) );
  NAND2X1 U412 ( .A(n75), .B(n82), .Y(n524) );
  NAND2X1 U413 ( .A(n37), .B(n662), .Y(n178) );
  NOR2X1 U414 ( .A(n123), .B(n522), .Y(n180) );
  XNOR2X1 U415 ( .A(n149), .B(n36), .Y(n527) );
  XNOR2X1 U416 ( .A(n94), .B(n153), .Y(n532) );
  XNOR2X1 U417 ( .A(writeptr[4]), .B(n84), .Y(n537) );
  AND2X2 U418 ( .A(n532), .B(n537), .Y(n179) );
  NAND3X1 U419 ( .A(n180), .B(n527), .C(n179), .Y(n181) );
  MUX2X1 U420 ( .B(n181), .A(n747), .S(RST), .Y(n1415) );
  INVX2 U421 ( .A(OUT_OPCODE[0]), .Y(n184) );
  INVX2 U422 ( .A(n1241), .Y(n183) );
  NAND2X1 U423 ( .A(n177), .B(state), .Y(n182) );
  MUX2X1 U424 ( .B(n184), .A(n183), .S(n137), .Y(n1030) );
  INVX2 U425 ( .A(OUT_OPCODE[1]), .Y(n186) );
  INVX2 U426 ( .A(n1214), .Y(n185) );
  MUX2X1 U427 ( .B(n186), .A(n185), .S(n138), .Y(n1031) );
  INVX2 U428 ( .A(DATA[0]), .Y(n188) );
  INVX2 U429 ( .A(n1187), .Y(n187) );
  MUX2X1 U430 ( .B(n188), .A(n187), .S(n137), .Y(n1032) );
  INVX2 U431 ( .A(DATA[1]), .Y(n190) );
  INVX2 U432 ( .A(n1064), .Y(n189) );
  MUX2X1 U433 ( .B(n190), .A(n189), .S(n138), .Y(n1033) );
  INVX2 U434 ( .A(DATA[2]), .Y(n192) );
  INVX2 U435 ( .A(n1025), .Y(n191) );
  MUX2X1 U436 ( .B(n192), .A(n191), .S(n137), .Y(n1034) );
  INVX2 U437 ( .A(DATA[3]), .Y(n194) );
  INVX2 U438 ( .A(n998), .Y(n193) );
  MUX2X1 U439 ( .B(n194), .A(n193), .S(n138), .Y(n1035) );
  INVX2 U440 ( .A(DATA[4]), .Y(n196) );
  INVX2 U441 ( .A(n971), .Y(n195) );
  MUX2X1 U442 ( .B(n196), .A(n195), .S(n137), .Y(n1036) );
  INVX2 U443 ( .A(DATA[5]), .Y(n198) );
  INVX2 U444 ( .A(n944), .Y(n197) );
  MUX2X1 U445 ( .B(n198), .A(n197), .S(n138), .Y(n1037) );
  INVX2 U446 ( .A(DATA[6]), .Y(n200) );
  INVX2 U447 ( .A(n917), .Y(n199) );
  MUX2X1 U448 ( .B(n200), .A(n199), .S(n137), .Y(n1038) );
  INVX2 U449 ( .A(DATA[7]), .Y(n202) );
  INVX2 U450 ( .A(n828), .Y(n201) );
  MUX2X1 U451 ( .B(n202), .A(n201), .S(n138), .Y(n1039) );
  NAND2X1 U452 ( .A(n30), .B(n215), .Y(n347) );
  INVX2 U453 ( .A(n347), .Y(n308) );
  INVX2 U454 ( .A(n54), .Y(n566) );
  NAND2X1 U455 ( .A(n107), .B(n151), .Y(n337) );
  NAND2X1 U456 ( .A(n555), .B(n149), .Y(n203) );
  NAND2X1 U457 ( .A(n337), .B(n203), .Y(n547) );
  NAND2X1 U458 ( .A(n149), .B(n29), .Y(n317) );
  NOR2X1 U459 ( .A(n87), .B(n85), .Y(n205) );
  XNOR2X1 U460 ( .A(n151), .B(n25), .Y(n553) );
  XNOR2X1 U461 ( .A(n553), .B(n594), .Y(n544) );
  NAND3X1 U462 ( .A(n94), .B(n86), .C(n149), .Y(n573) );
  AND2X2 U463 ( .A(n544), .B(n542), .Y(n204) );
  NAND3X1 U464 ( .A(n90), .B(n205), .C(n204), .Y(n277) );
  NAND2X1 U465 ( .A(W_ENABLE), .B(n277), .Y(n558) );
  NAND2X1 U466 ( .A(n566), .B(n581), .Y(n563) );
  NAND2X1 U467 ( .A(n96), .B(n117), .Y(n210) );
  NAND2X1 U468 ( .A(n94), .B(n177), .Y(n298) );
  INVX2 U469 ( .A(n298), .Y(n276) );
  NAND3X1 U470 ( .A(n118), .B(n103), .C(n53), .Y(n206) );
  NAND2X1 U471 ( .A(n239), .B(n569), .Y(n207) );
  MUX2X1 U472 ( .B(\opcode[31][0] ), .A(n171), .S(n365), .Y(n208) );
  NAND2X1 U473 ( .A(n210), .B(n208), .Y(n605) );
  MUX2X1 U474 ( .B(\opcode[31][1] ), .A(n175), .S(n365), .Y(n209) );
  NAND2X1 U475 ( .A(n210), .B(n209), .Y(n604) );
  OR2X2 U476 ( .A(n77), .B(n52), .Y(n556) );
  INVX2 U477 ( .A(n556), .Y(n220) );
  NAND2X1 U478 ( .A(n220), .B(n229), .Y(n565) );
  INVX2 U479 ( .A(n565), .Y(n353) );
  NAND2X1 U480 ( .A(n117), .B(n95), .Y(n214) );
  NAND3X1 U481 ( .A(n149), .B(n77), .C(n82), .Y(n322) );
  INVX2 U482 ( .A(n322), .Y(n283) );
  NAND2X1 U483 ( .A(n239), .B(n283), .Y(n211) );
  MUX2X1 U484 ( .B(\opcode[30][0] ), .A(n171), .S(n374), .Y(n212) );
  NAND2X1 U485 ( .A(n214), .B(n212), .Y(n617) );
  MUX2X1 U486 ( .B(\opcode[30][1] ), .A(n175), .S(n374), .Y(n213) );
  NAND2X1 U487 ( .A(n214), .B(n213), .Y(n616) );
  NAND2X1 U488 ( .A(n98), .B(n118), .Y(n219) );
  NAND3X1 U489 ( .A(n149), .B(n52), .C(n215), .Y(n327) );
  INVX2 U490 ( .A(n327), .Y(n288) );
  NAND2X1 U491 ( .A(n239), .B(n288), .Y(n216) );
  MUX2X1 U492 ( .B(\opcode[29][0] ), .A(n171), .S(n383), .Y(n217) );
  NAND2X1 U493 ( .A(n219), .B(n217), .Y(n633) );
  MUX2X1 U494 ( .B(\opcode[29][1] ), .A(n175), .S(n383), .Y(n218) );
  NAND2X1 U495 ( .A(n219), .B(n218), .Y(n632) );
  NAND2X1 U496 ( .A(n101), .B(n118), .Y(n224) );
  NAND2X1 U497 ( .A(n220), .B(n149), .Y(n332) );
  INVX2 U498 ( .A(n332), .Y(n293) );
  NAND2X1 U499 ( .A(n239), .B(n293), .Y(n221) );
  MUX2X1 U500 ( .B(\opcode[28][0] ), .A(n171), .S(n392), .Y(n222) );
  NAND2X1 U501 ( .A(n224), .B(n222), .Y(n645) );
  MUX2X1 U502 ( .B(\opcode[28][1] ), .A(n175), .S(n392), .Y(n223) );
  NAND2X1 U503 ( .A(n224), .B(n223), .Y(n644) );
  NAND2X1 U504 ( .A(n105), .B(n118), .Y(n228) );
  NAND2X1 U505 ( .A(n239), .B(n471), .Y(n225) );
  MUX2X1 U506 ( .B(\opcode[27][0] ), .A(n171), .S(n394), .Y(n226) );
  NAND2X1 U507 ( .A(n228), .B(n226), .Y(n651) );
  MUX2X1 U508 ( .B(\opcode[27][1] ), .A(n175), .S(n394), .Y(n227) );
  NAND2X1 U509 ( .A(n228), .B(n227), .Y(n650) );
  NAND2X1 U510 ( .A(n100), .B(n118), .Y(n234) );
  NAND3X1 U511 ( .A(n77), .B(n82), .C(n229), .Y(n342) );
  INVX2 U512 ( .A(n342), .Y(n303) );
  NAND2X1 U513 ( .A(n239), .B(n303), .Y(n231) );
  MUX2X1 U514 ( .B(\opcode[26][0] ), .A(n171), .S(n395), .Y(n232) );
  NAND2X1 U515 ( .A(n234), .B(n232), .Y(n631) );
  MUX2X1 U516 ( .B(\opcode[26][1] ), .A(n175), .S(n395), .Y(n233) );
  NAND2X1 U517 ( .A(n234), .B(n233), .Y(n630) );
  NAND2X1 U518 ( .A(n99), .B(n118), .Y(n238) );
  NAND2X1 U519 ( .A(n239), .B(n308), .Y(n235) );
  MUX2X1 U520 ( .B(\opcode[25][0] ), .A(n171), .S(n396), .Y(n236) );
  NAND2X1 U521 ( .A(n238), .B(n236), .Y(n657) );
  MUX2X1 U522 ( .B(\opcode[25][1] ), .A(n175), .S(n396), .Y(n237) );
  NAND2X1 U523 ( .A(n238), .B(n237), .Y(n656) );
  NAND2X1 U524 ( .A(n102), .B(n118), .Y(n242) );
  MUX2X1 U525 ( .B(\opcode[24][0] ), .A(n170), .S(n92), .Y(n240) );
  NAND2X1 U526 ( .A(n242), .B(n240), .Y(n607) );
  MUX2X1 U527 ( .B(\opcode[24][1] ), .A(n174), .S(n92), .Y(n241) );
  NAND2X1 U528 ( .A(n242), .B(n241), .Y(n606) );
  NAND2X1 U529 ( .A(n96), .B(n118), .Y(n247) );
  NAND3X1 U530 ( .A(n122), .B(n53), .C(n103), .Y(n243) );
  NAND2X1 U531 ( .A(n55), .B(n569), .Y(n244) );
  MUX2X1 U532 ( .B(\opcode[23][0] ), .A(n170), .S(n404), .Y(n245) );
  NAND2X1 U533 ( .A(n247), .B(n245), .Y(n619) );
  MUX2X1 U534 ( .B(\opcode[23][1] ), .A(n174), .S(n404), .Y(n246) );
  NAND2X1 U535 ( .A(n247), .B(n246), .Y(n618) );
  NAND2X1 U536 ( .A(n118), .B(n95), .Y(n251) );
  NAND2X1 U537 ( .A(n55), .B(n283), .Y(n248) );
  MUX2X1 U538 ( .B(\opcode[22][0] ), .A(n170), .S(n1), .Y(n249) );
  NAND2X1 U539 ( .A(n251), .B(n249), .Y(n621) );
  MUX2X1 U540 ( .B(\opcode[22][1] ), .A(n174), .S(n1), .Y(n250) );
  NAND2X1 U541 ( .A(n251), .B(n250), .Y(n620) );
  NAND2X1 U542 ( .A(n98), .B(n122), .Y(n255) );
  NAND2X1 U543 ( .A(n271), .B(n288), .Y(n252) );
  MUX2X1 U544 ( .B(\opcode[21][0] ), .A(n170), .S(n421), .Y(n253) );
  NAND2X1 U545 ( .A(n255), .B(n253), .Y(n661) );
  MUX2X1 U546 ( .B(\opcode[21][1] ), .A(n174), .S(n421), .Y(n254) );
  NAND2X1 U547 ( .A(n255), .B(n254), .Y(n660) );
  NAND2X1 U548 ( .A(n101), .B(n122), .Y(n259) );
  NAND2X1 U549 ( .A(n271), .B(n293), .Y(n256) );
  MUX2X1 U550 ( .B(\opcode[20][0] ), .A(n170), .S(n430), .Y(n257) );
  NAND2X1 U551 ( .A(n259), .B(n257), .Y(n659) );
  MUX2X1 U552 ( .B(\opcode[20][1] ), .A(n174), .S(n430), .Y(n258) );
  NAND2X1 U553 ( .A(n259), .B(n258), .Y(n658) );
  NAND2X1 U554 ( .A(n105), .B(n122), .Y(n263) );
  NAND2X1 U555 ( .A(n55), .B(n471), .Y(n260) );
  MUX2X1 U556 ( .B(\opcode[19][0] ), .A(n170), .S(n432), .Y(n261) );
  NAND2X1 U557 ( .A(n263), .B(n261), .Y(n629) );
  MUX2X1 U558 ( .B(\opcode[19][1] ), .A(n174), .S(n432), .Y(n262) );
  NAND2X1 U559 ( .A(n263), .B(n262), .Y(n628) );
  NAND2X1 U560 ( .A(n100), .B(n122), .Y(n267) );
  NAND2X1 U561 ( .A(n271), .B(n303), .Y(n264) );
  MUX2X1 U562 ( .B(\opcode[18][0] ), .A(n170), .S(n433), .Y(n265) );
  NAND2X1 U563 ( .A(n267), .B(n265), .Y(n603) );
  MUX2X1 U564 ( .B(\opcode[18][1] ), .A(n174), .S(n433), .Y(n266) );
  NAND2X1 U565 ( .A(n267), .B(n266), .Y(n602) );
  NAND2X1 U566 ( .A(n99), .B(n122), .Y(n270) );
  MUX2X1 U567 ( .B(\opcode[17][0] ), .A(n170), .S(n73), .Y(n268) );
  NAND2X1 U568 ( .A(n270), .B(n268), .Y(n613) );
  MUX2X1 U569 ( .B(\opcode[17][1] ), .A(n174), .S(n73), .Y(n269) );
  NAND2X1 U570 ( .A(n270), .B(n269), .Y(n612) );
  NAND2X1 U571 ( .A(n102), .B(n122), .Y(n275) );
  NAND2X1 U572 ( .A(n353), .B(n55), .Y(n272) );
  MUX2X1 U573 ( .B(\opcode[16][0] ), .A(n170), .S(n434), .Y(n273) );
  NAND2X1 U574 ( .A(n275), .B(n273), .Y(n627) );
  MUX2X1 U575 ( .B(\opcode[16][1] ), .A(n174), .S(n434), .Y(n274) );
  NAND2X1 U576 ( .A(n275), .B(n274), .Y(n626) );
  NAND2X1 U577 ( .A(n96), .B(n122), .Y(n282) );
  NAND3X1 U578 ( .A(n108), .B(n104), .C(n54), .Y(n278) );
  NAND2X1 U579 ( .A(n472), .B(n569), .Y(n279) );
  MUX2X1 U580 ( .B(\opcode[15][0] ), .A(n170), .S(n442), .Y(n280) );
  NAND2X1 U581 ( .A(n282), .B(n280), .Y(n649) );
  MUX2X1 U582 ( .B(\opcode[15][1] ), .A(n174), .S(n442), .Y(n281) );
  NAND2X1 U583 ( .A(n282), .B(n281), .Y(n648) );
  NAND2X1 U584 ( .A(n122), .B(n95), .Y(n287) );
  NAND2X1 U585 ( .A(n472), .B(n283), .Y(n284) );
  MUX2X1 U586 ( .B(\opcode[14][0] ), .A(n170), .S(n451), .Y(n285) );
  NAND2X1 U587 ( .A(n287), .B(n285), .Y(n637) );
  MUX2X1 U588 ( .B(\opcode[14][1] ), .A(n174), .S(n451), .Y(n286) );
  NAND2X1 U589 ( .A(n287), .B(n286), .Y(n636) );
  NAND2X1 U590 ( .A(n98), .B(n108), .Y(n292) );
  NAND2X1 U591 ( .A(n472), .B(n288), .Y(n289) );
  MUX2X1 U592 ( .B(\opcode[13][0] ), .A(n170), .S(n460), .Y(n290) );
  NAND2X1 U593 ( .A(n292), .B(n290), .Y(n639) );
  MUX2X1 U594 ( .B(\opcode[13][1] ), .A(n174), .S(n460), .Y(n291) );
  NAND2X1 U595 ( .A(n292), .B(n291), .Y(n638) );
  NAND2X1 U596 ( .A(n101), .B(n108), .Y(n297) );
  NAND2X1 U597 ( .A(n472), .B(n293), .Y(n294) );
  MUX2X1 U598 ( .B(\opcode[12][0] ), .A(n171), .S(n469), .Y(n295) );
  NAND2X1 U599 ( .A(n297), .B(n295), .Y(n643) );
  MUX2X1 U600 ( .B(\opcode[12][1] ), .A(n173), .S(n469), .Y(n296) );
  NAND2X1 U601 ( .A(n297), .B(n296), .Y(n642) );
  MUX2X1 U602 ( .B(n83), .A(n327), .S(n566), .Y(n300) );
  NOR2X1 U603 ( .A(n558), .B(n298), .Y(n299) );
  NAND3X1 U604 ( .A(n300), .B(n574), .C(n299), .Y(n301) );
  INVX2 U605 ( .A(n301), .Y(n302) );
  MUX2X1 U606 ( .B(n819), .A(n172), .S(n302), .Y(n1056) );
  MUX2X1 U607 ( .B(n818), .A(n176), .S(n302), .Y(n1057) );
  NAND2X1 U608 ( .A(n100), .B(n108), .Y(n307) );
  NAND2X1 U609 ( .A(n472), .B(n303), .Y(n304) );
  MUX2X1 U610 ( .B(\opcode[10][0] ), .A(n170), .S(n473), .Y(n305) );
  NAND2X1 U611 ( .A(n307), .B(n305), .Y(n647) );
  MUX2X1 U612 ( .B(\opcode[10][1] ), .A(n173), .S(n473), .Y(n306) );
  NAND2X1 U613 ( .A(n307), .B(n306), .Y(n646) );
  NAND2X1 U614 ( .A(n99), .B(n108), .Y(n312) );
  NAND2X1 U615 ( .A(n472), .B(n308), .Y(n309) );
  MUX2X1 U616 ( .B(\opcode[9][0] ), .A(n170), .S(n474), .Y(n310) );
  NAND2X1 U617 ( .A(n312), .B(n310), .Y(n623) );
  MUX2X1 U618 ( .B(\opcode[9][1] ), .A(n173), .S(n474), .Y(n311) );
  NAND2X1 U619 ( .A(n312), .B(n311), .Y(n622) );
  NAND2X1 U620 ( .A(n102), .B(n108), .Y(n316) );
  NAND2X1 U621 ( .A(n472), .B(n353), .Y(n313) );
  MUX2X1 U622 ( .B(\opcode[8][0] ), .A(n170), .S(n475), .Y(n314) );
  NAND2X1 U623 ( .A(n316), .B(n314), .Y(n635) );
  MUX2X1 U624 ( .B(\opcode[8][1] ), .A(n173), .S(n475), .Y(n315) );
  NAND2X1 U625 ( .A(n316), .B(n315), .Y(n634) );
  NAND2X1 U626 ( .A(n96), .B(n108), .Y(n321) );
  NAND3X1 U627 ( .A(n53), .B(n117), .C(n104), .Y(n352) );
  OR2X2 U628 ( .A(n126), .B(n78), .Y(n318) );
  MUX2X1 U629 ( .B(\opcode[7][0] ), .A(n170), .S(n483), .Y(n319) );
  NAND2X1 U630 ( .A(n321), .B(n319), .Y(n609) );
  MUX2X1 U631 ( .B(\opcode[7][1] ), .A(n173), .S(n483), .Y(n320) );
  NAND2X1 U632 ( .A(n321), .B(n320), .Y(n608) );
  NAND2X1 U633 ( .A(n108), .B(n95), .Y(n326) );
  OR2X2 U634 ( .A(n125), .B(n322), .Y(n323) );
  NAND2X1 U635 ( .A(n326), .B(n324), .Y(n601) );
  MUX2X1 U636 ( .B(\opcode[6][1] ), .A(n173), .S(n492), .Y(n325) );
  NAND2X1 U637 ( .A(n326), .B(n325), .Y(n600) );
  NAND2X1 U638 ( .A(n98), .B(n117), .Y(n331) );
  OR2X2 U639 ( .A(n125), .B(n327), .Y(n328) );
  MUX2X1 U640 ( .B(\opcode[5][0] ), .A(n170), .S(n501), .Y(n329) );
  NAND2X1 U641 ( .A(n331), .B(n329), .Y(n615) );
  MUX2X1 U642 ( .B(\opcode[5][1] ), .A(n173), .S(n501), .Y(n330) );
  NAND2X1 U643 ( .A(n331), .B(n330), .Y(n614) );
  NAND2X1 U644 ( .A(n101), .B(n117), .Y(n336) );
  OR2X2 U645 ( .A(n126), .B(n332), .Y(n333) );
  MUX2X1 U646 ( .B(\opcode[4][0] ), .A(n171), .S(n510), .Y(n334) );
  NAND2X1 U647 ( .A(n336), .B(n334), .Y(n641) );
  MUX2X1 U648 ( .B(\opcode[4][1] ), .A(n173), .S(n510), .Y(n335) );
  NAND2X1 U649 ( .A(n336), .B(n335), .Y(n640) );
  NAND2X1 U650 ( .A(n105), .B(n117), .Y(n341) );
  OR2X2 U651 ( .A(n126), .B(n83), .Y(n338) );
  MUX2X1 U652 ( .B(\opcode[3][0] ), .A(n170), .S(n512), .Y(n339) );
  NAND2X1 U653 ( .A(n341), .B(n339), .Y(n625) );
  MUX2X1 U654 ( .B(\opcode[3][1] ), .A(n173), .S(n512), .Y(n340) );
  NAND2X1 U655 ( .A(n341), .B(n340), .Y(n624) );
  NAND2X1 U656 ( .A(n100), .B(n117), .Y(n346) );
  OR2X2 U657 ( .A(n126), .B(n342), .Y(n343) );
  NAND2X1 U658 ( .A(n346), .B(n344), .Y(n655) );
  MUX2X1 U659 ( .B(\opcode[2][1] ), .A(n173), .S(n513), .Y(n345) );
  NAND2X1 U660 ( .A(n346), .B(n345), .Y(n654) );
  NAND2X1 U661 ( .A(n99), .B(n117), .Y(n351) );
  OR2X2 U662 ( .A(n126), .B(n347), .Y(n348) );
  MUX2X1 U663 ( .B(\opcode[1][0] ), .A(n170), .S(n514), .Y(n349) );
  NAND2X1 U664 ( .A(n351), .B(n349), .Y(n653) );
  MUX2X1 U665 ( .B(\opcode[1][1] ), .A(n173), .S(n514), .Y(n350) );
  NAND2X1 U666 ( .A(n351), .B(n350), .Y(n652) );
  NAND2X1 U667 ( .A(n102), .B(n117), .Y(n357) );
  INVX2 U668 ( .A(n125), .Y(n354) );
  MUX2X1 U669 ( .B(\opcode[0][0] ), .A(n170), .S(n69), .Y(n355) );
  NAND2X1 U670 ( .A(n357), .B(n355), .Y(n611) );
  MUX2X1 U671 ( .B(\opcode[0][1] ), .A(n173), .S(n69), .Y(n356) );
  NAND2X1 U672 ( .A(n357), .B(n356), .Y(n610) );
  INVX2 U673 ( .A(\memory[31][0] ), .Y(n358) );
  MUX2X1 U674 ( .B(n358), .A(n154), .S(n64), .Y(n1072) );
  INVX2 U675 ( .A(\memory[31][1] ), .Y(n359) );
  MUX2X1 U676 ( .B(n359), .A(n156), .S(n64), .Y(n1073) );
  INVX2 U677 ( .A(\memory[31][2] ), .Y(n360) );
  MUX2X1 U678 ( .B(n360), .A(n158), .S(n64), .Y(n1074) );
  INVX2 U679 ( .A(\memory[31][3] ), .Y(n361) );
  MUX2X1 U680 ( .B(n361), .A(n160), .S(n365), .Y(n1075) );
  INVX2 U681 ( .A(\memory[31][4] ), .Y(n362) );
  MUX2X1 U682 ( .B(n362), .A(n162), .S(n64), .Y(n1076) );
  INVX2 U683 ( .A(\memory[31][5] ), .Y(n363) );
  MUX2X1 U684 ( .B(n363), .A(n164), .S(n365), .Y(n1077) );
  INVX2 U685 ( .A(\memory[31][6] ), .Y(n364) );
  MUX2X1 U686 ( .B(n364), .A(n166), .S(n64), .Y(n1078) );
  INVX2 U687 ( .A(\memory[31][7] ), .Y(n366) );
  MUX2X1 U688 ( .B(n366), .A(n168), .S(n64), .Y(n1079) );
  INVX2 U689 ( .A(\memory[30][0] ), .Y(n367) );
  MUX2X1 U690 ( .B(n367), .A(n154), .S(n63), .Y(n1080) );
  INVX2 U691 ( .A(\memory[30][1] ), .Y(n368) );
  MUX2X1 U692 ( .B(n368), .A(n156), .S(n374), .Y(n1081) );
  INVX2 U693 ( .A(\memory[30][2] ), .Y(n369) );
  MUX2X1 U694 ( .B(n369), .A(n158), .S(n374), .Y(n1082) );
  INVX2 U695 ( .A(\memory[30][3] ), .Y(n370) );
  MUX2X1 U696 ( .B(n370), .A(n160), .S(n374), .Y(n1083) );
  INVX2 U697 ( .A(\memory[30][4] ), .Y(n371) );
  MUX2X1 U698 ( .B(n371), .A(n162), .S(n374), .Y(n1084) );
  INVX2 U699 ( .A(\memory[30][5] ), .Y(n372) );
  MUX2X1 U700 ( .B(n372), .A(n164), .S(n374), .Y(n1085) );
  INVX2 U701 ( .A(\memory[30][6] ), .Y(n373) );
  MUX2X1 U702 ( .B(n373), .A(n166), .S(n374), .Y(n1086) );
  INVX2 U703 ( .A(\memory[30][7] ), .Y(n375) );
  MUX2X1 U704 ( .B(n375), .A(n168), .S(n63), .Y(n1087) );
  INVX2 U705 ( .A(\memory[29][0] ), .Y(n376) );
  MUX2X1 U706 ( .B(n376), .A(n154), .S(n62), .Y(n1088) );
  INVX2 U707 ( .A(\memory[29][1] ), .Y(n377) );
  MUX2X1 U708 ( .B(n377), .A(n156), .S(n383), .Y(n1089) );
  INVX2 U709 ( .A(\memory[29][2] ), .Y(n378) );
  MUX2X1 U710 ( .B(n378), .A(n158), .S(n383), .Y(n1090) );
  INVX2 U711 ( .A(\memory[29][3] ), .Y(n379) );
  MUX2X1 U712 ( .B(n379), .A(n160), .S(n383), .Y(n1091) );
  INVX2 U713 ( .A(\memory[29][4] ), .Y(n380) );
  MUX2X1 U714 ( .B(n380), .A(n162), .S(n383), .Y(n1092) );
  INVX2 U715 ( .A(\memory[29][5] ), .Y(n381) );
  MUX2X1 U716 ( .B(n381), .A(n164), .S(n383), .Y(n1093) );
  INVX2 U717 ( .A(\memory[29][6] ), .Y(n382) );
  MUX2X1 U718 ( .B(n382), .A(n166), .S(n383), .Y(n1094) );
  INVX2 U719 ( .A(\memory[29][7] ), .Y(n384) );
  MUX2X1 U720 ( .B(n384), .A(n168), .S(n62), .Y(n1095) );
  INVX2 U721 ( .A(\memory[28][0] ), .Y(n385) );
  MUX2X1 U722 ( .B(n385), .A(n154), .S(n61), .Y(n1096) );
  INVX2 U723 ( .A(\memory[28][1] ), .Y(n386) );
  MUX2X1 U724 ( .B(n386), .A(n156), .S(n392), .Y(n1097) );
  INVX2 U725 ( .A(\memory[28][2] ), .Y(n387) );
  MUX2X1 U726 ( .B(n387), .A(n158), .S(n392), .Y(n1098) );
  INVX2 U727 ( .A(\memory[28][3] ), .Y(n388) );
  MUX2X1 U728 ( .B(n388), .A(n160), .S(n392), .Y(n1099) );
  INVX2 U729 ( .A(\memory[28][4] ), .Y(n389) );
  MUX2X1 U730 ( .B(n389), .A(n162), .S(n392), .Y(n1100) );
  INVX2 U731 ( .A(\memory[28][5] ), .Y(n390) );
  MUX2X1 U732 ( .B(n390), .A(n164), .S(n392), .Y(n1101) );
  INVX2 U733 ( .A(\memory[28][6] ), .Y(n391) );
  MUX2X1 U734 ( .B(n391), .A(n166), .S(n392), .Y(n1102) );
  INVX2 U735 ( .A(\memory[28][7] ), .Y(n393) );
  MUX2X1 U736 ( .B(n393), .A(n168), .S(n61), .Y(n1103) );
  MUX2X1 U737 ( .B(n689), .A(n154), .S(n24), .Y(n1293) );
  MUX2X1 U738 ( .B(n688), .A(n156), .S(n394), .Y(n1292) );
  MUX2X1 U739 ( .B(n687), .A(n158), .S(n24), .Y(n1291) );
  MUX2X1 U740 ( .B(n686), .A(n160), .S(n24), .Y(n1290) );
  MUX2X1 U741 ( .B(n685), .A(n162), .S(n394), .Y(n1289) );
  MUX2X1 U742 ( .B(n684), .A(n164), .S(n24), .Y(n1288) );
  MUX2X1 U743 ( .B(n683), .A(n166), .S(n24), .Y(n1287) );
  MUX2X1 U744 ( .B(n682), .A(n168), .S(n24), .Y(n1286) );
  MUX2X1 U745 ( .B(n697), .A(n154), .S(n60), .Y(n1301) );
  MUX2X1 U746 ( .B(n696), .A(n156), .S(n395), .Y(n1300) );
  MUX2X1 U747 ( .B(n695), .A(n158), .S(n395), .Y(n1299) );
  MUX2X1 U748 ( .B(n694), .A(n160), .S(n395), .Y(n1298) );
  MUX2X1 U749 ( .B(n693), .A(n162), .S(n395), .Y(n1297) );
  MUX2X1 U750 ( .B(n692), .A(n164), .S(n395), .Y(n1296) );
  MUX2X1 U751 ( .B(n691), .A(n166), .S(n395), .Y(n1295) );
  MUX2X1 U752 ( .B(n690), .A(n168), .S(n60), .Y(n1294) );
  MUX2X1 U753 ( .B(n705), .A(n154), .S(n59), .Y(n1309) );
  MUX2X1 U754 ( .B(n704), .A(n156), .S(n396), .Y(n1308) );
  MUX2X1 U755 ( .B(n703), .A(n158), .S(n396), .Y(n1307) );
  MUX2X1 U756 ( .B(n702), .A(n160), .S(n396), .Y(n1306) );
  MUX2X1 U757 ( .B(n701), .A(n162), .S(n396), .Y(n1305) );
  MUX2X1 U758 ( .B(n700), .A(n164), .S(n396), .Y(n1304) );
  MUX2X1 U759 ( .B(n699), .A(n166), .S(n396), .Y(n1303) );
  MUX2X1 U760 ( .B(n698), .A(n168), .S(n59), .Y(n1302) );
  MUX2X1 U761 ( .B(n713), .A(n154), .S(n93), .Y(n1317) );
  MUX2X1 U762 ( .B(n712), .A(n156), .S(n93), .Y(n1316) );
  MUX2X1 U763 ( .B(n711), .A(n158), .S(n93), .Y(n1315) );
  MUX2X1 U764 ( .B(n710), .A(n160), .S(n93), .Y(n1314) );
  MUX2X1 U765 ( .B(n709), .A(n162), .S(n93), .Y(n1313) );
  MUX2X1 U766 ( .B(n708), .A(n164), .S(n93), .Y(n1312) );
  MUX2X1 U767 ( .B(n707), .A(n166), .S(n93), .Y(n1311) );
  MUX2X1 U768 ( .B(n706), .A(n168), .S(n92), .Y(n1310) );
  INVX2 U769 ( .A(\memory[23][0] ), .Y(n397) );
  MUX2X1 U770 ( .B(n397), .A(n154), .S(n34), .Y(n1325) );
  INVX2 U771 ( .A(\memory[23][1] ), .Y(n398) );
  MUX2X1 U772 ( .B(n398), .A(n156), .S(n34), .Y(n1324) );
  INVX2 U773 ( .A(\memory[23][2] ), .Y(n399) );
  MUX2X1 U774 ( .B(n399), .A(n158), .S(n34), .Y(n1323) );
  INVX2 U775 ( .A(\memory[23][3] ), .Y(n400) );
  MUX2X1 U776 ( .B(n400), .A(n160), .S(n404), .Y(n1322) );
  INVX2 U777 ( .A(\memory[23][4] ), .Y(n401) );
  MUX2X1 U778 ( .B(n401), .A(n162), .S(n34), .Y(n1321) );
  INVX2 U779 ( .A(\memory[23][5] ), .Y(n402) );
  MUX2X1 U780 ( .B(n402), .A(n164), .S(n404), .Y(n1320) );
  INVX2 U781 ( .A(\memory[23][6] ), .Y(n403) );
  MUX2X1 U782 ( .B(n403), .A(n166), .S(n34), .Y(n1319) );
  INVX2 U783 ( .A(\memory[23][7] ), .Y(n405) );
  MUX2X1 U784 ( .B(n405), .A(n168), .S(n34), .Y(n1318) );
  INVX2 U785 ( .A(\memory[22][0] ), .Y(n406) );
  MUX2X1 U786 ( .B(n406), .A(n154), .S(n33), .Y(n1333) );
  INVX2 U787 ( .A(\memory[22][1] ), .Y(n407) );
  MUX2X1 U788 ( .B(n407), .A(n156), .S(n1), .Y(n1332) );
  INVX2 U789 ( .A(\memory[22][2] ), .Y(n408) );
  MUX2X1 U790 ( .B(n408), .A(n158), .S(n33), .Y(n1331) );
  INVX2 U791 ( .A(\memory[22][3] ), .Y(n409) );
  MUX2X1 U792 ( .B(n409), .A(n160), .S(n33), .Y(n1330) );
  INVX2 U793 ( .A(\memory[22][4] ), .Y(n410) );
  MUX2X1 U794 ( .B(n410), .A(n162), .S(n1), .Y(n1329) );
  INVX2 U795 ( .A(\memory[22][5] ), .Y(n411) );
  MUX2X1 U796 ( .B(n411), .A(n164), .S(n33), .Y(n1328) );
  INVX2 U797 ( .A(\memory[22][6] ), .Y(n412) );
  MUX2X1 U798 ( .B(n412), .A(n166), .S(n33), .Y(n1327) );
  INVX2 U799 ( .A(\memory[22][7] ), .Y(n413) );
  MUX2X1 U800 ( .B(n413), .A(n168), .S(n33), .Y(n1326) );
  INVX2 U801 ( .A(\memory[21][0] ), .Y(n414) );
  MUX2X1 U802 ( .B(n414), .A(n154), .S(n45), .Y(n1341) );
  INVX2 U803 ( .A(\memory[21][1] ), .Y(n415) );
  MUX2X1 U804 ( .B(n415), .A(n156), .S(n46), .Y(n1340) );
  INVX2 U805 ( .A(\memory[21][2] ), .Y(n416) );
  MUX2X1 U806 ( .B(n416), .A(n158), .S(n45), .Y(n1339) );
  INVX2 U807 ( .A(\memory[21][3] ), .Y(n417) );
  MUX2X1 U808 ( .B(n417), .A(n160), .S(n46), .Y(n1338) );
  INVX2 U809 ( .A(\memory[21][4] ), .Y(n418) );
  MUX2X1 U810 ( .B(n418), .A(n162), .S(n45), .Y(n1337) );
  INVX2 U811 ( .A(\memory[21][5] ), .Y(n419) );
  MUX2X1 U812 ( .B(n419), .A(n164), .S(n46), .Y(n1336) );
  INVX2 U813 ( .A(\memory[21][6] ), .Y(n420) );
  MUX2X1 U814 ( .B(n420), .A(n166), .S(n45), .Y(n1335) );
  INVX2 U815 ( .A(\memory[21][7] ), .Y(n422) );
  MUX2X1 U816 ( .B(n422), .A(n168), .S(n46), .Y(n1334) );
  INVX2 U817 ( .A(\memory[20][0] ), .Y(n423) );
  MUX2X1 U818 ( .B(n423), .A(n154), .S(n44), .Y(n1349) );
  INVX2 U819 ( .A(\memory[20][1] ), .Y(n424) );
  MUX2X1 U820 ( .B(n424), .A(n156), .S(n430), .Y(n1348) );
  INVX2 U821 ( .A(\memory[20][2] ), .Y(n425) );
  MUX2X1 U822 ( .B(n425), .A(n158), .S(n44), .Y(n1347) );
  INVX2 U823 ( .A(\memory[20][3] ), .Y(n426) );
  MUX2X1 U824 ( .B(n426), .A(n160), .S(n44), .Y(n1346) );
  INVX2 U825 ( .A(\memory[20][4] ), .Y(n427) );
  MUX2X1 U826 ( .B(n427), .A(n162), .S(n44), .Y(n1345) );
  INVX2 U827 ( .A(\memory[20][5] ), .Y(n428) );
  MUX2X1 U828 ( .B(n428), .A(n164), .S(n44), .Y(n1344) );
  INVX2 U829 ( .A(\memory[20][6] ), .Y(n429) );
  MUX2X1 U830 ( .B(n429), .A(n166), .S(n44), .Y(n1343) );
  INVX2 U831 ( .A(\memory[20][7] ), .Y(n431) );
  MUX2X1 U832 ( .B(n431), .A(n168), .S(n430), .Y(n1342) );
  MUX2X1 U833 ( .B(n811), .A(n154), .S(n56), .Y(n1104) );
  MUX2X1 U834 ( .B(n810), .A(n156), .S(n56), .Y(n1105) );
  MUX2X1 U835 ( .B(n809), .A(n159), .S(n56), .Y(n1106) );
  MUX2X1 U836 ( .B(n808), .A(n160), .S(n432), .Y(n1107) );
  MUX2X1 U837 ( .B(n807), .A(n162), .S(n56), .Y(n1108) );
  MUX2X1 U838 ( .B(n806), .A(n164), .S(n432), .Y(n1109) );
  MUX2X1 U839 ( .B(n805), .A(n166), .S(n56), .Y(n1110) );
  MUX2X1 U840 ( .B(n804), .A(n168), .S(n56), .Y(n1111) );
  MUX2X1 U841 ( .B(n803), .A(n154), .S(n42), .Y(n1112) );
  MUX2X1 U842 ( .B(n802), .A(n156), .S(n43), .Y(n1113) );
  MUX2X1 U843 ( .B(n801), .A(n159), .S(n42), .Y(n1114) );
  MUX2X1 U844 ( .B(n800), .A(n160), .S(n43), .Y(n1115) );
  MUX2X1 U845 ( .B(n799), .A(n162), .S(n42), .Y(n1116) );
  MUX2X1 U846 ( .B(n798), .A(n164), .S(n43), .Y(n1117) );
  MUX2X1 U847 ( .B(n797), .A(n166), .S(n42), .Y(n1118) );
  MUX2X1 U848 ( .B(n796), .A(n168), .S(n43), .Y(n1119) );
  MUX2X1 U849 ( .B(n795), .A(n154), .S(n73), .Y(n1120) );
  MUX2X1 U850 ( .B(n794), .A(n156), .S(n73), .Y(n1121) );
  MUX2X1 U851 ( .B(n793), .A(n159), .S(n32), .Y(n1122) );
  MUX2X1 U852 ( .B(n792), .A(n160), .S(n32), .Y(n1123) );
  MUX2X1 U853 ( .B(n791), .A(n162), .S(n32), .Y(n1124) );
  MUX2X1 U854 ( .B(n790), .A(n164), .S(n73), .Y(n1125) );
  MUX2X1 U855 ( .B(n789), .A(n166), .S(n32), .Y(n1126) );
  MUX2X1 U856 ( .B(n788), .A(n168), .S(n73), .Y(n1127) );
  MUX2X1 U857 ( .B(n787), .A(n154), .S(n31), .Y(n1128) );
  MUX2X1 U858 ( .B(n786), .A(n156), .S(n31), .Y(n1129) );
  MUX2X1 U859 ( .B(n785), .A(n159), .S(n31), .Y(n1130) );
  MUX2X1 U860 ( .B(n784), .A(n160), .S(n434), .Y(n1131) );
  MUX2X1 U861 ( .B(n783), .A(n162), .S(n31), .Y(n1132) );
  MUX2X1 U862 ( .B(n782), .A(n164), .S(n434), .Y(n1133) );
  MUX2X1 U863 ( .B(n781), .A(n166), .S(n31), .Y(n1134) );
  MUX2X1 U864 ( .B(n780), .A(n168), .S(n31), .Y(n1135) );
  INVX2 U865 ( .A(\memory[15][0] ), .Y(n435) );
  MUX2X1 U866 ( .B(n435), .A(n154), .S(n67), .Y(n1357) );
  INVX2 U867 ( .A(\memory[15][1] ), .Y(n436) );
  MUX2X1 U868 ( .B(n436), .A(n156), .S(n67), .Y(n1356) );
  INVX2 U869 ( .A(\memory[15][2] ), .Y(n437) );
  MUX2X1 U870 ( .B(n437), .A(n159), .S(n67), .Y(n1355) );
  INVX2 U871 ( .A(\memory[15][3] ), .Y(n438) );
  MUX2X1 U872 ( .B(n438), .A(n160), .S(n442), .Y(n1354) );
  INVX2 U873 ( .A(\memory[15][4] ), .Y(n439) );
  MUX2X1 U874 ( .B(n439), .A(n162), .S(n67), .Y(n1353) );
  INVX2 U875 ( .A(\memory[15][5] ), .Y(n440) );
  MUX2X1 U876 ( .B(n440), .A(n164), .S(n442), .Y(n1352) );
  INVX2 U877 ( .A(\memory[15][6] ), .Y(n441) );
  MUX2X1 U878 ( .B(n441), .A(n166), .S(n67), .Y(n1351) );
  INVX2 U879 ( .A(\memory[15][7] ), .Y(n443) );
  MUX2X1 U880 ( .B(n443), .A(n168), .S(n67), .Y(n1350) );
  INVX2 U881 ( .A(\memory[14][0] ), .Y(n444) );
  MUX2X1 U882 ( .B(n444), .A(n154), .S(n65), .Y(n1365) );
  INVX2 U883 ( .A(\memory[14][1] ), .Y(n445) );
  MUX2X1 U884 ( .B(n445), .A(n156), .S(n451), .Y(n1364) );
  INVX2 U885 ( .A(\memory[14][2] ), .Y(n446) );
  MUX2X1 U886 ( .B(n446), .A(n159), .S(n65), .Y(n1363) );
  INVX2 U887 ( .A(\memory[14][3] ), .Y(n447) );
  MUX2X1 U888 ( .B(n447), .A(n160), .S(n65), .Y(n1362) );
  INVX2 U889 ( .A(\memory[14][4] ), .Y(n448) );
  MUX2X1 U890 ( .B(n448), .A(n518), .S(n65), .Y(n1361) );
  INVX2 U891 ( .A(\memory[14][5] ), .Y(n449) );
  MUX2X1 U892 ( .B(n449), .A(n164), .S(n65), .Y(n1360) );
  INVX2 U893 ( .A(\memory[14][6] ), .Y(n450) );
  MUX2X1 U894 ( .B(n450), .A(n520), .S(n65), .Y(n1359) );
  INVX2 U895 ( .A(\memory[14][7] ), .Y(n452) );
  MUX2X1 U896 ( .B(n452), .A(n521), .S(n65), .Y(n1358) );
  INVX2 U897 ( .A(\memory[13][0] ), .Y(n453) );
  MUX2X1 U898 ( .B(n453), .A(n154), .S(n460), .Y(n1373) );
  INVX2 U899 ( .A(\memory[13][1] ), .Y(n454) );
  MUX2X1 U900 ( .B(n454), .A(n156), .S(n460), .Y(n1372) );
  INVX2 U901 ( .A(\memory[13][2] ), .Y(n455) );
  MUX2X1 U902 ( .B(n455), .A(n159), .S(n460), .Y(n1371) );
  INVX2 U903 ( .A(\memory[13][3] ), .Y(n456) );
  MUX2X1 U904 ( .B(n456), .A(n160), .S(n460), .Y(n1370) );
  INVX2 U905 ( .A(\memory[13][4] ), .Y(n457) );
  MUX2X1 U906 ( .B(n457), .A(n518), .S(n460), .Y(n1369) );
  INVX2 U907 ( .A(\memory[13][5] ), .Y(n458) );
  MUX2X1 U908 ( .B(n458), .A(n164), .S(n460), .Y(n1368) );
  INVX2 U909 ( .A(\memory[13][6] ), .Y(n459) );
  MUX2X1 U910 ( .B(n459), .A(n520), .S(n460), .Y(n1367) );
  INVX2 U911 ( .A(\memory[13][7] ), .Y(n461) );
  MUX2X1 U912 ( .B(n461), .A(n521), .S(n460), .Y(n1366) );
  INVX2 U913 ( .A(\memory[12][0] ), .Y(n462) );
  MUX2X1 U914 ( .B(n462), .A(n515), .S(n469), .Y(n1381) );
  INVX2 U915 ( .A(\memory[12][1] ), .Y(n463) );
  MUX2X1 U916 ( .B(n463), .A(n516), .S(n469), .Y(n1380) );
  INVX2 U917 ( .A(\memory[12][2] ), .Y(n464) );
  MUX2X1 U918 ( .B(n464), .A(n159), .S(n469), .Y(n1379) );
  INVX2 U919 ( .A(\memory[12][3] ), .Y(n465) );
  MUX2X1 U920 ( .B(n465), .A(n517), .S(n469), .Y(n1378) );
  INVX2 U921 ( .A(\memory[12][4] ), .Y(n466) );
  MUX2X1 U922 ( .B(n466), .A(n518), .S(n469), .Y(n1377) );
  INVX2 U923 ( .A(\memory[12][5] ), .Y(n467) );
  MUX2X1 U924 ( .B(n467), .A(n519), .S(n469), .Y(n1376) );
  INVX2 U925 ( .A(\memory[12][6] ), .Y(n468) );
  MUX2X1 U926 ( .B(n468), .A(n520), .S(n469), .Y(n1375) );
  INVX2 U927 ( .A(\memory[12][7] ), .Y(n470) );
  MUX2X1 U928 ( .B(n470), .A(n521), .S(n469), .Y(n1374) );
  MUX2X1 U929 ( .B(n779), .A(n515), .S(n97), .Y(n1136) );
  MUX2X1 U930 ( .B(n778), .A(n516), .S(n97), .Y(n1137) );
  MUX2X1 U931 ( .B(n777), .A(n159), .S(n97), .Y(n1138) );
  MUX2X1 U932 ( .B(n776), .A(n517), .S(n97), .Y(n1139) );
  MUX2X1 U933 ( .B(n775), .A(n518), .S(n97), .Y(n1140) );
  MUX2X1 U934 ( .B(n774), .A(n519), .S(n97), .Y(n1141) );
  MUX2X1 U935 ( .B(n773), .A(n520), .S(n97), .Y(n1142) );
  MUX2X1 U936 ( .B(n772), .A(n521), .S(n97), .Y(n1143) );
  MUX2X1 U937 ( .B(n771), .A(n515), .S(n473), .Y(n1144) );
  MUX2X1 U938 ( .B(n770), .A(n516), .S(n473), .Y(n1145) );
  MUX2X1 U939 ( .B(n769), .A(n159), .S(n473), .Y(n1146) );
  MUX2X1 U940 ( .B(n768), .A(n517), .S(n473), .Y(n1147) );
  MUX2X1 U941 ( .B(n767), .A(n518), .S(n473), .Y(n1148) );
  MUX2X1 U942 ( .B(n766), .A(n519), .S(n473), .Y(n1149) );
  MUX2X1 U943 ( .B(n765), .A(n520), .S(n473), .Y(n1150) );
  MUX2X1 U944 ( .B(n764), .A(n521), .S(n473), .Y(n1151) );
  MUX2X1 U945 ( .B(n763), .A(n154), .S(n474), .Y(n1152) );
  MUX2X1 U946 ( .B(n762), .A(n156), .S(n474), .Y(n1153) );
  MUX2X1 U947 ( .B(n761), .A(n159), .S(n474), .Y(n1154) );
  MUX2X1 U948 ( .B(n760), .A(n160), .S(n474), .Y(n1155) );
  MUX2X1 U949 ( .B(n759), .A(n518), .S(n474), .Y(n1156) );
  MUX2X1 U950 ( .B(n758), .A(n164), .S(n474), .Y(n1157) );
  MUX2X1 U951 ( .B(n757), .A(n520), .S(n474), .Y(n1158) );
  MUX2X1 U952 ( .B(n756), .A(n521), .S(n474), .Y(n1159) );
  MUX2X1 U953 ( .B(n755), .A(n154), .S(n475), .Y(n1160) );
  MUX2X1 U954 ( .B(n754), .A(n156), .S(n475), .Y(n1161) );
  MUX2X1 U955 ( .B(n753), .A(n159), .S(n475), .Y(n1162) );
  MUX2X1 U956 ( .B(n752), .A(n160), .S(n475), .Y(n1163) );
  MUX2X1 U957 ( .B(n751), .A(n518), .S(n475), .Y(n1164) );
  MUX2X1 U958 ( .B(n750), .A(n164), .S(n475), .Y(n1165) );
  MUX2X1 U959 ( .B(n749), .A(n520), .S(n475), .Y(n1166) );
  MUX2X1 U960 ( .B(n748), .A(n521), .S(n475), .Y(n1167) );
  INVX2 U961 ( .A(\memory[7][0] ), .Y(n476) );
  MUX2X1 U962 ( .B(n476), .A(n515), .S(n127), .Y(n906) );
  INVX2 U963 ( .A(\memory[7][1] ), .Y(n477) );
  MUX2X1 U964 ( .B(n477), .A(n516), .S(n127), .Y(n905) );
  INVX2 U965 ( .A(\memory[7][2] ), .Y(n478) );
  MUX2X1 U966 ( .B(n478), .A(n159), .S(n127), .Y(n904) );
  INVX2 U967 ( .A(\memory[7][3] ), .Y(n479) );
  MUX2X1 U968 ( .B(n479), .A(n517), .S(n127), .Y(n903) );
  INVX2 U969 ( .A(\memory[7][4] ), .Y(n480) );
  MUX2X1 U970 ( .B(n480), .A(n518), .S(n127), .Y(n902) );
  INVX2 U971 ( .A(\memory[7][5] ), .Y(n481) );
  MUX2X1 U972 ( .B(n481), .A(n519), .S(n127), .Y(n901) );
  INVX2 U973 ( .A(\memory[7][6] ), .Y(n482) );
  MUX2X1 U974 ( .B(n482), .A(n520), .S(n127), .Y(n900) );
  INVX2 U975 ( .A(\memory[7][7] ), .Y(n484) );
  MUX2X1 U976 ( .B(n484), .A(n521), .S(n127), .Y(n899) );
  INVX2 U977 ( .A(\memory[6][0] ), .Y(n485) );
  MUX2X1 U978 ( .B(n485), .A(n515), .S(n57), .Y(n896) );
  INVX2 U979 ( .A(\memory[6][1] ), .Y(n486) );
  MUX2X1 U980 ( .B(n486), .A(n516), .S(n492), .Y(n895) );
  INVX2 U981 ( .A(\memory[6][2] ), .Y(n487) );
  MUX2X1 U982 ( .B(n487), .A(n158), .S(n58), .Y(n894) );
  INVX2 U983 ( .A(\memory[6][3] ), .Y(n488) );
  MUX2X1 U984 ( .B(n488), .A(n517), .S(n57), .Y(n893) );
  INVX2 U985 ( .A(\memory[6][4] ), .Y(n489) );
  MUX2X1 U986 ( .B(n489), .A(n518), .S(n57), .Y(n892) );
  INVX2 U987 ( .A(\memory[6][5] ), .Y(n490) );
  MUX2X1 U988 ( .B(n490), .A(n519), .S(n58), .Y(n891) );
  INVX2 U989 ( .A(\memory[6][6] ), .Y(n491) );
  MUX2X1 U990 ( .B(n491), .A(n520), .S(n57), .Y(n890) );
  INVX2 U991 ( .A(\memory[6][7] ), .Y(n493) );
  MUX2X1 U992 ( .B(n493), .A(n521), .S(n58), .Y(n889) );
  INVX2 U993 ( .A(\memory[5][0] ), .Y(n494) );
  MUX2X1 U994 ( .B(n494), .A(n515), .S(n66), .Y(n886) );
  INVX2 U995 ( .A(\memory[5][1] ), .Y(n495) );
  MUX2X1 U996 ( .B(n495), .A(n516), .S(n66), .Y(n885) );
  INVX2 U997 ( .A(\memory[5][2] ), .Y(n496) );
  MUX2X1 U998 ( .B(n496), .A(n159), .S(n66), .Y(n884) );
  INVX2 U999 ( .A(\memory[5][3] ), .Y(n497) );
  MUX2X1 U1000 ( .B(n497), .A(n517), .S(n66), .Y(n883) );
  INVX2 U1001 ( .A(\memory[5][4] ), .Y(n498) );
  MUX2X1 U1002 ( .B(n498), .A(n518), .S(n66), .Y(n882) );
  INVX2 U1003 ( .A(\memory[5][5] ), .Y(n499) );
  MUX2X1 U1004 ( .B(n499), .A(n519), .S(n66), .Y(n881) );
  INVX2 U1005 ( .A(\memory[5][6] ), .Y(n500) );
  MUX2X1 U1006 ( .B(n500), .A(n520), .S(n66), .Y(n880) );
  INVX2 U1007 ( .A(\memory[5][7] ), .Y(n502) );
  MUX2X1 U1008 ( .B(n502), .A(n521), .S(n66), .Y(n879) );
  INVX2 U1009 ( .A(\memory[4][0] ), .Y(n503) );
  MUX2X1 U1010 ( .B(n503), .A(n515), .S(n39), .Y(n876) );
  INVX2 U1011 ( .A(\memory[4][1] ), .Y(n504) );
  MUX2X1 U1012 ( .B(n504), .A(n516), .S(n71), .Y(n875) );
  INVX2 U1013 ( .A(\memory[4][2] ), .Y(n505) );
  MUX2X1 U1014 ( .B(n505), .A(n158), .S(n39), .Y(n874) );
  INVX2 U1015 ( .A(\memory[4][3] ), .Y(n506) );
  MUX2X1 U1016 ( .B(n506), .A(n517), .S(n71), .Y(n873) );
  INVX2 U1017 ( .A(\memory[4][4] ), .Y(n507) );
  MUX2X1 U1018 ( .B(n507), .A(n518), .S(n510), .Y(n872) );
  INVX2 U1019 ( .A(\memory[4][5] ), .Y(n508) );
  MUX2X1 U1020 ( .B(n508), .A(n519), .S(n39), .Y(n871) );
  INVX2 U1021 ( .A(\memory[4][6] ), .Y(n509) );
  MUX2X1 U1022 ( .B(n509), .A(n520), .S(n71), .Y(n870) );
  INVX2 U1023 ( .A(\memory[4][7] ), .Y(n511) );
  MUX2X1 U1024 ( .B(n511), .A(n521), .S(n510), .Y(n869) );
  MUX2X1 U1025 ( .B(n738), .A(n515), .S(n47), .Y(n1406) );
  MUX2X1 U1026 ( .B(n739), .A(n516), .S(n3), .Y(n1407) );
  MUX2X1 U1027 ( .B(n740), .A(n159), .S(n3), .Y(n1408) );
  MUX2X1 U1028 ( .B(n741), .A(n517), .S(n3), .Y(n1409) );
  MUX2X1 U1029 ( .B(n742), .A(n162), .S(n47), .Y(n1410) );
  MUX2X1 U1030 ( .B(n743), .A(n519), .S(n3), .Y(n1411) );
  MUX2X1 U1031 ( .B(n744), .A(n166), .S(n47), .Y(n1412) );
  MUX2X1 U1032 ( .B(n745), .A(n168), .S(n3), .Y(n1413) );
  MUX2X1 U1033 ( .B(n730), .A(n515), .S(n513), .Y(n1398) );
  MUX2X1 U1034 ( .B(n731), .A(n516), .S(n513), .Y(n1399) );
  MUX2X1 U1035 ( .B(n732), .A(n158), .S(n40), .Y(n1400) );
  MUX2X1 U1036 ( .B(n733), .A(n517), .S(n40), .Y(n1401) );
  MUX2X1 U1037 ( .B(n734), .A(n162), .S(n513), .Y(n1402) );
  MUX2X1 U1038 ( .B(n735), .A(n519), .S(n40), .Y(n1403) );
  MUX2X1 U1039 ( .B(n736), .A(n166), .S(n513), .Y(n1404) );
  MUX2X1 U1040 ( .B(n737), .A(n168), .S(n40), .Y(n1405) );
  MUX2X1 U1041 ( .B(n722), .A(n515), .S(n48), .Y(n1390) );
  MUX2X1 U1042 ( .B(n723), .A(n516), .S(n4), .Y(n1391) );
  MUX2X1 U1043 ( .B(n724), .A(n159), .S(n4), .Y(n1392) );
  MUX2X1 U1044 ( .B(n725), .A(n517), .S(n4), .Y(n1393) );
  MUX2X1 U1045 ( .B(n726), .A(n162), .S(n48), .Y(n1394) );
  MUX2X1 U1046 ( .B(n727), .A(n519), .S(n4), .Y(n1395) );
  MUX2X1 U1047 ( .B(n728), .A(n166), .S(n48), .Y(n1396) );
  MUX2X1 U1048 ( .B(n729), .A(n168), .S(n4), .Y(n1397) );
  MUX2X1 U1049 ( .B(n714), .A(n515), .S(n79), .Y(n1382) );
  MUX2X1 U1050 ( .B(n715), .A(n516), .S(n80), .Y(n1383) );
  MUX2X1 U1051 ( .B(n716), .A(n158), .S(n70), .Y(n1384) );
  MUX2X1 U1052 ( .B(n717), .A(n517), .S(n80), .Y(n1385) );
  MUX2X1 U1053 ( .B(n718), .A(n162), .S(n79), .Y(n1386) );
  MUX2X1 U1054 ( .B(n719), .A(n519), .S(n70), .Y(n1387) );
  MUX2X1 U1055 ( .B(n720), .A(n166), .S(n70), .Y(n1388) );
  MUX2X1 U1056 ( .B(n721), .A(n168), .S(n80), .Y(n1389) );
  AND2X2 U1057 ( .A(state), .B(n522), .Y(N338) );
  XOR2X1 U1058 ( .A(n524), .B(n123), .Y(n523) );
  INVX2 U1059 ( .A(state), .Y(n598) );
  NOR2X1 U1060 ( .A(n523), .B(n598), .Y(N339) );
  NAND2X1 U1061 ( .A(n77), .B(n594), .Y(n526) );
  OAI21X1 U1062 ( .A(n77), .B(n594), .C(n524), .Y(n525) );
  AND2X2 U1063 ( .A(n526), .B(n525), .Y(n531) );
  XNOR2X1 U1064 ( .A(n531), .B(n527), .Y(n528) );
  AND2X2 U1065 ( .A(state), .B(n528), .Y(N340) );
  NOR2X1 U1066 ( .A(n149), .B(n663), .Y(n530) );
  NAND2X1 U1067 ( .A(n149), .B(n663), .Y(n529) );
  OAI21X1 U1068 ( .A(n531), .B(n530), .C(n529), .Y(n535) );
  XNOR2X1 U1069 ( .A(n535), .B(n532), .Y(n533) );
  NOR2X1 U1070 ( .A(n533), .B(n598), .Y(N341) );
  NAND2X1 U1071 ( .A(n153), .B(n568), .Y(n536) );
  NOR2X1 U1072 ( .A(n153), .B(n568), .Y(n534) );
  AOI21X1 U1073 ( .A(n536), .B(n535), .C(n534), .Y(n538) );
  XNOR2X1 U1074 ( .A(n538), .B(n28), .Y(n539) );
  AND2X2 U1075 ( .A(state), .B(n539), .Y(N342) );
  NOR2X1 U1076 ( .A(n85), .B(n540), .Y(n545) );
  AND2X2 U1077 ( .A(n6), .B(n541), .Y(n543) );
  NAND3X1 U1078 ( .A(n545), .B(n544), .C(n543), .Y(n546) );
  MUX2X1 U1079 ( .B(n546), .A(n746), .S(RST), .Y(n1414) );
  NAND2X1 U1080 ( .A(n89), .B(n38), .Y(n562) );
  INVX2 U1081 ( .A(n562), .Y(n576) );
  NAND2X1 U1082 ( .A(n576), .B(n27), .Y(n552) );
  NAND2X1 U1083 ( .A(n149), .B(n556), .Y(n548) );
  NAND2X1 U1084 ( .A(n548), .B(n565), .Y(n549) );
  NAND2X1 U1085 ( .A(n578), .B(n549), .Y(n551) );
  NAND2X1 U1086 ( .A(n149), .B(n558), .Y(n550) );
  NAND3X1 U1087 ( .A(n552), .B(n551), .C(n550), .Y(n854) );
  NAND2X1 U1088 ( .A(n576), .B(n554), .Y(n561) );
  NAND2X1 U1089 ( .A(n556), .B(n72), .Y(n557) );
  NAND2X1 U1090 ( .A(n578), .B(n557), .Y(n560) );
  NAND2X1 U1091 ( .A(n77), .B(n558), .Y(n559) );
  NAND3X1 U1092 ( .A(n561), .B(n560), .C(n559), .Y(n856) );
  MUX2X1 U1093 ( .B(n564), .A(n89), .S(n52), .Y(n858) );
  NAND2X1 U1094 ( .A(n566), .B(n565), .Y(n579) );
  NAND2X1 U1095 ( .A(n89), .B(n579), .Y(n567) );
  NAND2X1 U1096 ( .A(n94), .B(n567), .Y(n572) );
  XNOR2X1 U1097 ( .A(n569), .B(n568), .Y(n570) );
  NAND2X1 U1098 ( .A(n570), .B(n576), .Y(n571) );
  NAND3X1 U1099 ( .A(n572), .B(n577), .C(n571), .Y(n860) );
  XOR2X1 U1100 ( .A(n574), .B(n8), .Y(n575) );
  NAND2X1 U1101 ( .A(n576), .B(n575), .Y(n585) );
  NAND2X1 U1102 ( .A(n578), .B(n94), .Y(n580) );
  NAND3X1 U1103 ( .A(n89), .B(n580), .C(n579), .Y(n582) );
  MUX2X1 U1104 ( .B(n583), .A(n582), .S(n49), .Y(n584) );
  NAND2X1 U1105 ( .A(n585), .B(n584), .Y(n862) );
  NAND2X1 U1106 ( .A(n81), .B(n76), .Y(n595) );
  INVX2 U1107 ( .A(n595), .Y(n591) );
  NAND2X1 U1108 ( .A(n121), .B(n591), .Y(n589) );
  INVX2 U1109 ( .A(n589), .Y(n586) );
  NAND2X1 U1110 ( .A(n586), .B(n153), .Y(n587) );
  XNOR2X1 U1111 ( .A(n587), .B(n665), .Y(n588) );
  NOR2X1 U1112 ( .A(n598), .B(n588), .Y(N347) );
  XNOR2X1 U1113 ( .A(n589), .B(n664), .Y(n590) );
  NOR2X1 U1114 ( .A(n598), .B(n590), .Y(N346) );
  NAND2X1 U1115 ( .A(n120), .B(n591), .Y(n593) );
  OAI21X1 U1116 ( .A(n595), .B(n594), .C(n36), .Y(n592) );
  AOI21X1 U1117 ( .A(n593), .B(n592), .C(n598), .Y(N345) );
  XNOR2X1 U1118 ( .A(n595), .B(n594), .Y(n596) );
  NOR2X1 U1119 ( .A(n598), .B(n596), .Y(N344) );
  XNOR2X1 U1120 ( .A(n597), .B(n662), .Y(n599) );
  NOR2X1 U1121 ( .A(n599), .B(n598), .Y(N343) );
  INVX1 U1122 ( .A(FULL), .Y(n746) );
  INVX1 U1123 ( .A(EMPTY), .Y(n747) );
  NAND2X1 U1124 ( .A(n829), .B(n830), .Y(n828) );
  NOR2X1 U1125 ( .A(n831), .B(n832), .Y(n830) );
  NAND3X1 U1126 ( .A(n833), .B(n834), .C(n835), .Y(n832) );
  NOR2X1 U1127 ( .A(n836), .B(n837), .Y(n835) );
  OAI22X1 U1128 ( .A(n780), .B(n141), .C(n788), .D(n140), .Y(n837) );
  OAI22X1 U1129 ( .A(n796), .B(n128), .C(n804), .D(n130), .Y(n836) );
  AOI22X1 U1130 ( .A(n114), .B(\memory[23][7] ), .C(n110), .D(\memory[22][7] ), 
        .Y(n834) );
  AOI22X1 U1131 ( .A(n840), .B(\memory[21][7] ), .C(n841), .D(\memory[20][7] ), 
        .Y(n833) );
  NAND3X1 U1132 ( .A(n842), .B(n843), .C(n844), .Y(n831) );
  NOR2X1 U1133 ( .A(n845), .B(n846), .Y(n844) );
  OAI22X1 U1134 ( .A(n706), .B(n143), .C(n698), .D(n142), .Y(n846) );
  OAI22X1 U1135 ( .A(n690), .B(n131), .C(n682), .D(n132), .Y(n845) );
  AOI22X1 U1136 ( .A(n115), .B(\memory[31][7] ), .C(n112), .D(\memory[30][7] ), 
        .Y(n843) );
  AOI22X1 U1137 ( .A(n852), .B(\memory[29][7] ), .C(n865), .D(\memory[28][7] ), 
        .Y(n842) );
  NOR2X1 U1138 ( .A(n877), .B(n878), .Y(n829) );
  NAND3X1 U1139 ( .A(n887), .B(n888), .C(n897), .Y(n878) );
  NOR2X1 U1140 ( .A(n898), .B(n907), .Y(n897) );
  OAI22X1 U1141 ( .A(n745), .B(n133), .C(n737), .D(n134), .Y(n907) );
  OAI22X1 U1142 ( .A(n729), .B(n145), .C(n721), .D(n144), .Y(n898) );
  AOI22X1 U1143 ( .A(n908), .B(\memory[4][7] ), .C(n909), .D(\memory[5][7] ), 
        .Y(n888) );
  AOI22X1 U1144 ( .A(n116), .B(\memory[6][7] ), .C(n111), .D(\memory[7][7] ), 
        .Y(n887) );
  NAND3X1 U1145 ( .A(n910), .B(n911), .C(n912), .Y(n877) );
  NOR2X1 U1146 ( .A(n913), .B(n914), .Y(n912) );
  OAI22X1 U1147 ( .A(n748), .B(n147), .C(n756), .D(n146), .Y(n914) );
  OAI22X1 U1148 ( .A(n764), .B(n135), .C(n772), .D(n136), .Y(n913) );
  AOI22X1 U1149 ( .A(n113), .B(\memory[15][7] ), .C(n109), .D(\memory[14][7] ), 
        .Y(n911) );
  AOI22X1 U1150 ( .A(n915), .B(\memory[13][7] ), .C(n916), .D(\memory[12][7] ), 
        .Y(n910) );
  NAND2X1 U1151 ( .A(n918), .B(n919), .Y(n917) );
  NOR2X1 U1152 ( .A(n920), .B(n921), .Y(n919) );
  NAND3X1 U1153 ( .A(n922), .B(n923), .C(n924), .Y(n921) );
  NOR2X1 U1154 ( .A(n925), .B(n926), .Y(n924) );
  OAI22X1 U1155 ( .A(n781), .B(n141), .C(n789), .D(n140), .Y(n926) );
  OAI22X1 U1156 ( .A(n797), .B(n128), .C(n805), .D(n130), .Y(n925) );
  AOI22X1 U1157 ( .A(n114), .B(\memory[23][6] ), .C(n110), .D(\memory[22][6] ), 
        .Y(n923) );
  AOI22X1 U1158 ( .A(n840), .B(\memory[21][6] ), .C(n841), .D(\memory[20][6] ), 
        .Y(n922) );
  NAND3X1 U1159 ( .A(n927), .B(n928), .C(n929), .Y(n920) );
  NOR2X1 U1160 ( .A(n930), .B(n931), .Y(n929) );
  OAI22X1 U1161 ( .A(n707), .B(n143), .C(n699), .D(n142), .Y(n931) );
  OAI22X1 U1162 ( .A(n691), .B(n131), .C(n683), .D(n132), .Y(n930) );
  AOI22X1 U1163 ( .A(n115), .B(\memory[31][6] ), .C(n112), .D(\memory[30][6] ), 
        .Y(n928) );
  AOI22X1 U1164 ( .A(n852), .B(\memory[29][6] ), .C(n865), .D(\memory[28][6] ), 
        .Y(n927) );
  NOR2X1 U1165 ( .A(n932), .B(n933), .Y(n918) );
  NAND3X1 U1166 ( .A(n934), .B(n935), .C(n936), .Y(n933) );
  NOR2X1 U1167 ( .A(n937), .B(n938), .Y(n936) );
  OAI22X1 U1168 ( .A(n744), .B(n133), .C(n736), .D(n134), .Y(n938) );
  OAI22X1 U1169 ( .A(n728), .B(n145), .C(n720), .D(n144), .Y(n937) );
  AOI22X1 U1170 ( .A(n908), .B(\memory[4][6] ), .C(n909), .D(\memory[5][6] ), 
        .Y(n935) );
  AOI22X1 U1171 ( .A(n116), .B(\memory[6][6] ), .C(n111), .D(\memory[7][6] ), 
        .Y(n934) );
  NAND3X1 U1172 ( .A(n939), .B(n940), .C(n941), .Y(n932) );
  NOR2X1 U1173 ( .A(n942), .B(n943), .Y(n941) );
  OAI22X1 U1174 ( .A(n749), .B(n147), .C(n757), .D(n146), .Y(n943) );
  OAI22X1 U1175 ( .A(n765), .B(n135), .C(n773), .D(n136), .Y(n942) );
  AOI22X1 U1176 ( .A(n113), .B(\memory[15][6] ), .C(n109), .D(\memory[14][6] ), 
        .Y(n940) );
  AOI22X1 U1177 ( .A(n915), .B(\memory[13][6] ), .C(n916), .D(\memory[12][6] ), 
        .Y(n939) );
  NAND2X1 U1178 ( .A(n945), .B(n946), .Y(n944) );
  NOR2X1 U1179 ( .A(n947), .B(n948), .Y(n946) );
  NAND3X1 U1180 ( .A(n949), .B(n950), .C(n951), .Y(n948) );
  NOR2X1 U1181 ( .A(n952), .B(n953), .Y(n951) );
  OAI22X1 U1182 ( .A(n782), .B(n141), .C(n790), .D(n140), .Y(n953) );
  OAI22X1 U1183 ( .A(n798), .B(n128), .C(n806), .D(n130), .Y(n952) );
  AOI22X1 U1184 ( .A(n114), .B(\memory[23][5] ), .C(n110), .D(\memory[22][5] ), 
        .Y(n950) );
  AOI22X1 U1185 ( .A(n840), .B(\memory[21][5] ), .C(n841), .D(\memory[20][5] ), 
        .Y(n949) );
  NAND3X1 U1186 ( .A(n954), .B(n955), .C(n956), .Y(n947) );
  NOR2X1 U1187 ( .A(n957), .B(n958), .Y(n956) );
  OAI22X1 U1188 ( .A(n708), .B(n143), .C(n700), .D(n142), .Y(n958) );
  OAI22X1 U1189 ( .A(n692), .B(n131), .C(n684), .D(n132), .Y(n957) );
  AOI22X1 U1190 ( .A(n115), .B(\memory[31][5] ), .C(n112), .D(\memory[30][5] ), 
        .Y(n955) );
  AOI22X1 U1203 ( .A(n852), .B(\memory[29][5] ), .C(n865), .D(\memory[28][5] ), 
        .Y(n954) );
  NOR2X1 U1207 ( .A(n959), .B(n960), .Y(n945) );
  NAND3X1 U1208 ( .A(n961), .B(n962), .C(n963), .Y(n960) );
  NOR2X1 U1209 ( .A(n964), .B(n965), .Y(n963) );
  OAI22X1 U1210 ( .A(n743), .B(n133), .C(n735), .D(n134), .Y(n965) );
  OAI22X1 U1211 ( .A(n727), .B(n145), .C(n719), .D(n144), .Y(n964) );
  AOI22X1 U1212 ( .A(n908), .B(\memory[4][5] ), .C(n909), .D(\memory[5][5] ), 
        .Y(n962) );
  AOI22X1 U1213 ( .A(n116), .B(\memory[6][5] ), .C(n111), .D(\memory[7][5] ), 
        .Y(n961) );
  NAND3X1 U1214 ( .A(n966), .B(n967), .C(n968), .Y(n959) );
  NOR2X1 U1215 ( .A(n969), .B(n970), .Y(n968) );
  OAI22X1 U1216 ( .A(n750), .B(n147), .C(n758), .D(n146), .Y(n970) );
  OAI22X1 U1217 ( .A(n766), .B(n135), .C(n774), .D(n136), .Y(n969) );
  AOI22X1 U1218 ( .A(n113), .B(\memory[15][5] ), .C(n109), .D(\memory[14][5] ), 
        .Y(n967) );
  AOI22X1 U1219 ( .A(n915), .B(\memory[13][5] ), .C(n916), .D(\memory[12][5] ), 
        .Y(n966) );
  NAND2X1 U1220 ( .A(n972), .B(n973), .Y(n971) );
  NOR2X1 U1221 ( .A(n974), .B(n975), .Y(n973) );
  NAND3X1 U1222 ( .A(n976), .B(n977), .C(n978), .Y(n975) );
  NOR2X1 U1223 ( .A(n979), .B(n980), .Y(n978) );
  OAI22X1 U1224 ( .A(n783), .B(n141), .C(n791), .D(n140), .Y(n980) );
  OAI22X1 U1225 ( .A(n799), .B(n128), .C(n807), .D(n130), .Y(n979) );
  AOI22X1 U1226 ( .A(n114), .B(\memory[23][4] ), .C(n110), .D(\memory[22][4] ), 
        .Y(n977) );
  AOI22X1 U1227 ( .A(n840), .B(\memory[21][4] ), .C(n841), .D(\memory[20][4] ), 
        .Y(n976) );
  NAND3X1 U1228 ( .A(n981), .B(n982), .C(n983), .Y(n974) );
  NOR2X1 U1229 ( .A(n984), .B(n985), .Y(n983) );
  OAI22X1 U1230 ( .A(n709), .B(n143), .C(n701), .D(n142), .Y(n985) );
  OAI22X1 U1231 ( .A(n693), .B(n131), .C(n685), .D(n132), .Y(n984) );
  AOI22X1 U1232 ( .A(n115), .B(\memory[31][4] ), .C(n112), .D(\memory[30][4] ), 
        .Y(n982) );
  AOI22X1 U1233 ( .A(n852), .B(\memory[29][4] ), .C(n865), .D(\memory[28][4] ), 
        .Y(n981) );
  NOR2X1 U1234 ( .A(n986), .B(n987), .Y(n972) );
  NAND3X1 U1235 ( .A(n988), .B(n989), .C(n990), .Y(n987) );
  NOR2X1 U1236 ( .A(n991), .B(n992), .Y(n990) );
  OAI22X1 U1237 ( .A(n742), .B(n133), .C(n734), .D(n134), .Y(n992) );
  OAI22X1 U1238 ( .A(n726), .B(n145), .C(n718), .D(n144), .Y(n991) );
  AOI22X1 U1239 ( .A(n908), .B(\memory[4][4] ), .C(n909), .D(\memory[5][4] ), 
        .Y(n989) );
  AOI22X1 U1240 ( .A(n116), .B(\memory[6][4] ), .C(n111), .D(\memory[7][4] ), 
        .Y(n988) );
  NAND3X1 U1241 ( .A(n993), .B(n994), .C(n995), .Y(n986) );
  NOR2X1 U1242 ( .A(n996), .B(n997), .Y(n995) );
  OAI22X1 U1243 ( .A(n751), .B(n147), .C(n759), .D(n146), .Y(n997) );
  OAI22X1 U1244 ( .A(n767), .B(n135), .C(n775), .D(n136), .Y(n996) );
  AOI22X1 U1245 ( .A(n113), .B(\memory[15][4] ), .C(n109), .D(\memory[14][4] ), 
        .Y(n994) );
  AOI22X1 U1246 ( .A(n915), .B(\memory[13][4] ), .C(n916), .D(\memory[12][4] ), 
        .Y(n993) );
  NAND2X1 U1247 ( .A(n999), .B(n1000), .Y(n998) );
  NOR2X1 U1248 ( .A(n1001), .B(n1002), .Y(n1000) );
  NAND3X1 U1249 ( .A(n1003), .B(n1004), .C(n1005), .Y(n1002) );
  NOR2X1 U1250 ( .A(n1006), .B(n1007), .Y(n1005) );
  OAI22X1 U1251 ( .A(n784), .B(n141), .C(n792), .D(n140), .Y(n1007) );
  OAI22X1 U1252 ( .A(n800), .B(n128), .C(n808), .D(n130), .Y(n1006) );
  AOI22X1 U1253 ( .A(n114), .B(\memory[23][3] ), .C(n110), .D(\memory[22][3] ), 
        .Y(n1004) );
  AOI22X1 U1254 ( .A(n840), .B(\memory[21][3] ), .C(n841), .D(\memory[20][3] ), 
        .Y(n1003) );
  NAND3X1 U1255 ( .A(n1008), .B(n1009), .C(n1010), .Y(n1001) );
  NOR2X1 U1256 ( .A(n1011), .B(n1012), .Y(n1010) );
  OAI22X1 U1257 ( .A(n710), .B(n143), .C(n702), .D(n142), .Y(n1012) );
  OAI22X1 U1258 ( .A(n694), .B(n131), .C(n686), .D(n132), .Y(n1011) );
  AOI22X1 U1259 ( .A(n115), .B(\memory[31][3] ), .C(n112), .D(\memory[30][3] ), 
        .Y(n1009) );
  AOI22X1 U1260 ( .A(n852), .B(\memory[29][3] ), .C(n865), .D(\memory[28][3] ), 
        .Y(n1008) );
  NOR2X1 U1261 ( .A(n1013), .B(n1014), .Y(n999) );
  NAND3X1 U1262 ( .A(n1015), .B(n1016), .C(n1017), .Y(n1014) );
  NOR2X1 U1263 ( .A(n1018), .B(n1019), .Y(n1017) );
  OAI22X1 U1264 ( .A(n741), .B(n133), .C(n733), .D(n134), .Y(n1019) );
  OAI22X1 U1265 ( .A(n725), .B(n145), .C(n717), .D(n144), .Y(n1018) );
  AOI22X1 U1266 ( .A(n908), .B(\memory[4][3] ), .C(n909), .D(\memory[5][3] ), 
        .Y(n1016) );
  AOI22X1 U1267 ( .A(n116), .B(\memory[6][3] ), .C(n111), .D(\memory[7][3] ), 
        .Y(n1015) );
  NAND3X1 U1268 ( .A(n1020), .B(n1021), .C(n1022), .Y(n1013) );
  NOR2X1 U1269 ( .A(n1023), .B(n1024), .Y(n1022) );
  OAI22X1 U1270 ( .A(n752), .B(n147), .C(n760), .D(n146), .Y(n1024) );
  OAI22X1 U1271 ( .A(n768), .B(n135), .C(n776), .D(n136), .Y(n1023) );
  AOI22X1 U1272 ( .A(n113), .B(\memory[15][3] ), .C(n109), .D(\memory[14][3] ), 
        .Y(n1021) );
  AOI22X1 U1273 ( .A(n915), .B(\memory[13][3] ), .C(n916), .D(\memory[12][3] ), 
        .Y(n1020) );
  NAND2X1 U1274 ( .A(n1026), .B(n1027), .Y(n1025) );
  NOR2X1 U1275 ( .A(n1028), .B(n1029), .Y(n1027) );
  NAND3X1 U1276 ( .A(n1040), .B(n1041), .C(n1042), .Y(n1029) );
  NOR2X1 U1277 ( .A(n1043), .B(n1044), .Y(n1042) );
  OAI22X1 U1278 ( .A(n785), .B(n141), .C(n793), .D(n140), .Y(n1044) );
  OAI22X1 U1279 ( .A(n801), .B(n128), .C(n809), .D(n130), .Y(n1043) );
  AOI22X1 U1280 ( .A(n114), .B(\memory[23][2] ), .C(n110), .D(\memory[22][2] ), 
        .Y(n1041) );
  AOI22X1 U1281 ( .A(n840), .B(\memory[21][2] ), .C(n841), .D(\memory[20][2] ), 
        .Y(n1040) );
  NAND3X1 U1282 ( .A(n1045), .B(n1046), .C(n1047), .Y(n1028) );
  NOR2X1 U1283 ( .A(n1048), .B(n1049), .Y(n1047) );
  OAI22X1 U1284 ( .A(n711), .B(n143), .C(n703), .D(n142), .Y(n1049) );
  OAI22X1 U1285 ( .A(n695), .B(n131), .C(n687), .D(n132), .Y(n1048) );
  AOI22X1 U1286 ( .A(n115), .B(\memory[31][2] ), .C(n112), .D(\memory[30][2] ), 
        .Y(n1046) );
  AOI22X1 U1287 ( .A(n852), .B(\memory[29][2] ), .C(n865), .D(\memory[28][2] ), 
        .Y(n1045) );
  NOR2X1 U1288 ( .A(n1050), .B(n1051), .Y(n1026) );
  NAND3X1 U1289 ( .A(n1052), .B(n1053), .C(n1054), .Y(n1051) );
  NOR2X1 U1290 ( .A(n1055), .B(n1058), .Y(n1054) );
  OAI22X1 U1291 ( .A(n740), .B(n133), .C(n732), .D(n134), .Y(n1058) );
  OAI22X1 U1292 ( .A(n724), .B(n145), .C(n716), .D(n144), .Y(n1055) );
  AOI22X1 U1293 ( .A(n908), .B(\memory[4][2] ), .C(n909), .D(\memory[5][2] ), 
        .Y(n1053) );
  AOI22X1 U1294 ( .A(n116), .B(\memory[6][2] ), .C(n111), .D(\memory[7][2] ), 
        .Y(n1052) );
  NAND3X1 U1295 ( .A(n1059), .B(n1060), .C(n1061), .Y(n1050) );
  NOR2X1 U1296 ( .A(n1062), .B(n1063), .Y(n1061) );
  OAI22X1 U1297 ( .A(n753), .B(n147), .C(n761), .D(n146), .Y(n1063) );
  OAI22X1 U1298 ( .A(n769), .B(n135), .C(n777), .D(n136), .Y(n1062) );
  AOI22X1 U1299 ( .A(n113), .B(\memory[15][2] ), .C(n109), .D(\memory[14][2] ), 
        .Y(n1060) );
  AOI22X1 U1300 ( .A(n915), .B(\memory[13][2] ), .C(n916), .D(\memory[12][2] ), 
        .Y(n1059) );
  NAND2X1 U1301 ( .A(n1065), .B(n1066), .Y(n1064) );
  NOR2X1 U1302 ( .A(n1067), .B(n1068), .Y(n1066) );
  NAND3X1 U1303 ( .A(n1069), .B(n1070), .C(n1071), .Y(n1068) );
  NOR2X1 U1304 ( .A(n1168), .B(n1169), .Y(n1071) );
  OAI22X1 U1305 ( .A(n786), .B(n141), .C(n794), .D(n140), .Y(n1169) );
  OAI22X1 U1306 ( .A(n802), .B(n128), .C(n810), .D(n130), .Y(n1168) );
  AOI22X1 U1307 ( .A(n114), .B(\memory[23][1] ), .C(n110), .D(\memory[22][1] ), 
        .Y(n1070) );
  AOI22X1 U1308 ( .A(n840), .B(\memory[21][1] ), .C(n841), .D(\memory[20][1] ), 
        .Y(n1069) );
  NAND3X1 U1309 ( .A(n1170), .B(n1171), .C(n1172), .Y(n1067) );
  NOR2X1 U1310 ( .A(n1173), .B(n1174), .Y(n1172) );
  OAI22X1 U1311 ( .A(n712), .B(n143), .C(n704), .D(n142), .Y(n1174) );
  OAI22X1 U1312 ( .A(n696), .B(n131), .C(n688), .D(n132), .Y(n1173) );
  AOI22X1 U1313 ( .A(n115), .B(\memory[31][1] ), .C(n112), .D(\memory[30][1] ), 
        .Y(n1171) );
  AOI22X1 U1314 ( .A(n852), .B(\memory[29][1] ), .C(n865), .D(\memory[28][1] ), 
        .Y(n1170) );
  NOR2X1 U1315 ( .A(n1175), .B(n1176), .Y(n1065) );
  NAND3X1 U1316 ( .A(n1177), .B(n1178), .C(n1179), .Y(n1176) );
  NOR2X1 U1317 ( .A(n1180), .B(n1181), .Y(n1179) );
  OAI22X1 U1318 ( .A(n739), .B(n133), .C(n731), .D(n134), .Y(n1181) );
  OAI22X1 U1319 ( .A(n723), .B(n145), .C(n715), .D(n144), .Y(n1180) );
  AOI22X1 U1320 ( .A(n908), .B(\memory[4][1] ), .C(n909), .D(\memory[5][1] ), 
        .Y(n1178) );
  AOI22X1 U1321 ( .A(n116), .B(\memory[6][1] ), .C(n111), .D(\memory[7][1] ), 
        .Y(n1177) );
  NAND3X1 U1322 ( .A(n1182), .B(n1183), .C(n1184), .Y(n1175) );
  NOR2X1 U1323 ( .A(n1185), .B(n1186), .Y(n1184) );
  OAI22X1 U1324 ( .A(n754), .B(n147), .C(n762), .D(n146), .Y(n1186) );
  OAI22X1 U1325 ( .A(n770), .B(n135), .C(n778), .D(n136), .Y(n1185) );
  AOI22X1 U1326 ( .A(n113), .B(\memory[15][1] ), .C(n109), .D(\memory[14][1] ), 
        .Y(n1183) );
  AOI22X1 U1327 ( .A(n915), .B(\memory[13][1] ), .C(n916), .D(\memory[12][1] ), 
        .Y(n1182) );
  NAND2X1 U1328 ( .A(n1188), .B(n1189), .Y(n1187) );
  NOR2X1 U1329 ( .A(n1190), .B(n1191), .Y(n1189) );
  NAND3X1 U1330 ( .A(n1192), .B(n1193), .C(n1194), .Y(n1191) );
  NOR2X1 U1331 ( .A(n1195), .B(n1196), .Y(n1194) );
  OAI22X1 U1332 ( .A(n787), .B(n141), .C(n795), .D(n140), .Y(n1196) );
  OAI22X1 U1333 ( .A(n803), .B(n128), .C(n811), .D(n130), .Y(n1195) );
  AOI22X1 U1334 ( .A(n114), .B(\memory[23][0] ), .C(n110), .D(\memory[22][0] ), 
        .Y(n1193) );
  AOI22X1 U1335 ( .A(n840), .B(\memory[21][0] ), .C(n841), .D(\memory[20][0] ), 
        .Y(n1192) );
  NAND3X1 U1336 ( .A(n1197), .B(n1198), .C(n1199), .Y(n1190) );
  NOR2X1 U1337 ( .A(n1200), .B(n1201), .Y(n1199) );
  OAI22X1 U1338 ( .A(n713), .B(n143), .C(n705), .D(n142), .Y(n1201) );
  OAI22X1 U1339 ( .A(n697), .B(n131), .C(n689), .D(n132), .Y(n1200) );
  AOI22X1 U1340 ( .A(n115), .B(\memory[31][0] ), .C(n112), .D(\memory[30][0] ), 
        .Y(n1198) );
  AOI22X1 U1341 ( .A(n852), .B(\memory[29][0] ), .C(n865), .D(\memory[28][0] ), 
        .Y(n1197) );
  NOR2X1 U1342 ( .A(n1202), .B(n1203), .Y(n1188) );
  NAND3X1 U1343 ( .A(n1204), .B(n1205), .C(n1206), .Y(n1203) );
  NOR2X1 U1344 ( .A(n1207), .B(n1208), .Y(n1206) );
  OAI22X1 U1345 ( .A(n738), .B(n133), .C(n730), .D(n134), .Y(n1208) );
  OAI22X1 U1346 ( .A(n722), .B(n145), .C(n714), .D(n144), .Y(n1207) );
  AOI22X1 U1347 ( .A(n908), .B(\memory[4][0] ), .C(n909), .D(\memory[5][0] ), 
        .Y(n1205) );
  AOI22X1 U1348 ( .A(n116), .B(\memory[6][0] ), .C(n111), .D(\memory[7][0] ), 
        .Y(n1204) );
  NAND3X1 U1349 ( .A(n1209), .B(n1210), .C(n1211), .Y(n1202) );
  NOR2X1 U1350 ( .A(n1212), .B(n1213), .Y(n1211) );
  OAI22X1 U1351 ( .A(n755), .B(n147), .C(n763), .D(n146), .Y(n1213) );
  OAI22X1 U1352 ( .A(n771), .B(n135), .C(n779), .D(n136), .Y(n1212) );
  AOI22X1 U1353 ( .A(n113), .B(\memory[15][0] ), .C(n109), .D(\memory[14][0] ), 
        .Y(n1210) );
  AOI22X1 U1354 ( .A(n915), .B(\memory[13][0] ), .C(n916), .D(\memory[12][0] ), 
        .Y(n1209) );
  NAND2X1 U1355 ( .A(n1215), .B(n1216), .Y(n1214) );
  NOR2X1 U1356 ( .A(n1217), .B(n1218), .Y(n1216) );
  NAND3X1 U1357 ( .A(n1219), .B(n1220), .C(n1221), .Y(n1218) );
  NOR2X1 U1358 ( .A(n1222), .B(n1223), .Y(n1221) );
  OAI22X1 U1359 ( .A(n820), .B(n141), .C(n822), .D(n140), .Y(n1223) );
  OAI22X1 U1360 ( .A(n824), .B(n128), .C(n826), .D(n130), .Y(n1222) );
  AOI22X1 U1361 ( .A(n114), .B(\opcode[23][1] ), .C(n110), .D(\opcode[22][1] ), 
        .Y(n1220) );
  AOI22X1 U1362 ( .A(n840), .B(\opcode[21][1] ), .C(n841), .D(\opcode[20][1] ), 
        .Y(n1219) );
  NAND3X1 U1363 ( .A(n1224), .B(n1225), .C(n1226), .Y(n1217) );
  NOR2X1 U1364 ( .A(n1227), .B(n1228), .Y(n1226) );
  OAI22X1 U1365 ( .A(n672), .B(n143), .C(n670), .D(n142), .Y(n1228) );
  OAI22X1 U1366 ( .A(n668), .B(n131), .C(n666), .D(n132), .Y(n1227) );
  AOI22X1 U1367 ( .A(n115), .B(\opcode[31][1] ), .C(n112), .D(\opcode[30][1] ), 
        .Y(n1225) );
  AOI22X1 U1368 ( .A(n852), .B(\opcode[29][1] ), .C(n865), .D(\opcode[28][1] ), 
        .Y(n1224) );
  NOR2X1 U1369 ( .A(n1229), .B(n1230), .Y(n1215) );
  NAND3X1 U1370 ( .A(n1231), .B(n1232), .C(n1233), .Y(n1230) );
  NOR2X1 U1371 ( .A(n1234), .B(n1235), .Y(n1233) );
  OAI22X1 U1372 ( .A(n681), .B(n133), .C(n679), .D(n134), .Y(n1235) );
  OAI22X1 U1373 ( .A(n677), .B(n145), .C(n675), .D(n144), .Y(n1234) );
  AOI22X1 U1374 ( .A(n908), .B(\opcode[4][1] ), .C(n909), .D(\opcode[5][1] ), 
        .Y(n1232) );
  AOI22X1 U1375 ( .A(n116), .B(\opcode[6][1] ), .C(n111), .D(\opcode[7][1] ), 
        .Y(n1231) );
  NAND3X1 U1376 ( .A(n1236), .B(n1237), .C(n1238), .Y(n1229) );
  NOR2X1 U1377 ( .A(n1239), .B(n1240), .Y(n1238) );
  OAI22X1 U1378 ( .A(n812), .B(n147), .C(n814), .D(n146), .Y(n1240) );
  OAI22X1 U1379 ( .A(n816), .B(n135), .C(n818), .D(n136), .Y(n1239) );
  AOI22X1 U1380 ( .A(n113), .B(\opcode[15][1] ), .C(n109), .D(\opcode[14][1] ), 
        .Y(n1237) );
  AOI22X1 U1381 ( .A(n915), .B(\opcode[13][1] ), .C(n916), .D(\opcode[12][1] ), 
        .Y(n1236) );
  NAND2X1 U1382 ( .A(n1242), .B(n1243), .Y(n1241) );
  NOR2X1 U1383 ( .A(n1244), .B(n1245), .Y(n1243) );
  NAND3X1 U1384 ( .A(n1246), .B(n1247), .C(n1248), .Y(n1245) );
  NOR2X1 U1385 ( .A(n1249), .B(n1250), .Y(n1248) );
  OAI22X1 U1386 ( .A(n821), .B(n141), .C(n823), .D(n140), .Y(n1250) );
  NAND2X1 U1387 ( .A(n1251), .B(n1252), .Y(n838) );
  OAI22X1 U1388 ( .A(n825), .B(n128), .C(n827), .D(n130), .Y(n1249) );
  AOI22X1 U1389 ( .A(n114), .B(\opcode[23][0] ), .C(n110), .D(\opcode[22][0] ), 
        .Y(n1247) );
  AOI22X1 U1390 ( .A(n840), .B(\opcode[21][0] ), .C(n841), .D(\opcode[20][0] ), 
        .Y(n1246) );
  INVX1 U1391 ( .A(n1255), .Y(n1253) );
  NAND3X1 U1392 ( .A(n662), .B(n664), .C(n84), .Y(n1255) );
  INVX1 U1393 ( .A(n1256), .Y(n1251) );
  NAND3X1 U1394 ( .A(n76), .B(n664), .C(n84), .Y(n1256) );
  NAND3X1 U1395 ( .A(n1257), .B(n1258), .C(n1259), .Y(n1244) );
  NOR2X1 U1396 ( .A(n1260), .B(n1261), .Y(n1259) );
  OAI22X1 U1397 ( .A(n673), .B(n143), .C(n671), .D(n142), .Y(n1261) );
  OAI22X1 U1398 ( .A(n669), .B(n131), .C(n667), .D(n132), .Y(n1260) );
  AOI22X1 U1399 ( .A(n115), .B(\opcode[31][0] ), .C(n112), .D(\opcode[30][0] ), 
        .Y(n1258) );
  AOI22X1 U1400 ( .A(n852), .B(\opcode[29][0] ), .C(n865), .D(\opcode[28][0] ), 
        .Y(n1257) );
  INVX1 U1401 ( .A(n1264), .Y(n1263) );
  NAND3X1 U1402 ( .A(n153), .B(n662), .C(n84), .Y(n1264) );
  INVX1 U1403 ( .A(n1265), .Y(n1262) );
  NAND3X1 U1404 ( .A(n153), .B(n76), .C(n84), .Y(n1265) );
  NOR2X1 U1405 ( .A(n1266), .B(n1267), .Y(n1242) );
  NAND3X1 U1406 ( .A(n1268), .B(n1269), .C(n1270), .Y(n1267) );
  NOR2X1 U1407 ( .A(n1271), .B(n1272), .Y(n1270) );
  OAI22X1 U1408 ( .A(n680), .B(n133), .C(n678), .D(n134), .Y(n1272) );
  OAI22X1 U1409 ( .A(n676), .B(n145), .C(n674), .D(n144), .Y(n1271) );
  AOI22X1 U1410 ( .A(n908), .B(\opcode[4][0] ), .C(n909), .D(\opcode[5][0] ), 
        .Y(n1269) );
  AOI22X1 U1411 ( .A(n116), .B(\opcode[6][0] ), .C(n111), .D(\opcode[7][0] ), 
        .Y(n1268) );
  INVX1 U1412 ( .A(n1275), .Y(n1274) );
  NAND3X1 U1413 ( .A(n664), .B(n665), .C(n76), .Y(n1275) );
  INVX1 U1414 ( .A(n1276), .Y(n1273) );
  NAND3X1 U1415 ( .A(n664), .B(n665), .C(n662), .Y(n1276) );
  NAND3X1 U1416 ( .A(n1277), .B(n1278), .C(n1279), .Y(n1266) );
  NOR2X1 U1417 ( .A(n1280), .B(n1281), .Y(n1279) );
  OAI22X1 U1418 ( .A(n813), .B(n147), .C(n815), .D(n146), .Y(n1281) );
  NOR2X1 U1419 ( .A(n51), .B(readptr[2]), .Y(n1252) );
  OAI22X1 U1420 ( .A(n817), .B(n135), .C(n819), .D(n136), .Y(n1280) );
  AOI22X1 U1421 ( .A(n113), .B(\opcode[15][0] ), .C(n109), .D(\opcode[14][0] ), 
        .Y(n1278) );
  AOI22X1 U1422 ( .A(n915), .B(\opcode[13][0] ), .C(n916), .D(\opcode[12][0] ), 
        .Y(n1277) );
  INVX1 U1423 ( .A(n1284), .Y(n1283) );
  NAND3X1 U1424 ( .A(n662), .B(n665), .C(n153), .Y(n1284) );
  NOR2X1 U1425 ( .A(n663), .B(n51), .Y(n1254) );
  INVX1 U1426 ( .A(n1285), .Y(n1282) );
  NAND3X1 U1427 ( .A(n76), .B(n665), .C(n153), .Y(n1285) );
endmodule


module memoryblock_1 ( CLK, NEXT_BYTE, RCV_DATA, RCV_OPCODE, RST, W_ENABLE, 
        EOP, EMPTY, FULL, B_READY, PRGA_IN, PRGA_OPCODE );
  input [7:0] RCV_DATA;
  input [1:0] RCV_OPCODE;
  output [7:0] PRGA_IN;
  output [1:0] PRGA_OPCODE;
  input CLK, NEXT_BYTE, RST, W_ENABLE, EOP;
  output EMPTY, FULL, B_READY;
  wire   R_ENABLE;
  wire   [4:0] BYTE_COUNT;
  wire   [7:0] DATA;
  wire   [1:0] OUT_OPCODE;

  RBUFFER_1 U_0 ( .CLK(CLK), .RST(RST), .NEXT_BYTE(NEXT_BYTE), .DATA(DATA), 
        .OPCODE(OUT_OPCODE), .BYTE_COUNT(BYTE_COUNT), .EOP(EOP), .B_READY(
        B_READY), .R_ENABLE(R_ENABLE), .PRGA_IN(PRGA_IN), .PRGA_OPCODE(
        PRGA_OPCODE) );
  RFIFO_1 U_1 ( .CLK(CLK), .RST(RST), .W_ENABLE(W_ENABLE), .R_ENABLE(R_ENABLE), 
        .RCV_DATA(RCV_DATA), .RCV_OPCODE(RCV_OPCODE), .DATA(DATA), 
        .OUT_OPCODE(OUT_OPCODE), .BYTE_COUNT(BYTE_COUNT), .EMPTY(EMPTY), 
        .FULL(FULL) );
endmodule


module rx_CRC_CALC_1 ( CLK, RST, W_ENABLE, OPCODE, RCV_DATA, RX_CRC );
  input [1:0] OPCODE;
  input [7:0] RCV_DATA;
  output [15:0] RX_CRC;
  input CLK, RST, W_ENABLE;
  wire   n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n101, n103, n105, n107, n109, n111, n113, n115, n117,
         n119, n121, n123, n125, n127, n129, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n1,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n100, n102, n104, n106,
         n108, n110, n112, n114, n116, n118, n120, n122, n124, n126, n128,
         n130, n131, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172;
  wire   [15:0] current_crc;
  wire   [15:0] cache_1;

  DFFPOSX1 \cache_1_reg[0]  ( .D(n129), .CLK(CLK), .Q(cache_1[0]) );
  DFFPOSX1 \cache_1_reg[8]  ( .D(n127), .CLK(CLK), .Q(cache_1[8]) );
  DFFPOSX1 \cache_1_reg[15]  ( .D(n125), .CLK(CLK), .Q(cache_1[15]) );
  DFFPOSX1 \cache_1_reg[1]  ( .D(n123), .CLK(CLK), .Q(cache_1[1]) );
  DFFPOSX1 \cache_1_reg[9]  ( .D(n121), .CLK(CLK), .Q(cache_1[9]) );
  DFFPOSX1 \cache_1_reg[2]  ( .D(n119), .CLK(CLK), .Q(cache_1[2]) );
  DFFPOSX1 \cache_1_reg[10]  ( .D(n117), .CLK(CLK), .Q(cache_1[10]) );
  DFFPOSX1 \cache_1_reg[3]  ( .D(n115), .CLK(CLK), .Q(cache_1[3]) );
  DFFPOSX1 \cache_1_reg[11]  ( .D(n113), .CLK(CLK), .Q(cache_1[11]) );
  DFFPOSX1 \cache_1_reg[4]  ( .D(n111), .CLK(CLK), .Q(cache_1[4]) );
  DFFPOSX1 \cache_1_reg[12]  ( .D(n109), .CLK(CLK), .Q(cache_1[12]) );
  DFFPOSX1 \cache_1_reg[5]  ( .D(n107), .CLK(CLK), .Q(cache_1[5]) );
  DFFPOSX1 \cache_1_reg[13]  ( .D(n105), .CLK(CLK), .Q(cache_1[13]) );
  DFFPOSX1 \cache_1_reg[6]  ( .D(n103), .CLK(CLK), .Q(cache_1[6]) );
  DFFPOSX1 \cache_1_reg[14]  ( .D(n101), .CLK(CLK), .Q(cache_1[14]) );
  DFFPOSX1 \cache_1_reg[7]  ( .D(n99), .CLK(CLK), .Q(cache_1[7]) );
  DFFPOSX1 \cache_2_reg[15]  ( .D(n98), .CLK(CLK), .Q(RX_CRC[15]) );
  DFFPOSX1 \cache_2_reg[14]  ( .D(n97), .CLK(CLK), .Q(RX_CRC[14]) );
  DFFPOSX1 \cache_2_reg[13]  ( .D(n96), .CLK(CLK), .Q(RX_CRC[13]) );
  DFFPOSX1 \cache_2_reg[12]  ( .D(n95), .CLK(CLK), .Q(RX_CRC[12]) );
  DFFPOSX1 \cache_2_reg[11]  ( .D(n94), .CLK(CLK), .Q(RX_CRC[11]) );
  DFFPOSX1 \cache_2_reg[10]  ( .D(n93), .CLK(CLK), .Q(RX_CRC[10]) );
  DFFPOSX1 \cache_2_reg[9]  ( .D(n92), .CLK(CLK), .Q(RX_CRC[9]) );
  DFFPOSX1 \cache_2_reg[8]  ( .D(n91), .CLK(CLK), .Q(RX_CRC[8]) );
  DFFPOSX1 \cache_2_reg[7]  ( .D(n90), .CLK(CLK), .Q(RX_CRC[7]) );
  DFFPOSX1 \cache_2_reg[6]  ( .D(n89), .CLK(CLK), .Q(RX_CRC[6]) );
  DFFPOSX1 \cache_2_reg[5]  ( .D(n88), .CLK(CLK), .Q(RX_CRC[5]) );
  DFFPOSX1 \cache_2_reg[4]  ( .D(n87), .CLK(CLK), .Q(RX_CRC[4]) );
  DFFPOSX1 \cache_2_reg[3]  ( .D(n86), .CLK(CLK), .Q(RX_CRC[3]) );
  DFFPOSX1 \cache_2_reg[2]  ( .D(n85), .CLK(CLK), .Q(RX_CRC[2]) );
  DFFPOSX1 \cache_2_reg[1]  ( .D(n84), .CLK(CLK), .Q(RX_CRC[1]) );
  DFFPOSX1 \cache_2_reg[0]  ( .D(n83), .CLK(CLK), .Q(RX_CRC[0]) );
  DFFSR \current_crc_reg[15]  ( .D(n132), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[15]) );
  DFFSR \current_crc_reg[14]  ( .D(n133), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[14]) );
  DFFSR \current_crc_reg[13]  ( .D(n134), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[13]) );
  DFFSR \current_crc_reg[12]  ( .D(n135), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[12]) );
  DFFSR \current_crc_reg[11]  ( .D(n136), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[11]) );
  DFFSR \current_crc_reg[10]  ( .D(n137), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[10]) );
  DFFSR \current_crc_reg[9]  ( .D(n138), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[9]) );
  DFFSR \current_crc_reg[8]  ( .D(n139), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[8]) );
  DFFSR \current_crc_reg[7]  ( .D(n140), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[7]) );
  DFFSR \current_crc_reg[6]  ( .D(n141), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[6]) );
  DFFSR \current_crc_reg[5]  ( .D(n142), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[5]) );
  DFFSR \current_crc_reg[4]  ( .D(n143), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[4]) );
  DFFSR \current_crc_reg[3]  ( .D(n144), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[3]) );
  DFFSR \current_crc_reg[2]  ( .D(n145), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[2]) );
  DFFSR \current_crc_reg[1]  ( .D(n146), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[1]) );
  DFFSR \current_crc_reg[0]  ( .D(n147), .CLK(CLK), .R(n35), .S(1'b1), .Q(
        current_crc[0]) );
  INVX2 U3 ( .A(n28), .Y(n20) );
  XOR2X1 U4 ( .A(n27), .B(n25), .Y(n1) );
  INVX2 U21 ( .A(n53), .Y(n19) );
  INVX2 U22 ( .A(OPCODE[1]), .Y(n34) );
  AND2X2 U23 ( .A(n19), .B(n35), .Y(n18) );
  INVX4 U24 ( .A(n21), .Y(n33) );
  AND2X2 U25 ( .A(n19), .B(n35), .Y(n21) );
  INVX2 U26 ( .A(n22), .Y(n30) );
  INVX2 U27 ( .A(n22), .Y(n29) );
  AND2X2 U28 ( .A(n54), .B(n28), .Y(n22) );
  INVX2 U29 ( .A(RST), .Y(n35) );
  XNOR2X1 U30 ( .A(n63), .B(n27), .Y(n64) );
  XNOR2X1 U31 ( .A(RCV_DATA[6]), .B(current_crc[14]), .Y(n161) );
  XNOR2X1 U32 ( .A(RCV_DATA[7]), .B(current_crc[15]), .Y(n148) );
  XOR2X1 U33 ( .A(RCV_DATA[0]), .B(current_crc[8]), .Y(n23) );
  XNOR2X1 U34 ( .A(RCV_DATA[5]), .B(current_crc[13]), .Y(n63) );
  XOR2X1 U35 ( .A(RCV_DATA[1]), .B(current_crc[9]), .Y(n24) );
  XOR2X1 U36 ( .A(RCV_DATA[3]), .B(current_crc[11]), .Y(n25) );
  XOR2X1 U37 ( .A(RCV_DATA[2]), .B(current_crc[10]), .Y(n26) );
  XOR2X1 U38 ( .A(RCV_DATA[4]), .B(current_crc[12]), .Y(n27) );
  NAND3X1 U39 ( .A(OPCODE[0]), .B(W_ENABLE), .C(n34), .Y(n28) );
  INVX8 U40 ( .A(n33), .Y(n31) );
  INVX8 U41 ( .A(n33), .Y(n32) );
  INVX2 U42 ( .A(RX_CRC[0]), .Y(n36) );
  INVX2 U43 ( .A(cache_1[0]), .Y(n165) );
  NAND3X1 U44 ( .A(OPCODE[0]), .B(W_ENABLE), .C(n34), .Y(n53) );
  MUX2X1 U45 ( .B(n36), .A(n165), .S(n31), .Y(n83) );
  INVX2 U46 ( .A(RX_CRC[1]), .Y(n37) );
  INVX2 U47 ( .A(cache_1[1]), .Y(n130) );
  MUX2X1 U48 ( .B(n37), .A(n130), .S(n32), .Y(n84) );
  INVX2 U49 ( .A(RX_CRC[2]), .Y(n38) );
  INVX2 U50 ( .A(cache_1[2]), .Y(n114) );
  MUX2X1 U51 ( .B(n38), .A(n114), .S(n31), .Y(n85) );
  INVX2 U52 ( .A(RX_CRC[3]), .Y(n39) );
  INVX2 U53 ( .A(cache_1[3]), .Y(n100) );
  MUX2X1 U54 ( .B(n39), .A(n100), .S(n32), .Y(n86) );
  INVX2 U55 ( .A(RX_CRC[4]), .Y(n40) );
  INVX2 U56 ( .A(cache_1[4]), .Y(n76) );
  MUX2X1 U57 ( .B(n40), .A(n76), .S(n31), .Y(n87) );
  INVX2 U58 ( .A(RX_CRC[5]), .Y(n41) );
  INVX2 U59 ( .A(cache_1[5]), .Y(n70) );
  MUX2X1 U60 ( .B(n41), .A(n70), .S(n31), .Y(n88) );
  INVX2 U61 ( .A(RX_CRC[6]), .Y(n42) );
  INVX2 U62 ( .A(cache_1[6]), .Y(n62) );
  MUX2X1 U63 ( .B(n42), .A(n62), .S(n31), .Y(n89) );
  INVX2 U64 ( .A(RX_CRC[7]), .Y(n43) );
  INVX2 U65 ( .A(cache_1[7]), .Y(n52) );
  MUX2X1 U66 ( .B(n43), .A(n52), .S(n32), .Y(n90) );
  INVX2 U67 ( .A(RX_CRC[8]), .Y(n44) );
  INVX2 U68 ( .A(cache_1[8]), .Y(n160) );
  MUX2X1 U69 ( .B(n44), .A(n160), .S(n31), .Y(n91) );
  INVX2 U70 ( .A(RX_CRC[9]), .Y(n45) );
  INVX2 U71 ( .A(cache_1[9]), .Y(n122) );
  MUX2X1 U72 ( .B(n45), .A(n122), .S(n31), .Y(n92) );
  INVX2 U73 ( .A(RX_CRC[10]), .Y(n46) );
  INVX2 U74 ( .A(cache_1[10]), .Y(n108) );
  MUX2X1 U75 ( .B(n46), .A(n108), .S(n31), .Y(n93) );
  INVX2 U76 ( .A(RX_CRC[11]), .Y(n47) );
  INVX2 U77 ( .A(cache_1[11]), .Y(n80) );
  MUX2X1 U78 ( .B(n47), .A(n80), .S(n31), .Y(n94) );
  INVX2 U79 ( .A(RX_CRC[12]), .Y(n48) );
  INVX2 U80 ( .A(cache_1[12]), .Y(n73) );
  MUX2X1 U81 ( .B(n48), .A(n73), .S(n31), .Y(n95) );
  INVX2 U82 ( .A(RX_CRC[13]), .Y(n49) );
  INVX2 U83 ( .A(cache_1[13]), .Y(n67) );
  MUX2X1 U84 ( .B(n49), .A(n67), .S(n31), .Y(n96) );
  INVX2 U85 ( .A(RX_CRC[14]), .Y(n50) );
  INVX2 U86 ( .A(cache_1[14]), .Y(n59) );
  MUX2X1 U87 ( .B(n50), .A(n59), .S(n31), .Y(n97) );
  INVX2 U88 ( .A(RX_CRC[15]), .Y(n51) );
  INVX2 U89 ( .A(cache_1[15]), .Y(n153) );
  MUX2X1 U90 ( .B(n51), .A(n153), .S(n31), .Y(n98) );
  INVX2 U91 ( .A(current_crc[7]), .Y(n58) );
  MUX2X1 U92 ( .B(n52), .A(n58), .S(n18), .Y(n99) );
  NAND2X1 U93 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n54) );
  INVX2 U94 ( .A(n161), .Y(n55) );
  XOR2X1 U95 ( .A(n63), .B(n55), .Y(n168) );
  INVX2 U96 ( .A(n168), .Y(n56) );
  NAND2X1 U97 ( .A(n20), .B(n56), .Y(n57) );
  OAI21X1 U98 ( .A(n29), .B(n58), .C(n57), .Y(n140) );
  INVX2 U99 ( .A(current_crc[14]), .Y(n61) );
  MUX2X1 U100 ( .B(n59), .A(n61), .S(n18), .Y(n101) );
  NAND2X1 U101 ( .A(current_crc[6]), .B(n20), .Y(n60) );
  OAI21X1 U102 ( .A(n30), .B(n61), .C(n60), .Y(n133) );
  INVX2 U103 ( .A(current_crc[6]), .Y(n66) );
  MUX2X1 U104 ( .B(n62), .A(n66), .S(n32), .Y(n103) );
  NAND2X1 U105 ( .A(n20), .B(n64), .Y(n65) );
  OAI21X1 U106 ( .A(n29), .B(n66), .C(n65), .Y(n141) );
  INVX2 U107 ( .A(current_crc[13]), .Y(n69) );
  MUX2X1 U108 ( .B(n67), .A(n69), .S(n18), .Y(n105) );
  NAND2X1 U109 ( .A(current_crc[5]), .B(n20), .Y(n68) );
  OAI21X1 U110 ( .A(n30), .B(n69), .C(n68), .Y(n134) );
  INVX2 U111 ( .A(current_crc[5]), .Y(n72) );
  MUX2X1 U112 ( .B(n70), .A(n72), .S(n32), .Y(n107) );
  NAND2X1 U113 ( .A(n20), .B(n1), .Y(n71) );
  OAI21X1 U114 ( .A(n29), .B(n72), .C(n71), .Y(n142) );
  INVX2 U115 ( .A(current_crc[12]), .Y(n75) );
  MUX2X1 U116 ( .B(n73), .A(n75), .S(n32), .Y(n109) );
  NAND2X1 U117 ( .A(current_crc[4]), .B(n20), .Y(n74) );
  OAI21X1 U118 ( .A(n30), .B(n75), .C(n74), .Y(n135) );
  INVX2 U119 ( .A(current_crc[4]), .Y(n79) );
  MUX2X1 U120 ( .B(n76), .A(n79), .S(n32), .Y(n111) );
  XOR2X1 U121 ( .A(n25), .B(n26), .Y(n77) );
  NAND2X1 U122 ( .A(n20), .B(n77), .Y(n78) );
  OAI21X1 U123 ( .A(n29), .B(n79), .C(n78), .Y(n143) );
  INVX2 U124 ( .A(current_crc[11]), .Y(n82) );
  MUX2X1 U125 ( .B(n80), .A(n82), .S(n32), .Y(n113) );
  NAND2X1 U126 ( .A(current_crc[3]), .B(n20), .Y(n81) );
  OAI21X1 U127 ( .A(n30), .B(n82), .C(n81), .Y(n136) );
  INVX2 U128 ( .A(current_crc[3]), .Y(n106) );
  MUX2X1 U129 ( .B(n100), .A(n106), .S(n32), .Y(n115) );
  XNOR2X1 U130 ( .A(n26), .B(n24), .Y(n131) );
  INVX2 U131 ( .A(n131), .Y(n102) );
  NAND2X1 U132 ( .A(n20), .B(n102), .Y(n104) );
  OAI21X1 U133 ( .A(n29), .B(n106), .C(n104), .Y(n144) );
  INVX2 U134 ( .A(current_crc[10]), .Y(n112) );
  MUX2X1 U135 ( .B(n108), .A(n112), .S(n18), .Y(n117) );
  NAND2X1 U136 ( .A(current_crc[2]), .B(n20), .Y(n110) );
  OAI21X1 U137 ( .A(n30), .B(n112), .C(n110), .Y(n137) );
  INVX2 U138 ( .A(current_crc[2]), .Y(n120) );
  MUX2X1 U139 ( .B(n114), .A(n120), .S(n32), .Y(n119) );
  XOR2X1 U140 ( .A(n23), .B(n24), .Y(n116) );
  NAND2X1 U141 ( .A(n20), .B(n116), .Y(n118) );
  OAI21X1 U142 ( .A(n29), .B(n120), .C(n118), .Y(n145) );
  INVX2 U143 ( .A(current_crc[9]), .Y(n128) );
  MUX2X1 U144 ( .B(n122), .A(n128), .S(n32), .Y(n121) );
  INVX2 U145 ( .A(n148), .Y(n166) );
  INVX2 U146 ( .A(current_crc[1]), .Y(n152) );
  XNOR2X1 U147 ( .A(n166), .B(n152), .Y(n124) );
  NAND2X1 U148 ( .A(n20), .B(n124), .Y(n126) );
  OAI21X1 U149 ( .A(n30), .B(n128), .C(n126), .Y(n138) );
  MUX2X1 U150 ( .B(n130), .A(n152), .S(n18), .Y(n123) );
  XOR2X1 U151 ( .A(n131), .B(n1), .Y(n167) );
  INVX2 U152 ( .A(n167), .Y(n156) );
  XNOR2X1 U153 ( .A(n168), .B(n148), .Y(n149) );
  XNOR2X1 U154 ( .A(n156), .B(n149), .Y(n150) );
  NAND2X1 U155 ( .A(n20), .B(n150), .Y(n151) );
  OAI21X1 U156 ( .A(n29), .B(n152), .C(n151), .Y(n146) );
  INVX2 U157 ( .A(current_crc[15]), .Y(n159) );
  MUX2X1 U158 ( .B(n153), .A(n159), .S(n18), .Y(n125) );
  FAX1 U159 ( .A(current_crc[7]), .B(n23), .C(n166), .YS(n154) );
  XNOR2X1 U160 ( .A(n154), .B(n168), .Y(n155) );
  XOR2X1 U161 ( .A(n156), .B(n155), .Y(n157) );
  NAND2X1 U162 ( .A(n20), .B(n157), .Y(n158) );
  OAI21X1 U163 ( .A(n30), .B(n159), .C(n158), .Y(n132) );
  INVX2 U164 ( .A(current_crc[8]), .Y(n164) );
  MUX2X1 U165 ( .B(n160), .A(n164), .S(n32), .Y(n127) );
  INVX2 U166 ( .A(current_crc[0]), .Y(n172) );
  FAX1 U167 ( .A(n166), .B(n172), .C(n161), .YS(n162) );
  NAND2X1 U168 ( .A(n20), .B(n162), .Y(n163) );
  OAI21X1 U169 ( .A(n29), .B(n164), .C(n163), .Y(n139) );
  MUX2X1 U170 ( .B(n165), .A(n172), .S(n18), .Y(n129) );
  XOR2X1 U171 ( .A(n23), .B(n166), .Y(n169) );
  FAX1 U172 ( .A(n169), .B(n168), .C(n167), .YS(n170) );
  NAND2X1 U173 ( .A(n20), .B(n170), .Y(n171) );
  OAI21X1 U174 ( .A(n30), .B(n172), .C(n171), .Y(n147) );
endmodule


module rx_accumulator_1 ( CLK, RST, RCV_DATA, W_ENABLE, rx_CHECK_CRC );
  input [7:0] RCV_DATA;
  output [15:0] rx_CHECK_CRC;
  input CLK, RST, W_ENABLE;
  wire   n3, n4, n6, n7, n9, n10, n12, n13, n15, n16, n18, n19, n21, n22, n24,
         n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51,
         n53, n55, n58, n1, n2, n5, n8, n11, n14, n17, n20, n23, n56, n59, n60
;

  DFFSR \present_CHECK_CRC_reg[7]  ( .D(n58), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[7]) );
  DFFSR \present_CHECK_CRC_reg[15]  ( .D(n55), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[15]) );
  DFFSR \present_CHECK_CRC_reg[6]  ( .D(n53), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[6]) );
  DFFSR \present_CHECK_CRC_reg[14]  ( .D(n51), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[14]) );
  DFFSR \present_CHECK_CRC_reg[5]  ( .D(n49), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[5]) );
  DFFSR \present_CHECK_CRC_reg[13]  ( .D(n47), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[13]) );
  DFFSR \present_CHECK_CRC_reg[4]  ( .D(n45), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[4]) );
  DFFSR \present_CHECK_CRC_reg[12]  ( .D(n43), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[12]) );
  DFFSR \present_CHECK_CRC_reg[3]  ( .D(n41), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[3]) );
  DFFSR \present_CHECK_CRC_reg[11]  ( .D(n39), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[11]) );
  DFFSR \present_CHECK_CRC_reg[2]  ( .D(n37), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[2]) );
  DFFSR \present_CHECK_CRC_reg[10]  ( .D(n35), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[10]) );
  DFFSR \present_CHECK_CRC_reg[1]  ( .D(n33), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[1]) );
  DFFSR \present_CHECK_CRC_reg[9]  ( .D(n31), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[9]) );
  DFFSR \present_CHECK_CRC_reg[0]  ( .D(n29), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[0]) );
  DFFSR \present_CHECK_CRC_reg[8]  ( .D(n27), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[8]) );
  OAI21X1 U2 ( .A(n8), .B(n60), .C(n3), .Y(n27) );
  NAND2X1 U3 ( .A(rx_CHECK_CRC[8]), .B(n8), .Y(n3) );
  OAI21X1 U4 ( .A(n2), .B(n60), .C(n4), .Y(n29) );
  NAND2X1 U5 ( .A(RCV_DATA[0]), .B(n2), .Y(n4) );
  OAI21X1 U7 ( .A(n8), .B(n59), .C(n6), .Y(n31) );
  NAND2X1 U8 ( .A(rx_CHECK_CRC[9]), .B(n8), .Y(n6) );
  OAI21X1 U9 ( .A(n2), .B(n59), .C(n7), .Y(n33) );
  NAND2X1 U10 ( .A(RCV_DATA[1]), .B(n2), .Y(n7) );
  OAI21X1 U12 ( .A(n8), .B(n56), .C(n9), .Y(n35) );
  NAND2X1 U13 ( .A(rx_CHECK_CRC[10]), .B(n8), .Y(n9) );
  OAI21X1 U14 ( .A(n2), .B(n56), .C(n10), .Y(n37) );
  NAND2X1 U15 ( .A(RCV_DATA[2]), .B(n2), .Y(n10) );
  OAI21X1 U17 ( .A(n8), .B(n23), .C(n12), .Y(n39) );
  NAND2X1 U18 ( .A(rx_CHECK_CRC[11]), .B(n8), .Y(n12) );
  OAI21X1 U19 ( .A(n2), .B(n23), .C(n13), .Y(n41) );
  NAND2X1 U20 ( .A(RCV_DATA[3]), .B(n2), .Y(n13) );
  OAI21X1 U22 ( .A(n8), .B(n20), .C(n15), .Y(n43) );
  NAND2X1 U23 ( .A(rx_CHECK_CRC[12]), .B(n8), .Y(n15) );
  OAI21X1 U24 ( .A(n2), .B(n20), .C(n16), .Y(n45) );
  NAND2X1 U25 ( .A(RCV_DATA[4]), .B(n2), .Y(n16) );
  OAI21X1 U27 ( .A(n8), .B(n17), .C(n18), .Y(n47) );
  NAND2X1 U28 ( .A(rx_CHECK_CRC[13]), .B(n8), .Y(n18) );
  OAI21X1 U29 ( .A(n2), .B(n17), .C(n19), .Y(n49) );
  NAND2X1 U30 ( .A(RCV_DATA[5]), .B(n2), .Y(n19) );
  OAI21X1 U32 ( .A(n8), .B(n14), .C(n21), .Y(n51) );
  NAND2X1 U33 ( .A(rx_CHECK_CRC[14]), .B(n8), .Y(n21) );
  OAI21X1 U34 ( .A(n2), .B(n14), .C(n22), .Y(n53) );
  NAND2X1 U35 ( .A(RCV_DATA[6]), .B(n2), .Y(n22) );
  OAI21X1 U37 ( .A(n8), .B(n11), .C(n24), .Y(n55) );
  NAND2X1 U38 ( .A(rx_CHECK_CRC[15]), .B(n8), .Y(n24) );
  OAI21X1 U41 ( .A(n2), .B(n11), .C(n25), .Y(n58) );
  NAND2X1 U42 ( .A(RCV_DATA[7]), .B(n2), .Y(n25) );
  INVX4 U6 ( .A(n2), .Y(n8) );
  INVX4 U11 ( .A(n1), .Y(n2) );
  INVX2 U16 ( .A(W_ENABLE), .Y(n1) );
  INVX2 U21 ( .A(RST), .Y(n5) );
  INVX2 U26 ( .A(rx_CHECK_CRC[7]), .Y(n11) );
  INVX2 U31 ( .A(rx_CHECK_CRC[6]), .Y(n14) );
  INVX2 U36 ( .A(rx_CHECK_CRC[5]), .Y(n17) );
  INVX2 U39 ( .A(rx_CHECK_CRC[4]), .Y(n20) );
  INVX2 U40 ( .A(rx_CHECK_CRC[3]), .Y(n23) );
  INVX2 U43 ( .A(rx_CHECK_CRC[2]), .Y(n56) );
  INVX2 U60 ( .A(rx_CHECK_CRC[1]), .Y(n59) );
  INVX2 U61 ( .A(rx_CHECK_CRC[0]), .Y(n60) );
endmodule


module rx_decode_1 ( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP, D_ORIG, BITSTUFF, 
        BS_ERROR );
  input CLK, RST, DP1_RX, SHIFT_ENABLE, EOP;
  output D_ORIG, BITSTUFF, BS_ERROR;
  wire   DP_hold1, DP_hold2, N29, N30, N31, N32, n17, n19, n43, n44, n2, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n18, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42;
  wire   [3:0] state;

  DFFSR DP_hold2_reg ( .D(n44), .CLK(CLK), .R(1'b1), .S(n9), .Q(DP_hold2) );
  DFFSR \state_reg[3]  ( .D(N32), .CLK(CLK), .R(n9), .S(1'b1), .Q(state[3]) );
  DFFSR DP_hold1_reg ( .D(n43), .CLK(CLK), .R(1'b1), .S(n9), .Q(DP_hold1) );
  NAND2X1 U20 ( .A(n17), .B(n41), .Y(n43) );
  AOI22X1 U21 ( .A(DP_hold1), .B(n42), .C(DP1_RX), .D(n19), .Y(n17) );
  XNOR2X1 U25 ( .A(DP_hold1), .B(DP_hold2), .Y(D_ORIG) );
  DFFSR \state_reg[0]  ( .D(N29), .CLK(CLK), .R(n9), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[2]  ( .D(N31), .CLK(CLK), .R(n9), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[1]  ( .D(N30), .CLK(CLK), .R(n9), .S(1'b1), .Q(state[1]) );
  AND2X2 U4 ( .A(state[1]), .B(state[2]), .Y(n2) );
  INVX1 U10 ( .A(SHIFT_ENABLE), .Y(n31) );
  AND2X1 U11 ( .A(SHIFT_ENABLE), .B(state[0]), .Y(n22) );
  INVX2 U12 ( .A(RST), .Y(n9) );
  MUX2X1 U13 ( .B(DP_hold1), .A(DP_hold2), .S(n8), .Y(n40) );
  NAND2X1 U14 ( .A(SHIFT_ENABLE), .B(n19), .Y(n8) );
  INVX2 U15 ( .A(state[0]), .Y(n15) );
  NOR2X1 U16 ( .A(state[1]), .B(state[2]), .Y(n10) );
  NAND3X1 U17 ( .A(state[3]), .B(n15), .C(n10), .Y(n11) );
  INVX2 U18 ( .A(n11), .Y(BS_ERROR) );
  NAND2X1 U19 ( .A(n2), .B(n15), .Y(n19) );
  NOR2X1 U22 ( .A(state[3]), .B(n19), .Y(BITSTUFF) );
  INVX2 U23 ( .A(n19), .Y(n42) );
  OR2X2 U24 ( .A(EOP), .B(state[3]), .Y(n37) );
  INVX2 U26 ( .A(n37), .Y(n41) );
  INVX2 U27 ( .A(DP1_RX), .Y(n12) );
  XOR2X1 U28 ( .A(n12), .B(DP_hold2), .Y(n33) );
  INVX2 U29 ( .A(n33), .Y(n24) );
  NOR2X1 U30 ( .A(state[0]), .B(n24), .Y(n13) );
  MUX2X1 U31 ( .B(n13), .A(n24), .S(n2), .Y(n14) );
  MUX2X1 U32 ( .B(n15), .A(n14), .S(SHIFT_ENABLE), .Y(n16) );
  AND2X2 U33 ( .A(n41), .B(n16), .Y(N29) );
  INVX2 U34 ( .A(state[2]), .Y(n18) );
  NAND3X1 U35 ( .A(state[1]), .B(n33), .C(n18), .Y(n35) );
  INVX2 U36 ( .A(n35), .Y(n23) );
  INVX2 U37 ( .A(state[1]), .Y(n32) );
  NAND2X1 U38 ( .A(n33), .B(n32), .Y(n20) );
  AOI21X1 U39 ( .A(SHIFT_ENABLE), .B(n20), .C(n18), .Y(n21) );
  AOI21X1 U40 ( .A(n23), .B(n22), .C(n21), .Y(n25) );
  NAND2X1 U41 ( .A(n24), .B(n42), .Y(n29) );
  AOI21X1 U42 ( .A(n25), .B(n29), .C(n37), .Y(N31) );
  NAND3X1 U43 ( .A(n33), .B(n42), .C(SHIFT_ENABLE), .Y(n28) );
  INVX2 U44 ( .A(EOP), .Y(n26) );
  NAND2X1 U45 ( .A(BS_ERROR), .B(n26), .Y(n27) );
  OAI21X1 U46 ( .A(n37), .B(n28), .C(n27), .Y(N32) );
  INVX2 U47 ( .A(n29), .Y(n30) );
  AOI21X1 U48 ( .A(state[1]), .B(n31), .C(n30), .Y(n39) );
  NAND3X1 U49 ( .A(SHIFT_ENABLE), .B(n33), .C(n32), .Y(n34) );
  MUX2X1 U50 ( .B(n35), .A(n34), .S(state[0]), .Y(n36) );
  INVX2 U51 ( .A(n36), .Y(n38) );
  AOI21X1 U52 ( .A(n39), .B(n38), .C(n37), .Y(N30) );
  NAND2X1 U53 ( .A(n41), .B(n40), .Y(n44) );
endmodule


module rx_edgedetect_1 ( CLK, RST, DP1_RX, D_EDGE );
  input CLK, RST, DP1_RX;
  output D_EDGE;
  wire   DP_hold1, DP_hold2, n2, n4;

  DFFSR DP_hold1_reg ( .D(DP1_RX), .CLK(CLK), .R(1'b1), .S(n2), .Q(DP_hold1)
         );
  DFFSR DP_hold2_reg ( .D(DP_hold1), .CLK(CLK), .R(1'b1), .S(n2), .Q(DP_hold2)
         );
  INVX2 U4 ( .A(RST), .Y(n2) );
  XNOR2X1 U6 ( .A(DP_hold2), .B(DP_hold1), .Y(n4) );
  NOR2X1 U7 ( .A(RST), .B(n4), .Y(D_EDGE) );
endmodule


module rx_eopdetect_1 ( DP1_RX, DM1_RX, EOP );
  input DP1_RX, DM1_RX;
  output EOP;


  NOR2X1 U1 ( .A(DP1_RX), .B(DM1_RX), .Y(EOP) );
endmodule


module rx_rcu_1 ( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR, 
        RX_CRC, RX_CHECK_CRC, RCV_DATA, RCVING, W_ENABLE, R_ERROR, CRC_ERROR, 
        OPCODE );
  input [15:0] RX_CRC;
  input [15:0] RX_CHECK_CRC;
  input [7:0] RCV_DATA;
  output [1:0] OPCODE;
  input CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR;
  output RCVING, W_ENABLE, R_ERROR, CRC_ERROR;
  wire   nxtR_ERROR, curR_ERROR, curCRC_ERROR, N170, n37, n38, n41, n42, n83,
         n87, n88, n94, n150, n151, n161, n162, n163, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n39, n40,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84, n85,
         n86, n89, n90, n91, n92, n93, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n153, n154, n157, n160, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223;
  wire   [3:0] state;
  wire   [3:0] count;
  wire   [3:0] nextstate;

  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(CLK), .R(n51), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(CLK), .R(n51), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(CLK), .R(n51), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(CLK), .R(n51), .S(1'b1), .Q(
        state[1]) );
  DFFSR \count_reg[3]  ( .D(n163), .CLK(CLK), .R(n51), .S(1'b1), .Q(count[3])
         );
  DFFPOSX1 curCRC_ERROR_reg ( .D(n151), .CLK(CLK), .Q(curCRC_ERROR) );
  DFFPOSX1 curR_ERROR_reg ( .D(n150), .CLK(CLK), .Q(curR_ERROR) );
  DFFSR R_ERROR_reg ( .D(nxtR_ERROR), .CLK(CLK), .R(n51), .S(1'b1), .Q(R_ERROR) );
  DFFPOSX1 CRC_ERROR_reg ( .D(n218), .CLK(CLK), .Q(CRC_ERROR) );
  NAND2X1 U16 ( .A(n37), .B(n38), .Y(nextstate[2]) );
  OAI21X1 U19 ( .A(n222), .B(n42), .C(n47), .Y(n41) );
  NAND2X1 U20 ( .A(n184), .B(n185), .Y(n42) );
  AOI21X1 U52 ( .A(CRC_ERROR), .B(RST), .C(n88), .Y(n87) );
  OAI21X1 U56 ( .A(n51), .B(n220), .C(n94), .Y(n150) );
  NOR2X1 U79 ( .A(D_EDGE), .B(n49), .Y(n83) );
  DFFSR \count_reg[0]  ( .D(n217), .CLK(CLK), .R(n51), .S(1'b1), .Q(count[0])
         );
  DFFSR \count_reg[1]  ( .D(n161), .CLK(CLK), .R(n51), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n162), .CLK(CLK), .R(n51), .S(1'b1), .Q(count[2])
         );
  AND2X2 U3 ( .A(n5), .B(n48), .Y(n1) );
  AND2X1 U4 ( .A(n65), .B(n129), .Y(n2) );
  BUFX2 U5 ( .A(n39), .Y(n3) );
  BUFX2 U6 ( .A(n35), .Y(n4) );
  BUFX4 U7 ( .A(state[1]), .Y(n5) );
  AND2X2 U8 ( .A(n168), .B(n85), .Y(n6) );
  AND2X2 U9 ( .A(n19), .B(n35), .Y(n7) );
  AND2X2 U10 ( .A(n50), .B(n166), .Y(n8) );
  INVX2 U11 ( .A(n14), .Y(n170) );
  AND2X1 U12 ( .A(n70), .B(n16), .Y(n9) );
  AND2X2 U13 ( .A(n21), .B(n7), .Y(n10) );
  INVX2 U18 ( .A(n48), .Y(n14) );
  INVX4 U21 ( .A(n48), .Y(n49) );
  NAND2X1 U22 ( .A(n5), .B(n170), .Y(n15) );
  BUFX2 U23 ( .A(n129), .Y(n16) );
  BUFX2 U24 ( .A(n5), .Y(n47) );
  BUFX2 U25 ( .A(n46), .Y(n17) );
  AND2X2 U26 ( .A(n5), .B(n14), .Y(n52) );
  BUFX2 U27 ( .A(n33), .Y(n18) );
  NAND2X1 U28 ( .A(n32), .B(n2), .Y(W_ENABLE) );
  AND2X2 U29 ( .A(n64), .B(n63), .Y(n19) );
  INVX1 U30 ( .A(n19), .Y(n135) );
  INVX1 U31 ( .A(n54), .Y(n20) );
  BUFX2 U32 ( .A(n1), .Y(n21) );
  INVX4 U33 ( .A(n50), .Y(n54) );
  NAND2X1 U34 ( .A(n21), .B(n8), .Y(n22) );
  NAND2X1 U35 ( .A(n1), .B(n8), .Y(n123) );
  NAND2X1 U36 ( .A(n24), .B(n9), .Y(RCVING) );
  INVX2 U37 ( .A(n175), .Y(n23) );
  AND2X2 U38 ( .A(n25), .B(n43), .Y(n24) );
  INVX1 U39 ( .A(n24), .Y(n90) );
  NOR2X1 U40 ( .A(n36), .B(n23), .Y(n25) );
  NAND2X1 U41 ( .A(n1), .B(n7), .Y(n179) );
  AND2X2 U42 ( .A(SHIFT_ENABLE), .B(n103), .Y(n26) );
  AND2X1 U43 ( .A(n111), .B(n115), .Y(n112) );
  BUFX4 U44 ( .A(state[3]), .Y(n39) );
  AND2X1 U45 ( .A(n46), .B(n54), .Y(n27) );
  INVX1 U46 ( .A(n47), .Y(n73) );
  INVX2 U47 ( .A(n125), .Y(n28) );
  AND2X2 U48 ( .A(n39), .B(n50), .Y(n29) );
  INVX1 U49 ( .A(n29), .Y(n153) );
  NAND2X1 U50 ( .A(n65), .B(n129), .Y(OPCODE[0]) );
  AND2X1 U51 ( .A(n118), .B(n115), .Y(n31) );
  OR2X1 U53 ( .A(RCV_DATA[1]), .B(RCV_DATA[2]), .Y(n60) );
  AND2X2 U54 ( .A(n68), .B(n179), .Y(n32) );
  INVX2 U55 ( .A(RST), .Y(n51) );
  AND2X2 U57 ( .A(n39), .B(n54), .Y(n33) );
  AND2X2 U58 ( .A(SHIFT_ENABLE), .B(n103), .Y(n34) );
  NOR2X1 U59 ( .A(n50), .B(n39), .Y(n35) );
  NAND2X1 U60 ( .A(n69), .B(n68), .Y(n36) );
  INVX1 U61 ( .A(n111), .Y(n107) );
  INVX1 U62 ( .A(n105), .Y(n110) );
  INVX1 U63 ( .A(n67), .Y(n40) );
  INVX1 U64 ( .A(n40), .Y(n43) );
  INVX2 U65 ( .A(n71), .Y(n44) );
  INVX1 U66 ( .A(n8), .Y(n45) );
  AND2X2 U67 ( .A(state[2]), .B(n166), .Y(n46) );
  INVX1 U68 ( .A(n17), .Y(n71) );
  BUFX4 U69 ( .A(state[0]), .Y(n50) );
  INVX1 U70 ( .A(n178), .Y(n125) );
  INVX2 U71 ( .A(state[2]), .Y(n48) );
  INVX1 U72 ( .A(n167), .Y(n168) );
  INVX2 U73 ( .A(state[3]), .Y(n166) );
  NAND2X1 U74 ( .A(n52), .B(n8), .Y(n129) );
  NAND2X1 U75 ( .A(n17), .B(n54), .Y(n167) );
  NAND2X1 U76 ( .A(n27), .B(n47), .Y(n65) );
  INVX2 U77 ( .A(n5), .Y(n172) );
  NOR2X1 U78 ( .A(n49), .B(n172), .Y(n53) );
  NAND2X1 U80 ( .A(n53), .B(n29), .Y(n178) );
  NAND2X1 U81 ( .A(n178), .B(n123), .Y(n89) );
  INVX2 U82 ( .A(n89), .Y(n67) );
  NAND2X1 U83 ( .A(n33), .B(n49), .Y(n56) );
  OAI21X1 U84 ( .A(n50), .B(n170), .C(n166), .Y(n55) );
  MUX2X1 U85 ( .B(n56), .A(n55), .S(n47), .Y(n57) );
  NAND2X1 U86 ( .A(n57), .B(n67), .Y(OPCODE[1]) );
  NAND3X1 U87 ( .A(n33), .B(n49), .C(n172), .Y(n68) );
  INVX2 U88 ( .A(RCV_DATA[0]), .Y(n58) );
  NAND2X1 U89 ( .A(RCV_DATA[7]), .B(n58), .Y(n59) );
  NOR2X1 U90 ( .A(n60), .B(n59), .Y(n64) );
  NOR2X1 U91 ( .A(RCV_DATA[4]), .B(RCV_DATA[3]), .Y(n62) );
  NOR2X1 U92 ( .A(RCV_DATA[6]), .B(RCV_DATA[5]), .Y(n61) );
  AND2X2 U93 ( .A(n62), .B(n61), .Y(n63) );
  NAND3X1 U94 ( .A(n29), .B(n49), .C(n172), .Y(n177) );
  OAI21X1 U95 ( .A(n47), .B(n167), .C(n177), .Y(n121) );
  INVX2 U96 ( .A(n121), .Y(n70) );
  NOR2X1 U97 ( .A(n39), .B(n49), .Y(n66) );
  NAND3X1 U98 ( .A(n66), .B(n50), .C(n172), .Y(n175) );
  NAND2X1 U99 ( .A(n43), .B(n175), .Y(n104) );
  NAND2X1 U100 ( .A(n1), .B(n166), .Y(n69) );
  NAND2X1 U101 ( .A(n83), .B(n18), .Y(n81) );
  NAND2X1 U102 ( .A(n81), .B(n71), .Y(n72) );
  NAND3X1 U103 ( .A(curR_ERROR), .B(n73), .C(n72), .Y(n79) );
  NOR2X1 U104 ( .A(n20), .B(n15), .Y(n75) );
  NAND2X1 U105 ( .A(n19), .B(n166), .Y(n74) );
  NAND2X1 U106 ( .A(n75), .B(n74), .Y(n96) );
  NAND2X1 U107 ( .A(n28), .B(n175), .Y(n77) );
  NOR2X1 U108 ( .A(count[3]), .B(n172), .Y(n76) );
  NOR3X1 U109 ( .A(count[0]), .B(count[1]), .C(count[2]), .Y(n184) );
  NAND2X1 U110 ( .A(n76), .B(n184), .Y(n84) );
  AOI22X1 U111 ( .A(EOP), .B(n77), .C(n168), .D(n84), .Y(n78) );
  NAND3X1 U112 ( .A(n79), .B(n96), .C(n78), .Y(nxtR_ERROR) );
  INVX2 U113 ( .A(n79), .Y(n80) );
  OAI21X1 U114 ( .A(n51), .B(n80), .C(nxtR_ERROR), .Y(n94) );
  NAND2X1 U115 ( .A(curCRC_ERROR), .B(n51), .Y(n86) );
  NAND2X1 U116 ( .A(n8), .B(n49), .Y(n91) );
  NAND2X1 U117 ( .A(n91), .B(n81), .Y(n82) );
  NAND2X1 U118 ( .A(n82), .B(n172), .Y(n99) );
  INVX2 U119 ( .A(n84), .Y(n85) );
  NAND3X1 U120 ( .A(n222), .B(n51), .C(n6), .Y(n102) );
  OAI21X1 U121 ( .A(n86), .B(n99), .C(n102), .Y(n88) );
  INVX2 U122 ( .A(count[3]), .Y(n185) );
  NAND2X1 U123 ( .A(n184), .B(count[3]), .Y(n124) );
  INVX2 U124 ( .A(n124), .Y(n122) );
  AOI22X1 U125 ( .A(n90), .B(BS_ERROR), .C(n122), .D(n89), .Y(n95) );
  OAI22X1 U126 ( .A(n167), .B(EOP), .C(D_EDGE), .D(n91), .Y(n92) );
  MUX2X1 U127 ( .B(n92), .A(n18), .S(n47), .Y(n93) );
  AND2X2 U128 ( .A(n95), .B(n93), .Y(n37) );
  OAI21X1 U129 ( .A(n41), .B(n167), .C(n96), .Y(n98) );
  NAND2X1 U130 ( .A(EOP), .B(n104), .Y(n115) );
  NAND2X1 U131 ( .A(n115), .B(n177), .Y(n97) );
  NOR2X1 U132 ( .A(n98), .B(n97), .Y(n38) );
  INVX2 U133 ( .A(n99), .Y(n100) );
  OAI21X1 U134 ( .A(RST), .B(n100), .C(curCRC_ERROR), .Y(n101) );
  NAND2X1 U135 ( .A(n102), .B(n101), .Y(n151) );
  INVX2 U136 ( .A(BITSTUFF), .Y(n103) );
  NAND3X1 U137 ( .A(count[1]), .B(count[0]), .C(n34), .Y(n105) );
  NAND2X1 U138 ( .A(n104), .B(n124), .Y(n116) );
  INVX2 U139 ( .A(n116), .Y(n118) );
  NAND3X1 U140 ( .A(n110), .B(n31), .C(count[2]), .Y(n109) );
  NAND2X1 U141 ( .A(n118), .B(n105), .Y(n111) );
  OAI21X1 U142 ( .A(count[2]), .B(n116), .C(n115), .Y(n106) );
  NOR2X1 U143 ( .A(n107), .B(n106), .Y(n108) );
  MUX2X1 U144 ( .B(n109), .A(n108), .S(count[3]), .Y(n163) );
  NAND2X1 U145 ( .A(n31), .B(n110), .Y(n113) );
  MUX2X1 U146 ( .B(n113), .A(n112), .S(count[2]), .Y(n162) );
  NAND3X1 U147 ( .A(n26), .B(n118), .C(n115), .Y(n134) );
  INVX2 U148 ( .A(n134), .Y(n114) );
  NAND2X1 U149 ( .A(count[0]), .B(n114), .Y(n120) );
  INVX2 U150 ( .A(count[0]), .Y(n117) );
  OAI21X1 U151 ( .A(n26), .B(n116), .C(n115), .Y(n132) );
  AOI21X1 U152 ( .A(n118), .B(n117), .C(n132), .Y(n119) );
  MUX2X1 U153 ( .B(n120), .A(n119), .S(count[1]), .Y(n161) );
  NAND2X1 U154 ( .A(n121), .B(EOP), .Y(n131) );
  NAND2X1 U155 ( .A(n122), .B(n223), .Y(n140) );
  OAI21X1 U156 ( .A(n140), .B(n175), .C(n22), .Y(n128) );
  NAND3X1 U157 ( .A(n223), .B(n125), .C(n124), .Y(n126) );
  NAND2X1 U158 ( .A(n32), .B(n126), .Y(n127) );
  OAI21X1 U159 ( .A(n128), .B(n127), .C(n221), .Y(n130) );
  NAND3X1 U162 ( .A(n131), .B(n130), .C(n16), .Y(nextstate[1]) );
  INVX2 U163 ( .A(n132), .Y(n133) );
  MUX2X1 U166 ( .B(n134), .A(n133), .S(count[0]), .Y(n217) );
  NOR2X1 U169 ( .A(n223), .B(n45), .Y(n138) );
  NAND2X1 U170 ( .A(n4), .B(n135), .Y(n136) );
  OAI21X1 U171 ( .A(n153), .B(n140), .C(n136), .Y(n137) );
  OAI21X1 U172 ( .A(n138), .B(n137), .C(n221), .Y(n139) );
  NAND2X1 U173 ( .A(n1), .B(n139), .Y(n165) );
  NAND2X1 U174 ( .A(n29), .B(D_EDGE), .Y(n143) );
  INVX2 U175 ( .A(n140), .Y(n141) );
  NAND3X1 U176 ( .A(n8), .B(n141), .C(n221), .Y(n142) );
  NAND2X1 U177 ( .A(n143), .B(n142), .Y(n145) );
  NOR2X1 U178 ( .A(n153), .B(n223), .Y(n144) );
  MUX2X1 U179 ( .B(n145), .A(n144), .S(n49), .Y(n148) );
  OR2X2 U180 ( .A(n219), .B(n20), .Y(n147) );
  AOI21X1 U181 ( .A(D_EDGE), .B(n44), .C(n168), .Y(n146) );
  NAND3X1 U182 ( .A(n148), .B(n147), .C(n146), .Y(n157) );
  NAND2X1 U183 ( .A(n49), .B(n153), .Y(n154) );
  MUX2X1 U184 ( .B(n157), .A(n154), .S(n47), .Y(n160) );
  INVX2 U185 ( .A(n160), .Y(n164) );
  NAND2X1 U186 ( .A(n165), .B(n164), .Y(nextstate[0]) );
  NOR2X1 U187 ( .A(n219), .B(n166), .Y(n174) );
  AOI22X1 U188 ( .A(n3), .B(BS_ERROR), .C(D_EDGE), .D(n20), .Y(n171) );
  NAND2X1 U189 ( .A(n168), .B(EOP), .Y(n169) );
  OAI21X1 U190 ( .A(n171), .B(n170), .C(n169), .Y(n173) );
  OAI21X1 U191 ( .A(n174), .B(n173), .C(n172), .Y(n183) );
  OAI21X1 U192 ( .A(n18), .B(n15), .C(n175), .Y(n176) );
  AOI22X1 U193 ( .A(n6), .B(N170), .C(BS_ERROR), .D(n176), .Y(n182) );
  OAI21X1 U194 ( .A(EOP), .B(n28), .C(n177), .Y(n180) );
  NOR2X1 U195 ( .A(n180), .B(n10), .Y(n181) );
  NAND3X1 U196 ( .A(n183), .B(n182), .C(n181), .Y(nextstate[3]) );
  XNOR2X1 U197 ( .A(RX_CHECK_CRC[10]), .B(RX_CRC[10]), .Y(n190) );
  XNOR2X1 U198 ( .A(RX_CHECK_CRC[9]), .B(RX_CRC[9]), .Y(n189) );
  XOR2X1 U199 ( .A(RX_CHECK_CRC[7]), .B(RX_CRC[7]), .Y(n187) );
  XOR2X1 U200 ( .A(RX_CHECK_CRC[8]), .B(RX_CRC[8]), .Y(n186) );
  NOR2X1 U201 ( .A(n187), .B(n186), .Y(n188) );
  NAND3X1 U202 ( .A(n190), .B(n189), .C(n188), .Y(n197) );
  XNOR2X1 U203 ( .A(RX_CHECK_CRC[14]), .B(RX_CRC[14]), .Y(n195) );
  XNOR2X1 U204 ( .A(RX_CHECK_CRC[13]), .B(RX_CRC[13]), .Y(n194) );
  XOR2X1 U205 ( .A(RX_CHECK_CRC[11]), .B(RX_CRC[11]), .Y(n192) );
  XOR2X1 U206 ( .A(RX_CHECK_CRC[12]), .B(RX_CRC[12]), .Y(n191) );
  NOR2X1 U207 ( .A(n192), .B(n191), .Y(n193) );
  NAND3X1 U208 ( .A(n195), .B(n194), .C(n193), .Y(n196) );
  NOR2X1 U209 ( .A(n197), .B(n196), .Y(n213) );
  NOR2X1 U210 ( .A(n214), .B(RX_CHECK_CRC[0]), .Y(n198) );
  OAI22X1 U211 ( .A(RX_CRC[1]), .B(n198), .C(n198), .D(n216), .Y(n204) );
  AND2X1 U212 ( .A(RX_CHECK_CRC[0]), .B(n214), .Y(n199) );
  OAI22X1 U213 ( .A(n199), .B(n215), .C(RX_CHECK_CRC[1]), .D(n199), .Y(n203)
         );
  XOR2X1 U214 ( .A(RX_CHECK_CRC[15]), .B(RX_CRC[15]), .Y(n201) );
  XOR2X1 U215 ( .A(RX_CHECK_CRC[2]), .B(RX_CRC[2]), .Y(n200) );
  NOR2X1 U216 ( .A(n201), .B(n200), .Y(n202) );
  NAND3X1 U217 ( .A(n204), .B(n203), .C(n202), .Y(n211) );
  XNOR2X1 U218 ( .A(RX_CHECK_CRC[6]), .B(RX_CRC[6]), .Y(n209) );
  XNOR2X1 U219 ( .A(RX_CHECK_CRC[5]), .B(RX_CRC[5]), .Y(n208) );
  XOR2X1 U220 ( .A(RX_CHECK_CRC[3]), .B(RX_CRC[3]), .Y(n206) );
  XOR2X1 U221 ( .A(RX_CHECK_CRC[4]), .B(RX_CRC[4]), .Y(n205) );
  NOR2X1 U222 ( .A(n206), .B(n205), .Y(n207) );
  NAND3X1 U223 ( .A(n209), .B(n208), .C(n207), .Y(n210) );
  NOR2X1 U224 ( .A(n211), .B(n210), .Y(n212) );
  AND2X1 U225 ( .A(n213), .B(n212), .Y(N170) );
  INVX2 U226 ( .A(RX_CRC[0]), .Y(n214) );
  INVX2 U227 ( .A(RX_CRC[1]), .Y(n215) );
  INVX2 U228 ( .A(RX_CHECK_CRC[1]), .Y(n216) );
  INVX2 U229 ( .A(n87), .Y(n218) );
  INVX2 U230 ( .A(n83), .Y(n219) );
  INVX2 U231 ( .A(curR_ERROR), .Y(n220) );
  INVX2 U232 ( .A(BS_ERROR), .Y(n221) );
  INVX2 U233 ( .A(N170), .Y(n222) );
  INVX2 U234 ( .A(EOP), .Y(n223) );
endmodule


module rx_shift_reg_1 ( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF, RCV_DATA );
  output [7:0] RCV_DATA;
  input CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF;
  wire   n2, n6, n8, n10, n12, n14, n16, n18, n21, n23, n24, n26, n27, n29,
         n30, n32, n33, n35, n36, n38, n39, n41, n42, n44, n15, n17, n19, n20,
         n22, n25, n28, n31, n34, n37, n40, n43, n45, n46, n47, n48, n49, n50;
  wire   [7:0] present_val;

  DFFPOSX1 \RCV_DATA_reg[7]  ( .D(n42), .CLK(CLK), .Q(RCV_DATA[7]) );
  DFFPOSX1 \RCV_DATA_reg[6]  ( .D(n39), .CLK(CLK), .Q(RCV_DATA[6]) );
  DFFPOSX1 \RCV_DATA_reg[5]  ( .D(n36), .CLK(CLK), .Q(RCV_DATA[5]) );
  DFFPOSX1 \RCV_DATA_reg[4]  ( .D(n33), .CLK(CLK), .Q(RCV_DATA[4]) );
  DFFPOSX1 \RCV_DATA_reg[3]  ( .D(n30), .CLK(CLK), .Q(RCV_DATA[3]) );
  DFFPOSX1 \RCV_DATA_reg[2]  ( .D(n27), .CLK(CLK), .Q(RCV_DATA[2]) );
  DFFPOSX1 \RCV_DATA_reg[1]  ( .D(n24), .CLK(CLK), .Q(RCV_DATA[1]) );
  DFFPOSX1 \RCV_DATA_reg[0]  ( .D(n21), .CLK(CLK), .Q(RCV_DATA[0]) );
  OAI21X1 U2 ( .A(RST), .B(n50), .C(n2), .Y(n21) );
  NAND2X1 U3 ( .A(RCV_DATA[0]), .B(RST), .Y(n2) );
  OAI21X1 U6 ( .A(RST), .B(n49), .C(n6), .Y(n24) );
  NAND2X1 U7 ( .A(RCV_DATA[1]), .B(RST), .Y(n6) );
  OAI21X1 U10 ( .A(RST), .B(n48), .C(n8), .Y(n27) );
  NAND2X1 U11 ( .A(n25), .B(RST), .Y(n8) );
  OAI21X1 U14 ( .A(RST), .B(n47), .C(n10), .Y(n30) );
  NAND2X1 U15 ( .A(RCV_DATA[3]), .B(RST), .Y(n10) );
  OAI21X1 U18 ( .A(RST), .B(n46), .C(n12), .Y(n33) );
  NAND2X1 U19 ( .A(RCV_DATA[4]), .B(RST), .Y(n12) );
  OAI21X1 U22 ( .A(RST), .B(n45), .C(n14), .Y(n36) );
  NAND2X1 U23 ( .A(RCV_DATA[5]), .B(RST), .Y(n14) );
  OAI21X1 U26 ( .A(RST), .B(n43), .C(n16), .Y(n39) );
  NAND2X1 U27 ( .A(n17), .B(RST), .Y(n16) );
  OAI21X1 U30 ( .A(RST), .B(n40), .C(n18), .Y(n42) );
  NAND2X1 U31 ( .A(n20), .B(RST), .Y(n18) );
  DFFSR \present_val_reg[0]  ( .D(n23), .CLK(CLK), .R(n31), .S(1'b1), .Q(
        present_val[0]) );
  DFFSR \present_val_reg[7]  ( .D(n44), .CLK(CLK), .R(n31), .S(1'b1), .Q(
        present_val[7]) );
  DFFSR \present_val_reg[6]  ( .D(n41), .CLK(CLK), .R(n31), .S(1'b1), .Q(
        present_val[6]) );
  DFFSR \present_val_reg[5]  ( .D(n38), .CLK(CLK), .R(n31), .S(1'b1), .Q(
        present_val[5]) );
  DFFSR \present_val_reg[4]  ( .D(n35), .CLK(CLK), .R(n31), .S(1'b1), .Q(
        present_val[4]) );
  DFFSR \present_val_reg[3]  ( .D(n32), .CLK(CLK), .R(n31), .S(1'b1), .Q(
        present_val[3]) );
  DFFSR \present_val_reg[2]  ( .D(n29), .CLK(CLK), .R(n31), .S(1'b1), .Q(
        present_val[2]) );
  DFFSR \present_val_reg[1]  ( .D(n26), .CLK(CLK), .R(n31), .S(1'b1), .Q(
        present_val[1]) );
  INVX1 U20 ( .A(RCV_DATA[6]), .Y(n15) );
  INVX2 U21 ( .A(n15), .Y(n17) );
  INVX1 U24 ( .A(RCV_DATA[7]), .Y(n19) );
  INVX2 U25 ( .A(n19), .Y(n20) );
  INVX1 U28 ( .A(RCV_DATA[2]), .Y(n22) );
  INVX2 U29 ( .A(n22), .Y(n25) );
  INVX2 U32 ( .A(RST), .Y(n31) );
  AND2X2 U33 ( .A(SHIFT_ENABLE), .B(n34), .Y(n28) );
  INVX2 U34 ( .A(present_val[7]), .Y(n40) );
  INVX2 U35 ( .A(present_val[6]), .Y(n43) );
  INVX2 U36 ( .A(present_val[5]), .Y(n45) );
  INVX2 U37 ( .A(present_val[4]), .Y(n46) );
  INVX2 U38 ( .A(present_val[3]), .Y(n47) );
  INVX2 U39 ( .A(present_val[2]), .Y(n48) );
  INVX2 U40 ( .A(present_val[1]), .Y(n49) );
  INVX2 U41 ( .A(present_val[0]), .Y(n50) );
  INVX2 U42 ( .A(BITSTUFF), .Y(n34) );
  MUX2X1 U43 ( .B(n50), .A(n49), .S(n28), .Y(n23) );
  MUX2X1 U44 ( .B(n49), .A(n48), .S(n28), .Y(n26) );
  MUX2X1 U45 ( .B(n48), .A(n47), .S(n28), .Y(n29) );
  MUX2X1 U46 ( .B(n47), .A(n46), .S(n28), .Y(n32) );
  MUX2X1 U47 ( .B(n46), .A(n45), .S(n28), .Y(n35) );
  MUX2X1 U48 ( .B(n45), .A(n43), .S(n28), .Y(n38) );
  MUX2X1 U49 ( .B(n43), .A(n40), .S(n28), .Y(n41) );
  INVX2 U50 ( .A(D_ORIG), .Y(n37) );
  MUX2X1 U51 ( .B(n40), .A(n37), .S(n28), .Y(n44) );
endmodule


module rx_timer_1 ( CLK, RST, D_EDGE, RCVING, SHIFT_ENABLE );
  input CLK, RST, D_EDGE, RCVING;
  output SHIFT_ENABLE;
  wire   state, n15, n17, n18, n20, n21, n22, n23, n5, n7, n8, n9, n10, n11,
         n12, n13, n14, n16, n19, n24, n25, n26, n27;
  wire   [3:0] count;
  wire   [3:0] nextcount;

  DFFSR state_reg ( .D(n11), .CLK(CLK), .R(n12), .S(1'b1), .Q(state) );
  DFFSR \count_reg[0]  ( .D(nextcount[0]), .CLK(CLK), .R(n12), .S(1'b1), .Q(
        count[0]) );
  DFFSR \count_reg[1]  ( .D(nextcount[1]), .CLK(CLK), .R(n12), .S(1'b1), .Q(
        count[1]) );
  DFFSR \count_reg[2]  ( .D(nextcount[2]), .CLK(CLK), .R(n12), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[3]  ( .D(nextcount[3]), .CLK(CLK), .R(n12), .S(1'b1), .Q(
        count[3]) );
  XOR2X1 U19 ( .A(n18), .B(n25), .Y(n17) );
  NOR2X1 U20 ( .A(count[3]), .B(n26), .Y(n15) );
  XOR2X1 U22 ( .A(n21), .B(count[2]), .Y(n20) );
  NAND2X1 U24 ( .A(state), .B(n23), .Y(nextcount[0]) );
  OAI21X1 U25 ( .A(D_EDGE), .B(n27), .C(n11), .Y(n23) );
  NAND2X1 U30 ( .A(count[0]), .B(count[1]), .Y(n21) );
  XNOR2X1 U32 ( .A(count[0]), .B(count[1]), .Y(n22) );
  INVX2 U7 ( .A(n10), .Y(SHIFT_ENABLE) );
  INVX1 U9 ( .A(n7), .Y(nextcount[2]) );
  INVX2 U10 ( .A(RST), .Y(n12) );
  NOR2X1 U11 ( .A(n16), .B(n25), .Y(n5) );
  OAI21X1 U12 ( .A(n8), .B(D_EDGE), .C(n11), .Y(n7) );
  NAND2X1 U13 ( .A(n20), .B(state), .Y(n8) );
  NOR2X1 U14 ( .A(D_EDGE), .B(n14), .Y(n9) );
  NAND2X1 U15 ( .A(n5), .B(RCVING), .Y(n10) );
  BUFX2 U16 ( .A(RCVING), .Y(n11) );
  INVX2 U17 ( .A(count[2]), .Y(n13) );
  OAI21X1 U18 ( .A(n22), .B(n13), .C(n21), .Y(n18) );
  XOR2X1 U21 ( .A(n13), .B(n22), .Y(n25) );
  INVX2 U23 ( .A(state), .Y(n14) );
  INVX2 U26 ( .A(n18), .Y(n26) );
  NAND3X1 U27 ( .A(count[3]), .B(n9), .C(n26), .Y(n16) );
  AOI22X1 U28 ( .A(n15), .B(n25), .C(n17), .D(count[3]), .Y(n19) );
  NAND2X1 U29 ( .A(n11), .B(n9), .Y(n24) );
  NOR2X1 U31 ( .A(n19), .B(n24), .Y(nextcount[3]) );
  NOR2X1 U33 ( .A(n22), .B(n24), .Y(nextcount[1]) );
  INVX2 U34 ( .A(count[0]), .Y(n27) );
endmodule


module receiver_block_rewire_1 ( CLK, DM1_RX, DP1_RX, RST, BS_ERROR, CRC_ERROR, 
        EOP_external, OPCODE, RCV_DATA, R_ERROR, W_ENABLE );
  output [1:0] OPCODE;
  output [7:0] RCV_DATA;
  input CLK, DM1_RX, DP1_RX, RST;
  output BS_ERROR, CRC_ERROR, EOP_external, R_ERROR, W_ENABLE;
  wire   n8, SHIFT_ENABLE, BITSTUFF, D_ORIG, D_EDGE, RCVING, n1, n3, n4, n5,
         n6, n7;
  wire   [15:0] RX_CRC;
  wire   [15:0] rx_CHECK_CRC;

  rx_CRC_CALC_1 U_2 ( .CLK(CLK), .RST(RST), .W_ENABLE(n4), .OPCODE({n5, n7}), 
        .RCV_DATA(RCV_DATA), .RX_CRC(RX_CRC) );
  rx_accumulator_1 U_3 ( .CLK(CLK), .RST(RST), .RCV_DATA(RCV_DATA), .W_ENABLE(
        n4), .rx_CHECK_CRC(rx_CHECK_CRC) );
  rx_decode_1 U_1 ( .CLK(CLK), .RST(RST), .DP1_RX(DP1_RX), .SHIFT_ENABLE(n6), 
        .EOP(EOP_external), .D_ORIG(D_ORIG), .BITSTUFF(BITSTUFF), .BS_ERROR(
        BS_ERROR) );
  rx_edgedetect_1 U_0 ( .CLK(CLK), .RST(RST), .DP1_RX(DP1_RX), .D_EDGE(D_EDGE)
         );
  rx_eopdetect_1 U_4 ( .DP1_RX(DP1_RX), .DM1_RX(DM1_RX), .EOP(EOP_external) );
  rx_rcu_1 U_5 ( .CLK(CLK), .RST(RST), .D_EDGE(n1), .EOP(EOP_external), 
        .SHIFT_ENABLE(SHIFT_ENABLE), .BITSTUFF(BITSTUFF), .BS_ERROR(BS_ERROR), 
        .RX_CRC(RX_CRC), .RX_CHECK_CRC(rx_CHECK_CRC), .RCV_DATA({RCV_DATA[7:3], 
        n8, RCV_DATA[1:0]}), .RCVING(RCVING), .W_ENABLE(W_ENABLE), .R_ERROR(
        R_ERROR), .CRC_ERROR(CRC_ERROR), .OPCODE(OPCODE) );
  rx_shift_reg_1 U_6 ( .CLK(CLK), .RST(RST), .SHIFT_ENABLE(SHIFT_ENABLE), 
        .D_ORIG(D_ORIG), .BITSTUFF(BITSTUFF), .RCV_DATA({RCV_DATA[7:3], n8, 
        RCV_DATA[1:0]}) );
  rx_timer_1 U_7 ( .CLK(CLK), .RST(RST), .D_EDGE(D_EDGE), .RCVING(RCVING), 
        .SHIFT_ENABLE(SHIFT_ENABLE) );
  BUFX2 U1 ( .A(D_EDGE), .Y(n1) );
  BUFX2 U2 ( .A(n8), .Y(RCV_DATA[2]) );
  BUFX4 U3 ( .A(SHIFT_ENABLE), .Y(n6) );
  INVX1 U4 ( .A(W_ENABLE), .Y(n3) );
  INVX2 U5 ( .A(n3), .Y(n4) );
  BUFX2 U6 ( .A(OPCODE[1]), .Y(n5) );
  BUFX2 U7 ( .A(OPCODE[0]), .Y(n7) );
endmodule


module tx_CRC_CALC_1 ( CLK, RST, EOP, T_STROBE, PRGA_OPCODE, PRGA_OUT, TX_CRC
 );
  input [1:0] PRGA_OPCODE;
  input [7:0] PRGA_OUT;
  output [15:0] TX_CRC;
  input CLK, RST, EOP, T_STROBE;
  wire   n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n79, n80;

  DFFSR \current_crc_reg[8]  ( .D(n70), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[8]) );
  DFFSR \current_crc_reg[15]  ( .D(n63), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[15]) );
  DFFSR \current_crc_reg[9]  ( .D(n69), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[9]) );
  DFFSR \current_crc_reg[10]  ( .D(n68), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[10]) );
  DFFSR \current_crc_reg[11]  ( .D(n67), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[11]) );
  DFFSR \current_crc_reg[12]  ( .D(n66), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[12]) );
  DFFSR \current_crc_reg[13]  ( .D(n65), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[13]) );
  DFFSR \current_crc_reg[14]  ( .D(n64), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[14]) );
  DFFSR \current_crc_reg[7]  ( .D(n71), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[7]) );
  OAI22X1 U39 ( .A(n25), .B(n20), .C(n38), .D(n19), .Y(n63) );
  XNOR2X1 U40 ( .A(n40), .B(n79), .Y(n38) );
  OAI22X1 U41 ( .A(n37), .B(n20), .C(n19), .D(n36), .Y(n64) );
  OAI22X1 U42 ( .A(n35), .B(n20), .C(n19), .D(n34), .Y(n65) );
  OAI22X1 U43 ( .A(n33), .B(n20), .C(n19), .D(n32), .Y(n66) );
  OAI22X1 U44 ( .A(n31), .B(n20), .C(n19), .D(n30), .Y(n67) );
  OAI22X1 U45 ( .A(n29), .B(n20), .C(n19), .D(n28), .Y(n68) );
  OAI22X1 U46 ( .A(n27), .B(n20), .C(n41), .D(n19), .Y(n69) );
  XNOR2X1 U47 ( .A(TX_CRC[1]), .B(n42), .Y(n41) );
  OAI22X1 U48 ( .A(n24), .B(n20), .C(n43), .D(n19), .Y(n70) );
  XOR2X1 U49 ( .A(n44), .B(n45), .Y(n43) );
  XNOR2X1 U50 ( .A(TX_CRC[0]), .B(n42), .Y(n44) );
  OAI22X1 U51 ( .A(n79), .B(n20), .C(n46), .D(n19), .Y(n71) );
  OAI22X1 U52 ( .A(n20), .B(n36), .C(n47), .D(n19), .Y(n72) );
  XNOR2X1 U53 ( .A(n48), .B(n49), .Y(n47) );
  OAI22X1 U54 ( .A(n20), .B(n34), .C(n50), .D(n19), .Y(n73) );
  OAI22X1 U55 ( .A(n20), .B(n32), .C(n51), .D(n19), .Y(n74) );
  XNOR2X1 U56 ( .A(n52), .B(n53), .Y(n51) );
  OAI22X1 U57 ( .A(n20), .B(n30), .C(n54), .D(n19), .Y(n75) );
  OAI22X1 U58 ( .A(n20), .B(n28), .C(n55), .D(n19), .Y(n76) );
  XOR2X1 U59 ( .A(n56), .B(n57), .Y(n55) );
  OAI22X1 U60 ( .A(n20), .B(n26), .C(n58), .D(n19), .Y(n77) );
  XOR2X1 U61 ( .A(n59), .B(n60), .Y(n58) );
  XOR2X1 U62 ( .A(n42), .B(n46), .Y(n59) );
  OAI22X1 U63 ( .A(n20), .B(n23), .C(n40), .D(n19), .Y(n78) );
  XOR2X1 U64 ( .A(n61), .B(n62), .Y(n40) );
  XOR2X1 U65 ( .A(n57), .B(n42), .Y(n62) );
  XNOR2X1 U66 ( .A(n25), .B(PRGA_OUT[7]), .Y(n42) );
  XNOR2X1 U67 ( .A(n24), .B(PRGA_OUT[0]), .Y(n57) );
  XOR2X1 U68 ( .A(n46), .B(n60), .Y(n61) );
  XOR2X1 U69 ( .A(n54), .B(n50), .Y(n60) );
  XNOR2X1 U70 ( .A(n53), .B(n48), .Y(n50) );
  XOR2X1 U71 ( .A(TX_CRC[12]), .B(PRGA_OUT[4]), .Y(n48) );
  XOR2X1 U72 ( .A(TX_CRC[11]), .B(PRGA_OUT[3]), .Y(n53) );
  XOR2X1 U74 ( .A(TX_CRC[10]), .B(PRGA_OUT[2]), .Y(n52) );
  XNOR2X1 U75 ( .A(TX_CRC[9]), .B(PRGA_OUT[1]), .Y(n56) );
  XNOR2X1 U76 ( .A(n49), .B(n45), .Y(n46) );
  XNOR2X1 U77 ( .A(n37), .B(PRGA_OUT[6]), .Y(n45) );
  XOR2X1 U78 ( .A(TX_CRC[13]), .B(PRGA_OUT[5]), .Y(n49) );
  NAND3X1 U80 ( .A(PRGA_OPCODE[0]), .B(n80), .C(T_STROBE), .Y(n39) );
  DFFSR \current_crc_reg[6]  ( .D(n72), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[6]) );
  DFFSR \current_crc_reg[5]  ( .D(n73), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[5]) );
  DFFSR \current_crc_reg[4]  ( .D(n74), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[4]) );
  DFFSR \current_crc_reg[3]  ( .D(n75), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[3]) );
  DFFSR \current_crc_reg[2]  ( .D(n76), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[2]) );
  DFFSR \current_crc_reg[1]  ( .D(n77), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[1]) );
  DFFSR \current_crc_reg[0]  ( .D(n78), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[0]) );
  INVX4 U5 ( .A(n17), .Y(n20) );
  INVX1 U20 ( .A(EOP), .Y(n22) );
  INVX2 U21 ( .A(n39), .Y(n18) );
  AND2X2 U22 ( .A(n39), .B(n22), .Y(n17) );
  INVX2 U23 ( .A(RST), .Y(n21) );
  XOR2X1 U24 ( .A(n56), .B(n52), .Y(n54) );
  INVX2 U25 ( .A(n18), .Y(n19) );
  INVX2 U26 ( .A(TX_CRC[0]), .Y(n23) );
  INVX2 U27 ( .A(TX_CRC[8]), .Y(n24) );
  INVX2 U28 ( .A(TX_CRC[15]), .Y(n25) );
  INVX2 U29 ( .A(TX_CRC[1]), .Y(n26) );
  INVX2 U30 ( .A(TX_CRC[9]), .Y(n27) );
  INVX2 U31 ( .A(TX_CRC[2]), .Y(n28) );
  INVX2 U32 ( .A(TX_CRC[10]), .Y(n29) );
  INVX2 U33 ( .A(TX_CRC[3]), .Y(n30) );
  INVX2 U34 ( .A(TX_CRC[11]), .Y(n31) );
  INVX2 U35 ( .A(TX_CRC[4]), .Y(n32) );
  INVX2 U36 ( .A(TX_CRC[12]), .Y(n33) );
  INVX2 U37 ( .A(TX_CRC[5]), .Y(n34) );
  INVX2 U38 ( .A(TX_CRC[13]), .Y(n35) );
  INVX2 U73 ( .A(TX_CRC[6]), .Y(n36) );
  INVX2 U79 ( .A(TX_CRC[14]), .Y(n37) );
  INVX2 U81 ( .A(TX_CRC[7]), .Y(n79) );
  INVX2 U82 ( .A(PRGA_OPCODE[1]), .Y(n80) );
endmodule


module tx_encode_1 ( clk, rst, SHIFT_ENABLE_E, d_encode, EOP, t_bitstuff, 
        dp_tx_out, dm_tx_out );
  input clk, rst, SHIFT_ENABLE_E, d_encode, EOP;
  output t_bitstuff, dp_tx_out, dm_tx_out;
  wire   DE_holdout, DE_holdout_BS, DE_holdout_last, DE_holdout_nxt, dm_tx_nxt,
         n9, n12, n13, n14, n15, n18, n19, n20, n26, n27, n32, n37, n39, n40,
         n41, n43, n44, n49, n50, n61, n64, n1, n2, n3, n4, n5, n6, n7, n8,
         n10, n11, n16, n17, n21, n22, n23, n24, n25, n28, n29, n30, n31, n33,
         n34, n35, n36, n38, n42, n45, n46, n47, n48, n51, n52, n53, n63, n65,
         n66, n67;
  wire   [3:0] state;
  wire   [3:0] nextstate;

  DFFSR DE_holdout_reg ( .D(DE_holdout_nxt), .CLK(clk), .R(1'b1), .S(n6), .Q(
        DE_holdout) );
  DFFPOSX1 DE_holdout_last_reg ( .D(n61), .CLK(clk), .Q(DE_holdout_last) );
  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(clk), .R(n6), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n6), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n6), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n6), .S(1'b1), .Q(
        state[2]) );
  DFFSR DE_holdout_BS_reg ( .D(n64), .CLK(clk), .R(n6), .S(1'b1), .Q(
        DE_holdout_BS) );
  DFFSR dp_tx_out_reg ( .D(DE_holdout_nxt), .CLK(clk), .R(1'b1), .S(n6), .Q(
        dp_tx_out) );
  DFFSR dm_tx_out_reg ( .D(dm_tx_nxt), .CLK(clk), .R(n6), .S(1'b1), .Q(
        dm_tx_out) );
  OAI21X1 U9 ( .A(state[1]), .B(n9), .C(n13), .Y(nextstate[1]) );
  OAI21X1 U11 ( .A(n3), .B(n15), .C(n47), .Y(n14) );
  NAND3X1 U12 ( .A(SHIFT_ENABLE_E), .B(n53), .C(n3), .Y(n9) );
  OAI21X1 U14 ( .A(n2), .B(n47), .C(n18), .Y(nextstate[0]) );
  OAI21X1 U15 ( .A(n19), .B(n20), .C(SHIFT_ENABLE_E), .Y(n18) );
  NOR2X1 U18 ( .A(n3), .B(n15), .Y(n19) );
  NAND3X1 U19 ( .A(d_encode), .B(n26), .C(n27), .Y(n15) );
  XNOR2X1 U20 ( .A(n66), .B(n65), .Y(n27) );
  NOR2X1 U22 ( .A(n52), .B(SHIFT_ENABLE_E), .Y(n12) );
  OAI22X1 U23 ( .A(n6), .B(n66), .C(rst), .D(n65), .Y(n61) );
  OAI22X1 U26 ( .A(n5), .B(n67), .C(n65), .D(n32), .Y(n64) );
  NOR2X1 U36 ( .A(EOP), .B(state[3]), .Y(n26) );
  NOR2X1 U37 ( .A(n4), .B(n40), .Y(n37) );
  AOI22X1 U38 ( .A(n3), .B(n41), .C(n48), .D(n2), .Y(n40) );
  XNOR2X1 U40 ( .A(DE_holdout_BS), .B(n44), .Y(n41) );
  XOR2X1 U46 ( .A(DE_holdout), .B(SHIFT_ENABLE_E), .Y(n43) );
  XNOR2X1 U47 ( .A(n49), .B(n65), .Y(n39) );
  NAND2X1 U49 ( .A(SHIFT_ENABLE_E), .B(n63), .Y(n49) );
  NAND2X1 U55 ( .A(n44), .B(n67), .Y(n50) );
  NAND2X1 U57 ( .A(SHIFT_ENABLE_E), .B(d_encode), .Y(n44) );
  INVX1 U3 ( .A(n2), .Y(n3) );
  INVX2 U4 ( .A(state[0]), .Y(n2) );
  AND2X2 U5 ( .A(n27), .B(d_encode), .Y(n1) );
  AND2X2 U6 ( .A(n1), .B(n26), .Y(n53) );
  INVX2 U7 ( .A(n51), .Y(n4) );
  INVX1 U8 ( .A(EOP), .Y(n51) );
  INVX2 U10 ( .A(rst), .Y(n6) );
  NOR2X1 U13 ( .A(n42), .B(n8), .Y(n5) );
  INVX1 U16 ( .A(n5), .Y(n32) );
  NAND2X1 U17 ( .A(state[2]), .B(state[1]), .Y(n7) );
  NOR3X1 U21 ( .A(state[3]), .B(n7), .C(n2), .Y(t_bitstuff) );
  INVX2 U24 ( .A(n7), .Y(n25) );
  NAND3X1 U25 ( .A(n26), .B(n2), .C(n25), .Y(n42) );
  INVX2 U27 ( .A(SHIFT_ENABLE_E), .Y(n8) );
  NAND2X1 U28 ( .A(n63), .B(n25), .Y(n10) );
  OAI21X1 U29 ( .A(n52), .B(n10), .C(n42), .Y(n20) );
  INVX2 U30 ( .A(n42), .Y(n11) );
  AOI21X1 U31 ( .A(n14), .B(state[1]), .C(n11), .Y(n13) );
  INVX2 U32 ( .A(state[2]), .Y(n16) );
  INVX2 U33 ( .A(state[1]), .Y(n33) );
  NAND3X1 U34 ( .A(n2), .B(n16), .C(n33), .Y(n45) );
  NAND2X1 U35 ( .A(n45), .B(state[3]), .Y(n31) );
  INVX2 U39 ( .A(n39), .Y(n17) );
  NOR2X1 U41 ( .A(n52), .B(n17), .Y(n21) );
  MUX2X1 U42 ( .B(n21), .A(n37), .S(n25), .Y(n22) );
  NAND2X1 U43 ( .A(n31), .B(n22), .Y(dm_tx_nxt) );
  OAI21X1 U44 ( .A(n67), .B(n44), .C(n50), .Y(n24) );
  AND2X2 U45 ( .A(n43), .B(n2), .Y(n23) );
  AOI21X1 U48 ( .A(n3), .B(n24), .C(n23), .Y(n28) );
  MUX2X1 U50 ( .B(n39), .A(n28), .S(n25), .Y(n29) );
  OAI21X1 U51 ( .A(state[3]), .B(n29), .C(n51), .Y(n30) );
  NAND2X1 U52 ( .A(n31), .B(n30), .Y(DE_holdout_nxt) );
  NAND2X1 U53 ( .A(n46), .B(state[1]), .Y(n35) );
  AOI21X1 U54 ( .A(n53), .B(n33), .C(n12), .Y(n34) );
  MUX2X1 U56 ( .B(n35), .A(n34), .S(state[2]), .Y(n36) );
  INVX2 U58 ( .A(n36), .Y(n38) );
  NAND2X1 U59 ( .A(n42), .B(n38), .Y(nextstate[2]) );
  AOI21X1 U60 ( .A(state[3]), .B(n45), .C(n51), .Y(nextstate[3]) );
  INVX2 U61 ( .A(n9), .Y(n46) );
  INVX2 U62 ( .A(n12), .Y(n47) );
  INVX2 U63 ( .A(n43), .Y(n48) );
  INVX2 U64 ( .A(n26), .Y(n52) );
  INVX2 U65 ( .A(d_encode), .Y(n63) );
  INVX2 U74 ( .A(DE_holdout), .Y(n65) );
  INVX2 U75 ( .A(DE_holdout_last), .Y(n66) );
  INVX2 U76 ( .A(DE_holdout_BS), .Y(n67) );
endmodule


module tx_shiftreg_1 ( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe, 
        send_data, d_encode );
  input [7:0] send_data;
  input clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe;
  output d_encode;
  wire   n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n11, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69;
  wire   [7:1] present_val;
  wire   [2:0] count;

  DFFSR \count_reg[0]  ( .D(n53), .CLK(clk), .R(1'b1), .S(n17), .Q(count[0])
         );
  DFFSR \count_reg[1]  ( .D(n51), .CLK(clk), .R(1'b1), .S(n17), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n52), .CLK(clk), .R(1'b1), .S(n17), .Q(count[2])
         );
  DFFSR \present_val_reg[7]  ( .D(n44), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[7]) );
  DFFSR \present_val_reg[6]  ( .D(n45), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[6]) );
  DFFSR \present_val_reg[5]  ( .D(n46), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[5]) );
  DFFSR \present_val_reg[4]  ( .D(n47), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[4]) );
  DFFSR \present_val_reg[3]  ( .D(n48), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[3]) );
  DFFSR \present_val_reg[2]  ( .D(n49), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[2]) );
  DFFSR \present_val_reg[1]  ( .D(n50), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[1]) );
  DFFSR \present_val_reg[0]  ( .D(n43), .CLK(clk), .R(n17), .S(1'b1), .Q(
        d_encode) );
  AND2X2 U13 ( .A(n20), .B(n16), .Y(n11) );
  INVX4 U15 ( .A(n11), .Y(n68) );
  INVX4 U16 ( .A(n69), .Y(n65) );
  BUFX4 U17 ( .A(n11), .Y(n13) );
  BUFX2 U18 ( .A(n69), .Y(n14) );
  INVX2 U19 ( .A(rst), .Y(n17) );
  INVX4 U20 ( .A(n15), .Y(n16) );
  INVX2 U21 ( .A(n62), .Y(n15) );
  INVX2 U22 ( .A(t_bitstuff), .Y(n18) );
  NAND2X1 U23 ( .A(SHIFT_ENABLE_R), .B(n18), .Y(n20) );
  NAND2X1 U24 ( .A(count[1]), .B(count[0]), .Y(n64) );
  INVX2 U25 ( .A(n64), .Y(n19) );
  NAND3X1 U26 ( .A(SHIFT_ENABLE_R), .B(count[2]), .C(n19), .Y(n62) );
  NAND2X1 U27 ( .A(d_encode), .B(n13), .Y(n24) );
  NAND2X1 U28 ( .A(n68), .B(n16), .Y(n69) );
  NAND2X1 U29 ( .A(present_val[1]), .B(n65), .Y(n23) );
  INVX2 U30 ( .A(send_data[0]), .Y(n21) );
  OR2X2 U31 ( .A(n16), .B(n21), .Y(n22) );
  NAND3X1 U32 ( .A(n22), .B(n23), .C(n24), .Y(n43) );
  NAND2X1 U33 ( .A(present_val[1]), .B(n13), .Y(n28) );
  NAND2X1 U34 ( .A(present_val[2]), .B(n65), .Y(n27) );
  INVX2 U35 ( .A(send_data[1]), .Y(n25) );
  OR2X2 U36 ( .A(n16), .B(n25), .Y(n26) );
  NAND3X1 U37 ( .A(n28), .B(n27), .C(n26), .Y(n50) );
  NAND2X1 U38 ( .A(present_val[2]), .B(n13), .Y(n32) );
  NAND2X1 U39 ( .A(present_val[3]), .B(n65), .Y(n31) );
  INVX2 U40 ( .A(send_data[2]), .Y(n29) );
  OR2X2 U41 ( .A(n16), .B(n29), .Y(n30) );
  NAND3X1 U42 ( .A(n32), .B(n31), .C(n30), .Y(n49) );
  NAND2X1 U43 ( .A(present_val[3]), .B(n13), .Y(n36) );
  NAND2X1 U44 ( .A(present_val[4]), .B(n65), .Y(n35) );
  INVX2 U45 ( .A(send_data[3]), .Y(n33) );
  OR2X2 U46 ( .A(n16), .B(n33), .Y(n34) );
  NAND3X1 U47 ( .A(n36), .B(n35), .C(n34), .Y(n48) );
  NAND2X1 U48 ( .A(present_val[4]), .B(n13), .Y(n40) );
  NAND2X1 U49 ( .A(present_val[5]), .B(n65), .Y(n39) );
  INVX2 U50 ( .A(send_data[4]), .Y(n37) );
  OR2X2 U51 ( .A(n16), .B(n37), .Y(n38) );
  NAND3X1 U52 ( .A(n40), .B(n39), .C(n38), .Y(n47) );
  NAND2X1 U53 ( .A(present_val[5]), .B(n13), .Y(n55) );
  NAND2X1 U54 ( .A(present_val[6]), .B(n65), .Y(n54) );
  INVX2 U55 ( .A(send_data[5]), .Y(n41) );
  OR2X2 U56 ( .A(n16), .B(n41), .Y(n42) );
  NAND3X1 U57 ( .A(n55), .B(n54), .C(n42), .Y(n46) );
  NAND2X1 U58 ( .A(present_val[6]), .B(n13), .Y(n59) );
  NAND2X1 U59 ( .A(present_val[7]), .B(n65), .Y(n58) );
  INVX2 U60 ( .A(send_data[6]), .Y(n56) );
  OR2X2 U61 ( .A(n16), .B(n56), .Y(n57) );
  NAND3X1 U62 ( .A(n59), .B(n58), .C(n57), .Y(n45) );
  INVX2 U63 ( .A(present_val[7]), .Y(n61) );
  INVX2 U64 ( .A(send_data[7]), .Y(n60) );
  OAI22X1 U65 ( .A(n68), .B(n61), .C(n16), .D(n60), .Y(n44) );
  NAND2X1 U66 ( .A(count[2]), .B(n16), .Y(n63) );
  OAI21X1 U67 ( .A(n64), .B(n14), .C(n63), .Y(n52) );
  NAND2X1 U68 ( .A(n65), .B(count[0]), .Y(n67) );
  AND2X2 U69 ( .A(count[0]), .B(n68), .Y(n66) );
  MUX2X1 U70 ( .B(n67), .A(n66), .S(count[1]), .Y(n51) );
  MUX2X1 U71 ( .B(n14), .A(n68), .S(count[0]), .Y(n53) );
endmodule


module tx_tcu_1_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module tx_tcu_1 ( clk, rst, p_ready, t_bitstuff, PRGA_OUT, prga_opcode, t_crc, 
        sending, EOP, next_byte, send_data, t_strobe );
  input [7:0] PRGA_OUT;
  input [1:0] prga_opcode;
  input [15:0] t_crc;
  output [7:0] send_data;
  input clk, rst, p_ready, t_bitstuff;
  output sending, EOP, next_byte, t_strobe;
  wire   N59, N60, N61, N62, N63, N64, N65, N188, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n194, n195, n196, n197, n198, n199, n200, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256;
  wire   [2:0] state;
  wire   [6:0] count;
  wire   [2:0] nextstate;
  wire   [7:0] flop_data;
  wire   [7:0] current_send_data;

  DFFSR \count_reg[0]  ( .D(n200), .CLK(clk), .R(n25), .S(1'b1), .Q(count[0])
         );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n25), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n25), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n25), .S(1'b1), .Q(
        state[2]) );
  DFFSR \count_reg[6]  ( .D(n199), .CLK(clk), .R(n25), .S(1'b1), .Q(N188) );
  DFFSR \count_reg[1]  ( .D(n194), .CLK(clk), .R(n25), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[5]  ( .D(n198), .CLK(clk), .R(n25), .S(1'b1), .Q(count[5])
         );
  DFFSR \count_reg[2]  ( .D(n195), .CLK(clk), .R(n25), .S(1'b1), .Q(count[2])
         );
  DFFSR \count_reg[3]  ( .D(n196), .CLK(clk), .R(n25), .S(1'b1), .Q(count[3])
         );
  DFFSR \count_reg[4]  ( .D(n197), .CLK(clk), .R(n25), .S(1'b1), .Q(count[4])
         );
  DFFPOSX1 \flop_data_reg[7]  ( .D(n249), .CLK(clk), .Q(flop_data[7]) );
  DFFPOSX1 \current_send_data_reg[7]  ( .D(n173), .CLK(clk), .Q(
        current_send_data[7]) );
  DFFPOSX1 \flop_data_reg[6]  ( .D(n250), .CLK(clk), .Q(flop_data[6]) );
  DFFPOSX1 \current_send_data_reg[6]  ( .D(n172), .CLK(clk), .Q(
        current_send_data[6]) );
  DFFPOSX1 \flop_data_reg[5]  ( .D(n251), .CLK(clk), .Q(flop_data[5]) );
  DFFPOSX1 \current_send_data_reg[5]  ( .D(n171), .CLK(clk), .Q(
        current_send_data[5]) );
  DFFPOSX1 \flop_data_reg[4]  ( .D(n252), .CLK(clk), .Q(flop_data[4]) );
  DFFPOSX1 \current_send_data_reg[4]  ( .D(n170), .CLK(clk), .Q(
        current_send_data[4]) );
  DFFPOSX1 \flop_data_reg[3]  ( .D(n253), .CLK(clk), .Q(flop_data[3]) );
  DFFPOSX1 \current_send_data_reg[3]  ( .D(n169), .CLK(clk), .Q(
        current_send_data[3]) );
  DFFPOSX1 \flop_data_reg[2]  ( .D(n254), .CLK(clk), .Q(flop_data[2]) );
  DFFPOSX1 \current_send_data_reg[2]  ( .D(n168), .CLK(clk), .Q(
        current_send_data[2]) );
  DFFPOSX1 \flop_data_reg[1]  ( .D(n255), .CLK(clk), .Q(flop_data[1]) );
  DFFPOSX1 \current_send_data_reg[1]  ( .D(n167), .CLK(clk), .Q(
        current_send_data[1]) );
  DFFPOSX1 \flop_data_reg[0]  ( .D(n256), .CLK(clk), .Q(flop_data[0]) );
  DFFPOSX1 \current_send_data_reg[0]  ( .D(n166), .CLK(clk), .Q(
        current_send_data[0]) );
  DFFPOSX1 \send_data_reg[7]  ( .D(n165), .CLK(clk), .Q(send_data[7]) );
  DFFPOSX1 \send_data_reg[6]  ( .D(n164), .CLK(clk), .Q(send_data[6]) );
  DFFPOSX1 \send_data_reg[5]  ( .D(n163), .CLK(clk), .Q(send_data[5]) );
  DFFPOSX1 \send_data_reg[4]  ( .D(n162), .CLK(clk), .Q(send_data[4]) );
  DFFPOSX1 \send_data_reg[3]  ( .D(n161), .CLK(clk), .Q(send_data[3]) );
  DFFPOSX1 \send_data_reg[2]  ( .D(n160), .CLK(clk), .Q(send_data[2]) );
  DFFPOSX1 \send_data_reg[1]  ( .D(n159), .CLK(clk), .Q(send_data[1]) );
  DFFPOSX1 \send_data_reg[0]  ( .D(n158), .CLK(clk), .Q(send_data[0]) );
  tx_tcu_1_DW01_inc_0 r80 ( .A({n23, count[5], n1, n2, n5, count[1:0]}), .SUM(
        {N65, N64, N63, N62, N61, N60, N59}) );
  INVX2 U3 ( .A(count[2]), .Y(n186) );
  INVX2 U4 ( .A(n156), .Y(n10) );
  INVX2 U5 ( .A(count[0]), .Y(n150) );
  INVX2 U6 ( .A(n186), .Y(n5) );
  BUFX4 U7 ( .A(count[4]), .Y(n1) );
  BUFX4 U8 ( .A(count[3]), .Y(n2) );
  INVX2 U9 ( .A(n187), .Y(n3) );
  INVX2 U10 ( .A(n118), .Y(n4) );
  OR2X2 U11 ( .A(n104), .B(n13), .Y(n6) );
  INVX1 U12 ( .A(n134), .Y(n84) );
  INVX1 U13 ( .A(n11), .Y(n130) );
  NAND2X1 U14 ( .A(n147), .B(n146), .Y(n7) );
  NAND2X1 U15 ( .A(n8), .B(n247), .Y(n245) );
  INVX2 U16 ( .A(n7), .Y(n8) );
  INVX1 U17 ( .A(n120), .Y(n131) );
  OR2X1 U18 ( .A(n9), .B(n104), .Y(n114) );
  NAND2X1 U19 ( .A(n113), .B(n105), .Y(n9) );
  AND2X2 U20 ( .A(n5), .B(n20), .Y(n21) );
  INVX4 U21 ( .A(n24), .Y(n30) );
  INVX2 U22 ( .A(n11), .Y(n155) );
  OR2X2 U23 ( .A(n11), .B(n10), .Y(n133) );
  OR2X2 U24 ( .A(n188), .B(n189), .Y(n11) );
  AND2X2 U25 ( .A(n125), .B(n88), .Y(n12) );
  INVX4 U26 ( .A(n12), .Y(n140) );
  INVX1 U27 ( .A(n105), .Y(n13) );
  INVX1 U28 ( .A(n133), .Y(n119) );
  INVX2 U29 ( .A(state[1]), .Y(n14) );
  INVX1 U30 ( .A(n14), .Y(n15) );
  INVX4 U31 ( .A(n14), .Y(n16) );
  AND2X2 U32 ( .A(count[1]), .B(n18), .Y(n20) );
  AND2X1 U33 ( .A(n154), .B(n118), .Y(n17) );
  OR2X1 U34 ( .A(n30), .B(n29), .Y(n22) );
  INVX2 U35 ( .A(rst), .Y(n25) );
  NOR2X1 U36 ( .A(t_bitstuff), .B(n150), .Y(n18) );
  AND2X2 U37 ( .A(state[2]), .B(n16), .Y(n19) );
  BUFX4 U38 ( .A(N188), .Y(n23) );
  BUFX4 U39 ( .A(state[0]), .Y(n24) );
  XOR2X1 U40 ( .A(n18), .B(n3), .Y(n109) );
  XOR2X1 U41 ( .A(n21), .B(n2), .Y(n93) );
  XOR2X1 U42 ( .A(n20), .B(n5), .Y(n98) );
  OR2X2 U43 ( .A(n22), .B(n218), .Y(n27) );
  INVX1 U44 ( .A(n87), .Y(n118) );
  INVX1 U45 ( .A(n15), .Y(n26) );
  INVX2 U46 ( .A(n23), .Y(n145) );
  INVX2 U47 ( .A(state[2]), .Y(n58) );
  NAND3X1 U48 ( .A(n24), .B(n58), .C(n26), .Y(n82) );
  NAND3X1 U49 ( .A(n16), .B(n58), .C(n30), .Y(n87) );
  NAND2X1 U50 ( .A(n82), .B(n87), .Y(n63) );
  NAND2X1 U51 ( .A(n63), .B(n25), .Y(n50) );
  NAND2X1 U52 ( .A(state[2]), .B(n26), .Y(n29) );
  OAI21X1 U53 ( .A(n184), .B(n50), .C(n27), .Y(n216) );
  NAND2X1 U54 ( .A(n19), .B(n30), .Y(n59) );
  INVX2 U55 ( .A(n59), .Y(n28) );
  NAND2X1 U56 ( .A(n28), .B(n25), .Y(n33) );
  INVX2 U57 ( .A(n29), .Y(n62) );
  NAND2X1 U58 ( .A(n62), .B(n30), .Y(n120) );
  NAND2X1 U59 ( .A(n131), .B(n25), .Y(n32) );
  INVX2 U60 ( .A(t_crc[15]), .Y(n31) );
  OAI22X1 U61 ( .A(n157), .B(n33), .C(n32), .D(n31), .Y(n217) );
  INVX2 U62 ( .A(n32), .Y(n47) );
  INVX2 U63 ( .A(n33), .Y(n46) );
  AOI22X1 U64 ( .A(t_crc[14]), .B(n47), .C(PRGA_OUT[6]), .D(n46), .Y(n221) );
  INVX2 U65 ( .A(flop_data[6]), .Y(n80) );
  NAND3X1 U66 ( .A(n241), .B(n24), .C(n62), .Y(n49) );
  INVX2 U67 ( .A(t_crc[6]), .Y(n34) );
  OAI22X1 U68 ( .A(n50), .B(n80), .C(n49), .D(n34), .Y(n35) );
  INVX2 U69 ( .A(n35), .Y(n222) );
  AOI22X1 U70 ( .A(t_crc[13]), .B(n47), .C(PRGA_OUT[5]), .D(n46), .Y(n224) );
  INVX2 U71 ( .A(flop_data[5]), .Y(n78) );
  INVX2 U72 ( .A(t_crc[5]), .Y(n36) );
  OAI22X1 U73 ( .A(n50), .B(n78), .C(n49), .D(n36), .Y(n37) );
  INVX2 U74 ( .A(n37), .Y(n225) );
  AOI22X1 U75 ( .A(t_crc[12]), .B(n47), .C(PRGA_OUT[4]), .D(n46), .Y(n227) );
  INVX2 U76 ( .A(flop_data[4]), .Y(n76) );
  INVX2 U77 ( .A(t_crc[4]), .Y(n38) );
  OAI22X1 U78 ( .A(n50), .B(n76), .C(n49), .D(n38), .Y(n39) );
  INVX2 U79 ( .A(n39), .Y(n228) );
  AOI22X1 U80 ( .A(t_crc[11]), .B(n47), .C(PRGA_OUT[3]), .D(n46), .Y(n230) );
  INVX2 U81 ( .A(flop_data[3]), .Y(n74) );
  INVX2 U82 ( .A(t_crc[3]), .Y(n40) );
  OAI22X1 U83 ( .A(n50), .B(n74), .C(n49), .D(n40), .Y(n41) );
  INVX2 U84 ( .A(n41), .Y(n231) );
  AOI22X1 U85 ( .A(t_crc[10]), .B(n47), .C(PRGA_OUT[2]), .D(n46), .Y(n233) );
  INVX2 U86 ( .A(flop_data[2]), .Y(n72) );
  INVX2 U87 ( .A(t_crc[2]), .Y(n42) );
  OAI22X1 U88 ( .A(n50), .B(n72), .C(n49), .D(n42), .Y(n43) );
  INVX2 U89 ( .A(n43), .Y(n234) );
  AOI22X1 U90 ( .A(t_crc[9]), .B(n47), .C(PRGA_OUT[1]), .D(n46), .Y(n236) );
  INVX2 U91 ( .A(flop_data[1]), .Y(n70) );
  INVX2 U92 ( .A(t_crc[1]), .Y(n44) );
  OAI22X1 U93 ( .A(n50), .B(n70), .C(n49), .D(n44), .Y(n45) );
  INVX2 U94 ( .A(n45), .Y(n237) );
  AOI22X1 U95 ( .A(t_crc[8]), .B(n47), .C(PRGA_OUT[0]), .D(n46), .Y(n239) );
  INVX2 U96 ( .A(flop_data[0]), .Y(n68) );
  INVX2 U97 ( .A(t_crc[0]), .Y(n48) );
  OAI22X1 U98 ( .A(n50), .B(n68), .C(n49), .D(n48), .Y(n51) );
  INVX2 U99 ( .A(n51), .Y(n240) );
  INVX2 U100 ( .A(count[4]), .Y(n147) );
  INVX2 U101 ( .A(count[5]), .Y(n146) );
  INVX2 U102 ( .A(n82), .Y(n132) );
  NAND2X1 U103 ( .A(n149), .B(n132), .Y(n52) );
  NOR2X1 U104 ( .A(n148), .B(n52), .Y(t_strobe) );
  NOR3X1 U105 ( .A(n16), .B(n24), .C(state[2]), .Y(n124) );
  INVX2 U106 ( .A(p_ready), .Y(n53) );
  NAND2X1 U107 ( .A(n124), .B(n53), .Y(n64) );
  OAI21X1 U108 ( .A(n156), .B(n4), .C(n64), .Y(n54) );
  AOI21X1 U109 ( .A(n19), .B(n24), .C(n54), .Y(n55) );
  INVX2 U110 ( .A(n55), .Y(next_byte) );
  NAND2X1 U111 ( .A(n243), .B(n23), .Y(n57) );
  INVX2 U112 ( .A(n244), .Y(n56) );
  NAND2X1 U113 ( .A(n62), .B(n56), .Y(n134) );
  OAI22X1 U114 ( .A(n57), .B(n134), .C(n154), .D(n4), .Y(EOP) );
  NAND2X1 U115 ( .A(n62), .B(n145), .Y(n61) );
  NAND3X1 U116 ( .A(n24), .B(n16), .C(n58), .Y(n86) );
  NAND2X1 U117 ( .A(n59), .B(n86), .Y(n135) );
  NOR2X1 U118 ( .A(n135), .B(n63), .Y(n60) );
  NAND3X1 U119 ( .A(n120), .B(n61), .C(n60), .Y(sending) );
  INVX2 U120 ( .A(PRGA_OUT[0]), .Y(n67) );
  NOR3X1 U121 ( .A(n63), .B(n19), .C(n62), .Y(n66) );
  AND2X2 U122 ( .A(n64), .B(n25), .Y(n65) );
  AND2X2 U123 ( .A(n66), .B(n65), .Y(n81) );
  MUX2X1 U124 ( .B(n68), .A(n67), .S(n81), .Y(n256) );
  INVX2 U125 ( .A(PRGA_OUT[1]), .Y(n69) );
  MUX2X1 U126 ( .B(n70), .A(n69), .S(n81), .Y(n255) );
  INVX2 U127 ( .A(PRGA_OUT[2]), .Y(n71) );
  MUX2X1 U128 ( .B(n72), .A(n71), .S(n81), .Y(n254) );
  INVX2 U129 ( .A(PRGA_OUT[3]), .Y(n73) );
  MUX2X1 U130 ( .B(n74), .A(n73), .S(n81), .Y(n253) );
  INVX2 U131 ( .A(PRGA_OUT[4]), .Y(n75) );
  MUX2X1 U132 ( .B(n76), .A(n75), .S(n81), .Y(n252) );
  INVX2 U133 ( .A(PRGA_OUT[5]), .Y(n77) );
  MUX2X1 U134 ( .B(n78), .A(n77), .S(n81), .Y(n251) );
  INVX2 U135 ( .A(PRGA_OUT[6]), .Y(n79) );
  MUX2X1 U136 ( .B(n80), .A(n79), .S(n81), .Y(n250) );
  MUX2X1 U137 ( .B(n184), .A(n157), .S(n81), .Y(n249) );
  OAI21X1 U138 ( .A(n155), .B(n120), .C(n82), .Y(n83) );
  NAND2X1 U139 ( .A(t_bitstuff), .B(n132), .Y(n94) );
  OAI21X1 U140 ( .A(n84), .B(n83), .C(n94), .Y(n85) );
  INVX2 U141 ( .A(n85), .Y(n139) );
  NAND2X1 U142 ( .A(N63), .B(n139), .Y(n92) );
  NAND2X1 U143 ( .A(n2), .B(n21), .Y(n102) );
  OR2X2 U144 ( .A(n155), .B(n86), .Y(n125) );
  NAND2X1 U145 ( .A(n118), .B(n133), .Y(n88) );
  NOR2X1 U146 ( .A(n102), .B(n12), .Y(n90) );
  NAND2X1 U147 ( .A(n102), .B(n140), .Y(n89) );
  NAND2X1 U148 ( .A(n89), .B(n94), .Y(n104) );
  MUX2X1 U149 ( .B(n90), .A(n104), .S(n1), .Y(n91) );
  NAND2X1 U150 ( .A(n92), .B(n91), .Y(n197) );
  NAND2X1 U151 ( .A(N62), .B(n139), .Y(n97) );
  NAND2X1 U152 ( .A(n93), .B(n140), .Y(n96) );
  INVX2 U153 ( .A(n94), .Y(n142) );
  NAND2X1 U154 ( .A(n142), .B(n2), .Y(n95) );
  NAND3X1 U155 ( .A(n97), .B(n96), .C(n95), .Y(n196) );
  NAND2X1 U156 ( .A(N61), .B(n139), .Y(n101) );
  NAND2X1 U157 ( .A(n98), .B(n140), .Y(n100) );
  NAND2X1 U158 ( .A(n142), .B(n5), .Y(n99) );
  NAND3X1 U159 ( .A(n101), .B(n100), .C(n99), .Y(n195) );
  NAND2X1 U160 ( .A(N64), .B(n139), .Y(n108) );
  INVX2 U161 ( .A(n102), .Y(n103) );
  NAND3X1 U162 ( .A(n103), .B(n1), .C(n140), .Y(n112) );
  INVX2 U163 ( .A(n112), .Y(n106) );
  NAND2X1 U164 ( .A(n140), .B(n147), .Y(n105) );
  MUX2X1 U165 ( .B(n106), .A(n6), .S(count[5]), .Y(n107) );
  NAND2X1 U166 ( .A(n108), .B(n107), .Y(n198) );
  AOI22X1 U167 ( .A(n109), .B(n140), .C(N60), .D(n139), .Y(n111) );
  NAND2X1 U168 ( .A(n142), .B(n3), .Y(n110) );
  NAND2X1 U169 ( .A(n111), .B(n110), .Y(n194) );
  NAND2X1 U170 ( .A(N65), .B(n139), .Y(n117) );
  NOR2X1 U171 ( .A(n146), .B(n112), .Y(n115) );
  NAND2X1 U172 ( .A(n140), .B(n146), .Y(n113) );
  MUX2X1 U173 ( .B(n115), .A(n114), .S(n23), .Y(n116) );
  NAND2X1 U174 ( .A(n117), .B(n116), .Y(n199) );
  NAND2X1 U175 ( .A(n151), .B(p_ready), .Y(n123) );
  NAND2X1 U176 ( .A(n119), .B(n17), .Y(n122) );
  AND2X2 U177 ( .A(n120), .B(n134), .Y(n121) );
  NAND3X1 U178 ( .A(n123), .B(n122), .C(n121), .Y(nextstate[2]) );
  NAND2X1 U179 ( .A(n124), .B(p_ready), .Y(n129) );
  NAND2X1 U180 ( .A(n17), .B(n133), .Y(n128) );
  INVX2 U181 ( .A(n125), .Y(n126) );
  AOI21X1 U182 ( .A(n152), .B(n132), .C(n126), .Y(n127) );
  NAND3X1 U183 ( .A(n129), .B(n128), .C(n127), .Y(nextstate[1]) );
  AOI22X1 U184 ( .A(n153), .B(n132), .C(n131), .D(n130), .Y(n138) );
  NAND3X1 U185 ( .A(n17), .B(n133), .C(p_ready), .Y(n137) );
  NOR2X1 U186 ( .A(n135), .B(n84), .Y(n136) );
  NAND3X1 U187 ( .A(n138), .B(n137), .C(n136), .Y(nextstate[0]) );
  XOR2X1 U188 ( .A(n150), .B(t_bitstuff), .Y(n141) );
  AOI22X1 U189 ( .A(n141), .B(n140), .C(N59), .D(n139), .Y(n144) );
  NAND2X1 U190 ( .A(n142), .B(count[0]), .Y(n143) );
  NAND2X1 U191 ( .A(n144), .B(n143), .Y(n200) );
  NAND2X1 U192 ( .A(n145), .B(n150), .Y(n148) );
  NOR2X1 U203 ( .A(n16), .B(n24), .Y(n151) );
  INVX1 U204 ( .A(n153), .Y(n152) );
  NAND3X1 U205 ( .A(n149), .B(n145), .C(count[0]), .Y(n153) );
  AND2X1 U206 ( .A(prga_opcode[1]), .B(prga_opcode[0]), .Y(n156) );
  NAND3X1 U207 ( .A(n1), .B(count[1]), .C(count[5]), .Y(n189) );
  NAND3X1 U208 ( .A(count[0]), .B(n2), .C(n190), .Y(n188) );
  NOR2X1 U209 ( .A(n23), .B(n186), .Y(n190) );
  INVX1 U210 ( .A(count[1]), .Y(n187) );
  OAI21X1 U211 ( .A(n191), .B(n192), .C(n193), .Y(n173) );
  INVX1 U212 ( .A(current_send_data[7]), .Y(n192) );
  OAI21X1 U213 ( .A(n191), .B(n201), .C(n202), .Y(n172) );
  INVX1 U214 ( .A(current_send_data[6]), .Y(n201) );
  OAI21X1 U215 ( .A(n191), .B(n203), .C(n204), .Y(n171) );
  INVX1 U216 ( .A(current_send_data[5]), .Y(n203) );
  OAI21X1 U217 ( .A(n191), .B(n205), .C(n206), .Y(n170) );
  INVX1 U218 ( .A(current_send_data[4]), .Y(n205) );
  OAI21X1 U219 ( .A(n191), .B(n207), .C(n208), .Y(n169) );
  INVX1 U220 ( .A(current_send_data[3]), .Y(n207) );
  OAI21X1 U221 ( .A(n191), .B(n209), .C(n210), .Y(n168) );
  INVX1 U222 ( .A(current_send_data[2]), .Y(n209) );
  OAI21X1 U223 ( .A(n191), .B(n211), .C(n212), .Y(n167) );
  INVX1 U224 ( .A(current_send_data[1]), .Y(n211) );
  OAI21X1 U225 ( .A(n191), .B(n213), .C(n214), .Y(n166) );
  INVX1 U226 ( .A(current_send_data[0]), .Y(n213) );
  AOI21X1 U227 ( .A(n24), .B(n16), .C(rst), .Y(n191) );
  NAND2X1 U228 ( .A(n215), .B(n193), .Y(n165) );
  NOR2X1 U229 ( .A(n216), .B(n217), .Y(n193) );
  INVX1 U230 ( .A(PRGA_OUT[7]), .Y(n157) );
  OAI21X1 U231 ( .A(n23), .B(t_crc[7]), .C(n25), .Y(n218) );
  INVX1 U232 ( .A(flop_data[7]), .Y(n184) );
  AOI22X1 U233 ( .A(n219), .B(current_send_data[7]), .C(send_data[7]), .D(rst), 
        .Y(n215) );
  NAND2X1 U234 ( .A(n220), .B(n202), .Y(n164) );
  AND2X1 U235 ( .A(n221), .B(n222), .Y(n202) );
  AOI22X1 U236 ( .A(n219), .B(current_send_data[6]), .C(send_data[6]), .D(rst), 
        .Y(n220) );
  NAND2X1 U237 ( .A(n223), .B(n204), .Y(n163) );
  AND2X1 U238 ( .A(n224), .B(n225), .Y(n204) );
  AOI22X1 U239 ( .A(n219), .B(current_send_data[5]), .C(send_data[5]), .D(rst), 
        .Y(n223) );
  NAND2X1 U240 ( .A(n226), .B(n206), .Y(n162) );
  AND2X1 U241 ( .A(n227), .B(n228), .Y(n206) );
  AOI22X1 U242 ( .A(n219), .B(current_send_data[4]), .C(send_data[4]), .D(rst), 
        .Y(n226) );
  NAND2X1 U243 ( .A(n229), .B(n208), .Y(n161) );
  AND2X1 U244 ( .A(n230), .B(n231), .Y(n208) );
  AOI22X1 U245 ( .A(n219), .B(current_send_data[3]), .C(send_data[3]), .D(rst), 
        .Y(n229) );
  NAND2X1 U246 ( .A(n232), .B(n210), .Y(n160) );
  AND2X1 U247 ( .A(n233), .B(n234), .Y(n210) );
  AOI22X1 U248 ( .A(n219), .B(current_send_data[2]), .C(send_data[2]), .D(rst), 
        .Y(n232) );
  NAND2X1 U249 ( .A(n235), .B(n212), .Y(n159) );
  AND2X1 U250 ( .A(n236), .B(n237), .Y(n212) );
  AOI22X1 U251 ( .A(n219), .B(current_send_data[1]), .C(send_data[1]), .D(rst), 
        .Y(n235) );
  NAND2X1 U252 ( .A(n238), .B(n214), .Y(n158) );
  AND2X1 U253 ( .A(n239), .B(n240), .Y(n214) );
  NOR2X1 U254 ( .A(rst), .B(n23), .Y(n241) );
  AOI22X1 U255 ( .A(n219), .B(current_send_data[0]), .C(send_data[0]), .D(rst), 
        .Y(n238) );
  INVX1 U256 ( .A(n242), .Y(n219) );
  NAND3X1 U257 ( .A(n24), .B(n25), .C(n16), .Y(n242) );
  OAI21X1 U258 ( .A(n245), .B(n246), .C(n24), .Y(n244) );
  NAND3X1 U259 ( .A(n5), .B(n23), .C(n2), .Y(n246) );
  NOR2X1 U260 ( .A(count[1]), .B(count[0]), .Y(n247) );
  NAND3X1 U261 ( .A(n149), .B(n150), .C(n23), .Y(n154) );
  NOR2X1 U262 ( .A(n243), .B(count[1]), .Y(n149) );
  NAND3X1 U263 ( .A(n186), .B(n185), .C(n248), .Y(n243) );
  NOR2X1 U264 ( .A(count[5]), .B(n1), .Y(n248) );
  INVX1 U265 ( .A(count[3]), .Y(n185) );
endmodule


module tx_timer_1 ( CLK, RST, SENDING, SHIFT_ENABLE_R, SHIFT_ENABLE_E );
  input CLK, RST, SENDING;
  output SHIFT_ENABLE_R, SHIFT_ENABLE_E;
  wire   state, nxt_SHIFT_ENABLE_E, n12, n13, n14, n15, n16, n17, n18, n6, n8,
         n9, n10, n11, n19, n20, n21, n22;
  wire   [3:0] count;
  wire   [3:0] nextcount;
  assign SHIFT_ENABLE_R = nxt_SHIFT_ENABLE_E;

  DFFSR state_reg ( .D(n8), .CLK(CLK), .R(n9), .S(1'b1), .Q(state) );
  DFFSR \count_reg[0]  ( .D(nextcount[0]), .CLK(CLK), .R(n9), .S(1'b1), .Q(
        count[0]) );
  DFFSR \count_reg[2]  ( .D(nextcount[2]), .CLK(CLK), .R(n9), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[1]  ( .D(nextcount[1]), .CLK(CLK), .R(n9), .S(1'b1), .Q(
        count[1]) );
  DFFSR \count_reg[3]  ( .D(nextcount[3]), .CLK(CLK), .R(n9), .S(1'b1), .Q(
        count[3]) );
  DFFSR SHIFT_ENABLE_E_reg ( .D(nxt_SHIFT_ENABLE_E), .CLK(CLK), .R(n9), .S(
        1'b1), .Q(SHIFT_ENABLE_E) );
  NOR2X1 U14 ( .A(n12), .B(n13), .Y(nextcount[3]) );
  XNOR2X1 U15 ( .A(count[3]), .B(n14), .Y(n12) );
  NOR2X1 U16 ( .A(n15), .B(n21), .Y(n14) );
  AOI21X1 U17 ( .A(n16), .B(state), .C(n22), .Y(nextcount[2]) );
  XNOR2X1 U18 ( .A(n15), .B(n21), .Y(n16) );
  NAND2X1 U19 ( .A(count[1]), .B(count[0]), .Y(n15) );
  NOR2X1 U20 ( .A(n17), .B(n13), .Y(nextcount[1]) );
  NAND3X1 U21 ( .A(n8), .B(n18), .C(state), .Y(n13) );
  XNOR2X1 U22 ( .A(count[0]), .B(count[1]), .Y(n17) );
  OAI21X1 U23 ( .A(count[0]), .B(n22), .C(state), .Y(nextcount[0]) );
  AND2X1 U8 ( .A(n20), .B(n19), .Y(n6) );
  AND2X2 U10 ( .A(SENDING), .B(n6), .Y(nxt_SHIFT_ENABLE_E) );
  INVX2 U11 ( .A(n22), .Y(n8) );
  INVX1 U12 ( .A(SENDING), .Y(n22) );
  INVX2 U13 ( .A(RST), .Y(n9) );
  NOR2X1 U24 ( .A(count[0]), .B(count[2]), .Y(n11) );
  INVX2 U25 ( .A(count[1]), .Y(n10) );
  NAND2X1 U26 ( .A(n11), .B(n10), .Y(n18) );
  INVX2 U27 ( .A(n18), .Y(n20) );
  AND2X2 U28 ( .A(count[3]), .B(state), .Y(n19) );
  INVX2 U29 ( .A(count[2]), .Y(n21) );
endmodule


module transmitter_block_1 ( PRGA_OUT, clk, p_ready, prga_opcode, rst, SENDING, 
        dm_tx_out, dp_tx_out, NEXT_BYTE );
  input [7:0] PRGA_OUT;
  input [1:0] prga_opcode;
  input clk, p_ready, rst;
  output SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE;
  wire   t_strobe, EOP, SHIFT_ENABLE_E, d_encode, t_bitstuff, SHIFT_ENABLE_R;
  wire   [15:0] TX_CRC;
  wire   [7:0] send_data;

  tx_CRC_CALC_1 U_1 ( .CLK(clk), .RST(rst), .EOP(EOP), .T_STROBE(t_strobe), 
        .PRGA_OPCODE(prga_opcode), .PRGA_OUT(PRGA_OUT), .TX_CRC(TX_CRC) );
  tx_encode_1 U_0 ( .clk(clk), .rst(rst), .SHIFT_ENABLE_E(SHIFT_ENABLE_E), 
        .d_encode(d_encode), .EOP(EOP), .t_bitstuff(t_bitstuff), .dp_tx_out(
        dp_tx_out), .dm_tx_out(dm_tx_out) );
  tx_shiftreg_1 U_2 ( .clk(clk), .rst(rst), .SHIFT_ENABLE_R(SHIFT_ENABLE_R), 
        .t_bitstuff(t_bitstuff), .t_strobe(t_strobe), .send_data(send_data), 
        .d_encode(d_encode) );
  tx_tcu_1 U_3 ( .clk(clk), .rst(rst), .p_ready(p_ready), .t_bitstuff(
        t_bitstuff), .PRGA_OUT(PRGA_OUT), .prga_opcode(prga_opcode), .t_crc(
        TX_CRC), .sending(SENDING), .EOP(EOP), .next_byte(NEXT_BYTE), 
        .send_data(send_data), .t_strobe(t_strobe) );
  tx_timer_1 U_4 ( .CLK(clk), .RST(rst), .SENDING(SENDING), .SHIFT_ENABLE_R(
        SHIFT_ENABLE_R), .SHIFT_ENABLE_E(SHIFT_ENABLE_E) );
endmodule


module RMEDT_REWIRE_1 ( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN, DATA_IN, BS_ERROR, 
        CRC_ERROR, EMPTY, FULL, KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, 
        R_ERROR, SENDING, dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE, DATA, 
        ADDR );
  input [7:0] DATA_IN;
  output [7:0] DATA;
  output [7:0] ADDR;
  input CLK, DM1_RX, DP1_RX, RST, SERIAL_IN;
  output BS_ERROR, CRC_ERROR, EMPTY, FULL, KEY_ERROR, PROG_ERROR, PARITY_ERROR,
         RBUF_FULL, R_ERROR, SENDING, dm_tx_out, dp_tx_out, W_ENABLE_R,
         R_ENABLE;
  wire   B_READY, PDATA_READY, EOP_external, NEXT_BYTE, W_ENABLE;
  wire   [7:0] PRGA_IN;
  wire   [1:0] PRGA_OPCODE;
  wire   [7:0] PROCESSED_DATA;
  wire   [7:0] RCV_DATA;
  wire   [1:0] OPCODE;

  EDBlock_1 U_0 ( .BYTE(PRGA_IN), .BYTE_READY(B_READY), .CLK(CLK), .OPCODE(
        PRGA_OPCODE), .RST(RST), .SERIAL_IN(SERIAL_IN), .DATA_IN(DATA_IN), 
        .KEY_ERROR(KEY_ERROR), .PARITY_ERROR(PARITY_ERROR), .PDATA_READY(
        PDATA_READY), .PROCESSED_DATA(PROCESSED_DATA), .PROG_ERROR(PROG_ERROR), 
        .RBUF_FULL(RBUF_FULL), .W_ENABLE(W_ENABLE_R), .R_ENABLE(R_ENABLE), 
        .DATA(DATA), .ADDR(ADDR) );
  memoryblock_1 U_1 ( .CLK(CLK), .NEXT_BYTE(NEXT_BYTE), .RCV_DATA(RCV_DATA), 
        .RCV_OPCODE(OPCODE), .RST(RST), .W_ENABLE(W_ENABLE), .EOP(EOP_external), .EMPTY(EMPTY), .FULL(FULL), .B_READY(B_READY), .PRGA_IN(PRGA_IN), 
        .PRGA_OPCODE(PRGA_OPCODE) );
  receiver_block_rewire_1 U_2 ( .CLK(CLK), .DM1_RX(DM1_RX), .DP1_RX(DP1_RX), 
        .RST(RST), .BS_ERROR(BS_ERROR), .CRC_ERROR(CRC_ERROR), .EOP_external(
        EOP_external), .OPCODE(OPCODE), .RCV_DATA(RCV_DATA), .R_ERROR(R_ERROR), 
        .W_ENABLE(W_ENABLE) );
  transmitter_block_1 U_3 ( .PRGA_OUT(PROCESSED_DATA), .clk(CLK), .p_ready(
        PDATA_READY), .prga_opcode(PRGA_OPCODE), .rst(RST), .SENDING(SENDING), 
        .dm_tx_out(dm_tx_out), .dp_tx_out(dp_tx_out), .NEXT_BYTE(NEXT_BYTE) );
endmodule


module KSA_0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_0_DW01_add_6 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;

  AND2X2 U2 ( .A(n18), .B(n14), .Y(n1) );
  NAND2X1 U3 ( .A(n33), .B(n34), .Y(n19) );
  INVX2 U4 ( .A(n38), .Y(SUM[0]) );
  XNOR2X1 U5 ( .A(n2), .B(n3), .Y(SUM[7]) );
  XOR2X1 U6 ( .A(B[7]), .B(A[7]), .Y(n3) );
  AOI21X1 U7 ( .A(n4), .B(n5), .C(n6), .Y(n2) );
  INVX2 U8 ( .A(n7), .Y(n6) );
  XNOR2X1 U9 ( .A(n4), .B(n8), .Y(SUM[6]) );
  NAND2X1 U10 ( .A(n5), .B(n7), .Y(n8) );
  NAND2X1 U11 ( .A(B[6]), .B(A[6]), .Y(n7) );
  OR2X2 U12 ( .A(A[6]), .B(B[6]), .Y(n5) );
  NAND2X1 U13 ( .A(n9), .B(n10), .Y(n4) );
  NAND2X1 U14 ( .A(n11), .B(n12), .Y(n10) );
  XNOR2X1 U15 ( .A(n11), .B(n13), .Y(SUM[5]) );
  NAND2X1 U16 ( .A(n9), .B(n12), .Y(n13) );
  OR2X2 U17 ( .A(A[5]), .B(B[5]), .Y(n12) );
  NAND2X1 U18 ( .A(B[5]), .B(A[5]), .Y(n9) );
  NAND3X1 U19 ( .A(n14), .B(n15), .C(n16), .Y(n11) );
  NAND3X1 U20 ( .A(n17), .B(n18), .C(n19), .Y(n16) );
  INVX2 U21 ( .A(n20), .Y(n17) );
  NAND3X1 U22 ( .A(n21), .B(n18), .C(n22), .Y(n15) );
  XOR2X1 U23 ( .A(n23), .B(n1), .Y(SUM[4]) );
  NAND2X1 U24 ( .A(B[4]), .B(A[4]), .Y(n14) );
  OR2X2 U25 ( .A(A[4]), .B(B[4]), .Y(n18) );
  OAI21X1 U26 ( .A(n24), .B(n20), .C(n25), .Y(n23) );
  NAND2X1 U27 ( .A(n21), .B(n22), .Y(n25) );
  NAND2X1 U28 ( .A(n26), .B(n27), .Y(n22) );
  NAND2X1 U29 ( .A(n28), .B(n21), .Y(n20) );
  INVX2 U30 ( .A(n19), .Y(n24) );
  XNOR2X1 U31 ( .A(n29), .B(n30), .Y(SUM[3]) );
  AND2X2 U32 ( .A(n21), .B(n26), .Y(n30) );
  NAND2X1 U33 ( .A(B[3]), .B(A[3]), .Y(n26) );
  OR2X2 U34 ( .A(A[3]), .B(B[3]), .Y(n21) );
  AOI21X1 U35 ( .A(n19), .B(n28), .C(n31), .Y(n29) );
  INVX2 U36 ( .A(n27), .Y(n31) );
  XNOR2X1 U37 ( .A(n32), .B(n19), .Y(SUM[2]) );
  NAND3X1 U38 ( .A(A[0]), .B(B[0]), .C(n35), .Y(n34) );
  NAND2X1 U39 ( .A(n28), .B(n27), .Y(n32) );
  NAND2X1 U40 ( .A(B[2]), .B(A[2]), .Y(n27) );
  OR2X2 U41 ( .A(A[2]), .B(B[2]), .Y(n28) );
  XOR2X1 U42 ( .A(n36), .B(n37), .Y(SUM[1]) );
  NAND2X1 U43 ( .A(n35), .B(n33), .Y(n36) );
  NAND2X1 U44 ( .A(B[1]), .B(A[1]), .Y(n33) );
  OR2X2 U45 ( .A(A[1]), .B(B[1]), .Y(n35) );
  OAI21X1 U46 ( .A(A[0]), .B(B[0]), .C(n37), .Y(n38) );
  NAND2X1 U47 ( .A(B[0]), .B(A[0]), .Y(n37) );
endmodule


module KSA_0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  NAND2X1 U2 ( .A(n35), .B(n36), .Y(n30) );
  INVX2 U3 ( .A(n40), .Y(SUM[0]) );
  XNOR2X1 U4 ( .A(n1), .B(n2), .Y(SUM[7]) );
  XOR2X1 U5 ( .A(B[7]), .B(A[7]), .Y(n2) );
  AOI21X1 U6 ( .A(n3), .B(n4), .C(n5), .Y(n1) );
  INVX2 U7 ( .A(n6), .Y(n5) );
  XNOR2X1 U8 ( .A(n3), .B(n7), .Y(SUM[6]) );
  NAND2X1 U9 ( .A(n4), .B(n6), .Y(n7) );
  NAND2X1 U10 ( .A(B[6]), .B(A[6]), .Y(n6) );
  OR2X2 U11 ( .A(A[6]), .B(B[6]), .Y(n4) );
  NAND2X1 U12 ( .A(n8), .B(n9), .Y(n3) );
  NAND2X1 U13 ( .A(n10), .B(n11), .Y(n9) );
  XNOR2X1 U14 ( .A(n10), .B(n12), .Y(SUM[5]) );
  NAND2X1 U15 ( .A(n8), .B(n11), .Y(n12) );
  OR2X2 U16 ( .A(A[5]), .B(B[5]), .Y(n11) );
  NAND2X1 U17 ( .A(B[5]), .B(A[5]), .Y(n8) );
  OAI21X1 U18 ( .A(n13), .B(n14), .C(n15), .Y(n10) );
  AOI21X1 U19 ( .A(n16), .B(n17), .C(n18), .Y(n15) );
  INVX2 U20 ( .A(n19), .Y(n18) );
  INVX2 U21 ( .A(n20), .Y(n16) );
  NAND2X1 U22 ( .A(n21), .B(n17), .Y(n14) );
  INVX2 U23 ( .A(n22), .Y(n21) );
  XNOR2X1 U24 ( .A(n23), .B(n24), .Y(SUM[4]) );
  OAI21X1 U25 ( .A(n13), .B(n22), .C(n20), .Y(n24) );
  OAI21X1 U26 ( .A(n25), .B(n26), .C(n27), .Y(n20) );
  INVX2 U27 ( .A(n28), .Y(n26) );
  NAND2X1 U28 ( .A(n29), .B(n27), .Y(n22) );
  INVX2 U29 ( .A(n30), .Y(n13) );
  NAND2X1 U30 ( .A(n17), .B(n19), .Y(n23) );
  NAND2X1 U31 ( .A(B[4]), .B(A[4]), .Y(n19) );
  OR2X2 U32 ( .A(A[4]), .B(B[4]), .Y(n17) );
  XNOR2X1 U33 ( .A(n31), .B(n32), .Y(SUM[3]) );
  AND2X2 U34 ( .A(n27), .B(n28), .Y(n32) );
  NAND2X1 U35 ( .A(B[3]), .B(A[3]), .Y(n28) );
  OR2X2 U36 ( .A(A[3]), .B(B[3]), .Y(n27) );
  AOI21X1 U37 ( .A(n30), .B(n29), .C(n25), .Y(n31) );
  INVX2 U38 ( .A(n33), .Y(n25) );
  XNOR2X1 U39 ( .A(n34), .B(n30), .Y(SUM[2]) );
  NAND3X1 U40 ( .A(A[0]), .B(B[0]), .C(n37), .Y(n36) );
  NAND2X1 U41 ( .A(n29), .B(n33), .Y(n34) );
  NAND2X1 U42 ( .A(B[2]), .B(A[2]), .Y(n33) );
  OR2X2 U43 ( .A(A[2]), .B(B[2]), .Y(n29) );
  XOR2X1 U44 ( .A(n38), .B(n39), .Y(SUM[1]) );
  NAND2X1 U45 ( .A(n37), .B(n35), .Y(n38) );
  NAND2X1 U46 ( .A(B[1]), .B(A[1]), .Y(n35) );
  OR2X2 U47 ( .A(A[1]), .B(B[1]), .Y(n37) );
  OAI21X1 U48 ( .A(A[0]), .B(B[0]), .C(n39), .Y(n40) );
  NAND2X1 U49 ( .A(B[0]), .B(A[0]), .Y(n39) );
endmodule


module KSA_0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49;

  OAI21X1 U2 ( .A(n17), .B(n18), .C(n19), .Y(n1) );
  XNOR2X1 U3 ( .A(n6), .B(n10), .Y(SUM[6]) );
  XNOR2X1 U4 ( .A(n27), .B(n2), .Y(SUM[4]) );
  NAND2X1 U5 ( .A(n21), .B(n23), .Y(n2) );
  XOR2X1 U6 ( .A(n48), .B(n47), .Y(SUM[1]) );
  XOR2X1 U7 ( .A(n35), .B(n36), .Y(SUM[3]) );
  AND2X2 U8 ( .A(n33), .B(n31), .Y(n3) );
  INVX2 U9 ( .A(n39), .Y(n38) );
  NAND2X1 U10 ( .A(n45), .B(n42), .Y(n43) );
  INVX2 U11 ( .A(n49), .Y(SUM[0]) );
  XNOR2X1 U12 ( .A(n4), .B(n5), .Y(SUM[7]) );
  XOR2X1 U13 ( .A(B[7]), .B(A[7]), .Y(n5) );
  AOI21X1 U14 ( .A(n6), .B(n7), .C(n8), .Y(n4) );
  INVX2 U15 ( .A(n9), .Y(n8) );
  NAND2X1 U16 ( .A(n7), .B(n9), .Y(n10) );
  NAND2X1 U17 ( .A(B[6]), .B(A[6]), .Y(n9) );
  OR2X2 U18 ( .A(A[6]), .B(B[6]), .Y(n7) );
  OAI21X1 U19 ( .A(n11), .B(n12), .C(n13), .Y(n6) );
  INVX2 U20 ( .A(n14), .Y(n12) );
  INVX2 U21 ( .A(n15), .Y(n11) );
  XNOR2X1 U22 ( .A(n16), .B(n1), .Y(SUM[5]) );
  OAI21X1 U23 ( .A(n17), .B(n18), .C(n19), .Y(n14) );
  AOI21X1 U24 ( .A(n20), .B(n21), .C(n22), .Y(n19) );
  INVX2 U25 ( .A(n23), .Y(n22) );
  NAND2X1 U26 ( .A(n24), .B(n25), .Y(n20) );
  NAND3X1 U27 ( .A(n26), .B(n21), .C(n3), .Y(n18) );
  NAND2X1 U28 ( .A(n13), .B(n15), .Y(n16) );
  OR2X2 U29 ( .A(A[5]), .B(B[5]), .Y(n15) );
  NAND2X1 U30 ( .A(B[5]), .B(A[5]), .Y(n13) );
  NAND2X1 U31 ( .A(B[4]), .B(A[4]), .Y(n23) );
  OR2X2 U32 ( .A(A[4]), .B(B[4]), .Y(n21) );
  OAI21X1 U33 ( .A(n17), .B(n28), .C(n29), .Y(n27) );
  AND2X2 U34 ( .A(n24), .B(n25), .Y(n29) );
  NAND2X1 U35 ( .A(n30), .B(n31), .Y(n24) );
  INVX2 U36 ( .A(n32), .Y(n30) );
  NAND2X1 U37 ( .A(n3), .B(n26), .Y(n28) );
  AOI21X1 U38 ( .A(B[0]), .B(A[0]), .C(n34), .Y(n17) );
  NAND2X1 U39 ( .A(n25), .B(n31), .Y(n36) );
  OR2X2 U40 ( .A(A[3]), .B(B[3]), .Y(n31) );
  NAND2X1 U41 ( .A(B[3]), .B(A[3]), .Y(n25) );
  NOR2X1 U42 ( .A(n37), .B(n38), .Y(n35) );
  NAND3X1 U43 ( .A(n26), .B(n33), .C(n40), .Y(n39) );
  AND2X2 U44 ( .A(B[0]), .B(A[0]), .Y(n40) );
  NAND2X1 U45 ( .A(n41), .B(n32), .Y(n37) );
  NAND2X1 U46 ( .A(n34), .B(n33), .Y(n41) );
  INVX2 U47 ( .A(n42), .Y(n34) );
  XNOR2X1 U48 ( .A(n43), .B(n44), .Y(SUM[2]) );
  NAND2X1 U49 ( .A(n33), .B(n32), .Y(n44) );
  NAND2X1 U50 ( .A(B[2]), .B(A[2]), .Y(n32) );
  OR2X2 U51 ( .A(A[2]), .B(B[2]), .Y(n33) );
  NAND2X1 U52 ( .A(n46), .B(n26), .Y(n45) );
  AND2X2 U53 ( .A(A[0]), .B(B[0]), .Y(n46) );
  NAND2X1 U54 ( .A(n42), .B(n26), .Y(n47) );
  OR2X2 U55 ( .A(A[1]), .B(B[1]), .Y(n26) );
  NAND2X1 U56 ( .A(B[1]), .B(A[1]), .Y(n42) );
  OAI21X1 U57 ( .A(A[0]), .B(B[0]), .C(n48), .Y(n49) );
  NAND2X1 U58 ( .A(B[0]), .B(A[0]), .Y(n48) );
endmodule


module KSA_0_DW01_add_9 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59;

  INVX2 U2 ( .A(n17), .Y(n1) );
  INVX1 U3 ( .A(n5), .Y(n21) );
  AND2X2 U4 ( .A(n27), .B(n11), .Y(n2) );
  NAND2X1 U5 ( .A(n3), .B(n37), .Y(n15) );
  AND2X2 U6 ( .A(n38), .B(n39), .Y(n3) );
  AND2X2 U7 ( .A(B[0]), .B(A[0]), .Y(n4) );
  OAI21X1 U8 ( .A(B[6]), .B(A[6]), .C(n11), .Y(n5) );
  OR2X2 U9 ( .A(A[6]), .B(B[6]), .Y(n12) );
  INVX2 U10 ( .A(n37), .Y(n34) );
  INVX2 U11 ( .A(n59), .Y(SUM[0]) );
  XOR2X1 U12 ( .A(n6), .B(n7), .Y(SUM[7]) );
  XOR2X1 U13 ( .A(B[7]), .B(A[7]), .Y(n7) );
  NAND3X1 U14 ( .A(n8), .B(n9), .C(n10), .Y(n6) );
  NAND3X1 U15 ( .A(n11), .B(n12), .C(n13), .Y(n10) );
  NAND3X1 U16 ( .A(n14), .B(n11), .C(n15), .Y(n9) );
  AOI21X1 U17 ( .A(n16), .B(n17), .C(n18), .Y(n14) );
  NAND2X1 U18 ( .A(n19), .B(n20), .Y(n18) );
  INVX2 U19 ( .A(B[6]), .Y(n17) );
  INVX2 U20 ( .A(A[6]), .Y(n16) );
  AOI21X1 U21 ( .A(n21), .B(n22), .C(n23), .Y(n8) );
  NAND2X1 U22 ( .A(n24), .B(n25), .Y(n23) );
  OAI21X1 U23 ( .A(A[6]), .B(B[6]), .C(n26), .Y(n25) );
  INVX2 U24 ( .A(n27), .Y(n26) );
  XOR2X1 U25 ( .A(n28), .B(n29), .Y(SUM[6]) );
  INVX2 U26 ( .A(n30), .Y(n29) );
  OAI21X1 U27 ( .A(n1), .B(A[6]), .C(n24), .Y(n30) );
  NAND2X1 U28 ( .A(B[6]), .B(A[6]), .Y(n24) );
  NAND3X1 U29 ( .A(n27), .B(n31), .C(n32), .Y(n28) );
  OAI21X1 U30 ( .A(n33), .B(n34), .C(n35), .Y(n32) );
  AND2X2 U31 ( .A(n36), .B(n11), .Y(n35) );
  NAND2X1 U32 ( .A(n38), .B(n39), .Y(n33) );
  AOI22X1 U33 ( .A(n22), .B(n11), .C(n13), .D(n11), .Y(n31) );
  INVX2 U34 ( .A(n40), .Y(n13) );
  INVX2 U35 ( .A(n41), .Y(n22) );
  XNOR2X1 U36 ( .A(n42), .B(n2), .Y(SUM[5]) );
  OR2X2 U37 ( .A(A[5]), .B(B[5]), .Y(n11) );
  NAND2X1 U38 ( .A(B[5]), .B(A[5]), .Y(n27) );
  AOI21X1 U39 ( .A(n36), .B(n15), .C(n43), .Y(n42) );
  NAND2X1 U40 ( .A(n40), .B(n41), .Y(n43) );
  NAND3X1 U41 ( .A(A[3]), .B(B[3]), .C(n19), .Y(n40) );
  INVX2 U42 ( .A(n44), .Y(n36) );
  OAI21X1 U43 ( .A(A[4]), .B(B[4]), .C(n20), .Y(n44) );
  XNOR2X1 U44 ( .A(n45), .B(n46), .Y(SUM[4]) );
  AND2X2 U45 ( .A(n19), .B(n41), .Y(n46) );
  NAND2X1 U46 ( .A(B[4]), .B(A[4]), .Y(n41) );
  OR2X2 U47 ( .A(A[4]), .B(B[4]), .Y(n19) );
  AOI21X1 U48 ( .A(n15), .B(n20), .C(n47), .Y(n45) );
  INVX2 U49 ( .A(n48), .Y(n47) );
  XNOR2X1 U50 ( .A(n15), .B(n49), .Y(SUM[3]) );
  NAND2X1 U51 ( .A(n20), .B(n48), .Y(n49) );
  NAND2X1 U52 ( .A(B[3]), .B(A[3]), .Y(n48) );
  OR2X2 U53 ( .A(A[3]), .B(B[3]), .Y(n20) );
  NAND3X1 U54 ( .A(n50), .B(n51), .C(n52), .Y(n37) );
  AND2X2 U55 ( .A(B[0]), .B(A[0]), .Y(n52) );
  NAND3X1 U56 ( .A(A[1]), .B(B[1]), .C(n51), .Y(n38) );
  XOR2X1 U57 ( .A(n53), .B(n54), .Y(SUM[2]) );
  AOI21X1 U58 ( .A(n4), .B(n50), .C(n55), .Y(n54) );
  INVX2 U59 ( .A(n56), .Y(n55) );
  NAND2X1 U60 ( .A(n51), .B(n39), .Y(n53) );
  NAND2X1 U61 ( .A(B[2]), .B(A[2]), .Y(n39) );
  OR2X2 U62 ( .A(A[2]), .B(B[2]), .Y(n51) );
  XNOR2X1 U63 ( .A(n57), .B(n4), .Y(SUM[1]) );
  NAND2X1 U64 ( .A(n50), .B(n56), .Y(n57) );
  NAND2X1 U65 ( .A(B[1]), .B(A[1]), .Y(n56) );
  OR2X2 U66 ( .A(A[1]), .B(B[1]), .Y(n50) );
  OAI21X1 U67 ( .A(A[0]), .B(B[0]), .C(n58), .Y(n59) );
  NAND2X1 U68 ( .A(B[0]), .B(A[0]), .Y(n58) );
endmodule


module KSA_0_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  XOR2X1 U2 ( .A(n3), .B(A[6]), .Y(SUM[6]) );
  XOR2X1 U3 ( .A(n5), .B(A[4]), .Y(SUM[4]) );
  AND2X2 U4 ( .A(A[1]), .B(A[0]), .Y(n1) );
  XOR2X1 U5 ( .A(n1), .B(A[2]), .Y(SUM[2]) );
  XNOR2X1 U6 ( .A(A[7]), .B(n2), .Y(SUM[7]) );
  NAND2X1 U7 ( .A(A[6]), .B(n3), .Y(n2) );
  INVX2 U8 ( .A(n4), .Y(n3) );
  NAND3X1 U9 ( .A(A[4]), .B(A[5]), .C(n5), .Y(n4) );
  XNOR2X1 U10 ( .A(A[5]), .B(n6), .Y(SUM[5]) );
  NAND2X1 U11 ( .A(A[4]), .B(n5), .Y(n6) );
  INVX2 U12 ( .A(n7), .Y(n5) );
  NAND3X1 U13 ( .A(A[2]), .B(A[3]), .C(n1), .Y(n7) );
  XNOR2X1 U14 ( .A(A[3]), .B(n8), .Y(SUM[3]) );
  NAND2X1 U15 ( .A(A[2]), .B(n1), .Y(n8) );
  XOR2X1 U16 ( .A(A[1]), .B(A[0]), .Y(SUM[1]) );
  INVX2 U17 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module KSA_0 ( KEY, CLK, RST, KEY_ERROR, BYTE_READY, BYTE, OPCODE, DATA_IN, 
        PROCESSED_DATA, PDATA_READY, W_ENABLE, R_ENABLE, ADDR, DATA );
  input [63:0] KEY;
  input [7:0] BYTE;
  input [1:0] OPCODE;
  input [7:0] DATA_IN;
  output [7:0] PROCESSED_DATA;
  output [7:0] ADDR;
  output [7:0] DATA;
  input CLK, RST, KEY_ERROR, BYTE_READY;
  output PDATA_READY, W_ENABLE, R_ENABLE;
  wire   permuteComplete, \keyTable[0][7] , \keyTable[0][6] , \keyTable[0][5] ,
         \keyTable[0][4] , \keyTable[0][3] , \keyTable[0][2] ,
         \keyTable[0][1] , \keyTable[0][0] , \keyTable[1][7] ,
         \keyTable[1][6] , \keyTable[1][5] , \keyTable[1][4] ,
         \keyTable[1][3] , \keyTable[1][2] , \keyTable[1][1] ,
         \keyTable[1][0] , \keyTable[2][7] , \keyTable[2][6] ,
         \keyTable[2][5] , \keyTable[2][4] , \keyTable[2][3] ,
         \keyTable[2][2] , \keyTable[2][1] , \keyTable[2][0] ,
         \keyTable[3][7] , \keyTable[3][6] , \keyTable[3][5] ,
         \keyTable[3][4] , \keyTable[3][3] , \keyTable[3][2] ,
         \keyTable[3][1] , \keyTable[3][0] , \keyTable[4][7] ,
         \keyTable[4][6] , \keyTable[4][5] , \keyTable[4][4] ,
         \keyTable[4][3] , \keyTable[4][2] , \keyTable[4][1] ,
         \keyTable[4][0] , \keyTable[5][7] , \keyTable[5][6] ,
         \keyTable[5][5] , \keyTable[5][4] , \keyTable[5][3] ,
         \keyTable[5][2] , \keyTable[5][1] , \keyTable[5][0] ,
         \keyTable[6][7] , \keyTable[6][6] , \keyTable[6][5] ,
         \keyTable[6][4] , \keyTable[6][3] , \keyTable[6][2] ,
         \keyTable[6][1] , \keyTable[6][0] , \keyTable[7][7] ,
         \keyTable[7][6] , \keyTable[7][5] , \keyTable[7][4] ,
         \keyTable[7][3] , \keyTable[7][2] , \keyTable[7][1] ,
         \keyTable[7][0] , fw_enable, fr_enable, N407, N408, N409, N410, N411,
         N412, N413, N414, N424, N425, N426, N427, N428, N429, N430, N431,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N496, N497, N498, N499, N500, N501,
         N502, N503, N512, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N522, N523, N524, N525, N526, N527, N456, N455, N454, N453,
         N452, N451, N450, N449, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n125, n127, n129, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n156, n157, n160, n161,
         n162, n164, n166, n167, n169, n170, n171, n172, n175, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n692, n701, n746, n748, n750, n752, n754, n756, n758,
         n760, n765, n766, n767, n768, n769, n771, n772, n773, n774, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n864, n865, n866,
         n867, n868, n869, n870, n871, n883, n884, n885, n886, n887, n888,
         n889, n890, n898, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
  wire   [4:0] state;
  wire   [7:0] si;
  wire   [7:0] sj;
  wire   [7:0] currentProcessedData;
  wire   [4:0] nextState;
  wire   [7:0] inti;
  wire   [7:0] intj;
  wire   [2:0] keyi;
  wire   [7:0] temp;
  wire   [7:0] extratemp;
  wire   [7:0] nextProcessedData;
  wire   [7:0] delaydata;
  wire   [7:0] prefillCounter;
  wire   [7:0] faddr;
  wire   [7:0] fdata;
  tri   [7:0] nfaddr;
  tri   [7:0] nfdata;

  DFFPOSX1 \prefillCounter_reg[0]  ( .D(n1138), .CLK(CLK), .Q(
        prefillCounter[0]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n242), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n242), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[4]  ( .D(nextState[4]), .CLK(CLK), .R(n241), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n241), .S(1'b1), .Q(
        state[0]) );
  DFFPOSX1 permuteComplete_reg ( .D(n1154), .CLK(CLK), .Q(permuteComplete) );
  DFFSR \state_reg[3]  ( .D(nextState[3]), .CLK(CLK), .R(n241), .S(1'b1), .Q(
        state[3]) );
  DFFSR PDATA_READY_reg ( .D(n1134), .CLK(CLK), .R(n241), .S(1'b1), .Q(
        PDATA_READY) );
  DFFPOSX1 \extratemp_reg[7]  ( .D(n1133), .CLK(CLK), .Q(extratemp[7]) );
  DFFPOSX1 \extratemp_reg[6]  ( .D(n1132), .CLK(CLK), .Q(extratemp[6]) );
  DFFPOSX1 \extratemp_reg[5]  ( .D(n1131), .CLK(CLK), .Q(extratemp[5]) );
  DFFPOSX1 \extratemp_reg[4]  ( .D(n1130), .CLK(CLK), .Q(extratemp[4]) );
  DFFPOSX1 \extratemp_reg[3]  ( .D(n1129), .CLK(CLK), .Q(extratemp[3]) );
  DFFPOSX1 \extratemp_reg[2]  ( .D(n1128), .CLK(CLK), .Q(extratemp[2]) );
  DFFPOSX1 \extratemp_reg[1]  ( .D(n1127), .CLK(CLK), .Q(extratemp[1]) );
  DFFPOSX1 \extratemp_reg[0]  ( .D(n1126), .CLK(CLK), .Q(extratemp[0]) );
  DFFPOSX1 \keyTable_reg[7][0]  ( .D(n1244), .CLK(CLK), .Q(\keyTable[7][0] )
         );
  DFFPOSX1 \keyTable_reg[7][1]  ( .D(n1243), .CLK(CLK), .Q(\keyTable[7][1] )
         );
  DFFPOSX1 \keyTable_reg[7][2]  ( .D(n1242), .CLK(CLK), .Q(\keyTable[7][2] )
         );
  DFFPOSX1 \keyTable_reg[7][3]  ( .D(n1241), .CLK(CLK), .Q(\keyTable[7][3] )
         );
  DFFPOSX1 \keyTable_reg[7][4]  ( .D(n1240), .CLK(CLK), .Q(\keyTable[7][4] )
         );
  DFFPOSX1 \keyTable_reg[7][5]  ( .D(n1239), .CLK(CLK), .Q(\keyTable[7][5] )
         );
  DFFPOSX1 \keyTable_reg[7][6]  ( .D(n1238), .CLK(CLK), .Q(\keyTable[7][6] )
         );
  DFFPOSX1 \keyTable_reg[7][7]  ( .D(n1237), .CLK(CLK), .Q(\keyTable[7][7] )
         );
  DFFPOSX1 \keyTable_reg[6][0]  ( .D(n1236), .CLK(CLK), .Q(\keyTable[6][0] )
         );
  DFFPOSX1 \keyTable_reg[6][1]  ( .D(n1235), .CLK(CLK), .Q(\keyTable[6][1] )
         );
  DFFPOSX1 \keyTable_reg[6][2]  ( .D(n1234), .CLK(CLK), .Q(\keyTable[6][2] )
         );
  DFFPOSX1 \keyTable_reg[6][3]  ( .D(n1233), .CLK(CLK), .Q(\keyTable[6][3] )
         );
  DFFPOSX1 \keyTable_reg[6][4]  ( .D(n1232), .CLK(CLK), .Q(\keyTable[6][4] )
         );
  DFFPOSX1 \keyTable_reg[6][5]  ( .D(n1231), .CLK(CLK), .Q(\keyTable[6][5] )
         );
  DFFPOSX1 \keyTable_reg[6][6]  ( .D(n1230), .CLK(CLK), .Q(\keyTable[6][6] )
         );
  DFFPOSX1 \keyTable_reg[6][7]  ( .D(n1229), .CLK(CLK), .Q(\keyTable[6][7] )
         );
  DFFPOSX1 \keyTable_reg[5][0]  ( .D(n1228), .CLK(CLK), .Q(\keyTable[5][0] )
         );
  DFFPOSX1 \keyTable_reg[5][1]  ( .D(n1227), .CLK(CLK), .Q(\keyTable[5][1] )
         );
  DFFPOSX1 \keyTable_reg[5][2]  ( .D(n1226), .CLK(CLK), .Q(\keyTable[5][2] )
         );
  DFFPOSX1 \keyTable_reg[5][3]  ( .D(n1225), .CLK(CLK), .Q(\keyTable[5][3] )
         );
  DFFPOSX1 \keyTable_reg[5][4]  ( .D(n1224), .CLK(CLK), .Q(\keyTable[5][4] )
         );
  DFFPOSX1 \keyTable_reg[5][5]  ( .D(n1223), .CLK(CLK), .Q(\keyTable[5][5] )
         );
  DFFPOSX1 \keyTable_reg[5][6]  ( .D(n1222), .CLK(CLK), .Q(\keyTable[5][6] )
         );
  DFFPOSX1 \keyTable_reg[5][7]  ( .D(n1221), .CLK(CLK), .Q(\keyTable[5][7] )
         );
  DFFPOSX1 \keyTable_reg[4][0]  ( .D(n1220), .CLK(CLK), .Q(\keyTable[4][0] )
         );
  DFFPOSX1 \keyTable_reg[4][1]  ( .D(n1219), .CLK(CLK), .Q(\keyTable[4][1] )
         );
  DFFPOSX1 \keyTable_reg[4][2]  ( .D(n1218), .CLK(CLK), .Q(\keyTable[4][2] )
         );
  DFFPOSX1 \keyTable_reg[4][3]  ( .D(n1217), .CLK(CLK), .Q(\keyTable[4][3] )
         );
  DFFPOSX1 \keyTable_reg[4][4]  ( .D(n1216), .CLK(CLK), .Q(\keyTable[4][4] )
         );
  DFFPOSX1 \keyTable_reg[4][5]  ( .D(n1215), .CLK(CLK), .Q(\keyTable[4][5] )
         );
  DFFPOSX1 \keyTable_reg[4][6]  ( .D(n1214), .CLK(CLK), .Q(\keyTable[4][6] )
         );
  DFFPOSX1 \keyTable_reg[4][7]  ( .D(n1213), .CLK(CLK), .Q(\keyTable[4][7] )
         );
  DFFPOSX1 \keyTable_reg[3][0]  ( .D(n1212), .CLK(CLK), .Q(\keyTable[3][0] )
         );
  DFFPOSX1 \keyTable_reg[3][1]  ( .D(n1211), .CLK(CLK), .Q(\keyTable[3][1] )
         );
  DFFPOSX1 \keyTable_reg[3][2]  ( .D(n1210), .CLK(CLK), .Q(\keyTable[3][2] )
         );
  DFFPOSX1 \keyTable_reg[3][3]  ( .D(n1209), .CLK(CLK), .Q(\keyTable[3][3] )
         );
  DFFPOSX1 \keyTable_reg[3][4]  ( .D(n1208), .CLK(CLK), .Q(\keyTable[3][4] )
         );
  DFFPOSX1 \keyTable_reg[3][5]  ( .D(n1207), .CLK(CLK), .Q(\keyTable[3][5] )
         );
  DFFPOSX1 \keyTable_reg[3][6]  ( .D(n1206), .CLK(CLK), .Q(\keyTable[3][6] )
         );
  DFFPOSX1 \keyTable_reg[3][7]  ( .D(n1205), .CLK(CLK), .Q(\keyTable[3][7] )
         );
  DFFPOSX1 \keyTable_reg[2][0]  ( .D(n1204), .CLK(CLK), .Q(\keyTable[2][0] )
         );
  DFFPOSX1 \keyTable_reg[2][1]  ( .D(n1203), .CLK(CLK), .Q(\keyTable[2][1] )
         );
  DFFPOSX1 \keyTable_reg[2][2]  ( .D(n1202), .CLK(CLK), .Q(\keyTable[2][2] )
         );
  DFFPOSX1 \keyTable_reg[2][3]  ( .D(n1201), .CLK(CLK), .Q(\keyTable[2][3] )
         );
  DFFPOSX1 \keyTable_reg[2][4]  ( .D(n1200), .CLK(CLK), .Q(\keyTable[2][4] )
         );
  DFFPOSX1 \keyTable_reg[2][5]  ( .D(n1199), .CLK(CLK), .Q(\keyTable[2][5] )
         );
  DFFPOSX1 \keyTable_reg[2][6]  ( .D(n1198), .CLK(CLK), .Q(\keyTable[2][6] )
         );
  DFFPOSX1 \keyTable_reg[2][7]  ( .D(n1197), .CLK(CLK), .Q(\keyTable[2][7] )
         );
  DFFPOSX1 \keyTable_reg[1][0]  ( .D(n1196), .CLK(CLK), .Q(\keyTable[1][0] )
         );
  DFFPOSX1 \keyTable_reg[1][1]  ( .D(n1195), .CLK(CLK), .Q(\keyTable[1][1] )
         );
  DFFPOSX1 \keyTable_reg[1][2]  ( .D(n1194), .CLK(CLK), .Q(\keyTable[1][2] )
         );
  DFFPOSX1 \keyTable_reg[1][3]  ( .D(n1193), .CLK(CLK), .Q(\keyTable[1][3] )
         );
  DFFPOSX1 \keyTable_reg[1][4]  ( .D(n1192), .CLK(CLK), .Q(\keyTable[1][4] )
         );
  DFFPOSX1 \keyTable_reg[1][5]  ( .D(n1191), .CLK(CLK), .Q(\keyTable[1][5] )
         );
  DFFPOSX1 \keyTable_reg[1][6]  ( .D(n1190), .CLK(CLK), .Q(\keyTable[1][6] )
         );
  DFFPOSX1 \keyTable_reg[0][6]  ( .D(n1189), .CLK(CLK), .Q(\keyTable[0][6] )
         );
  DFFPOSX1 \keyTable_reg[0][5]  ( .D(n1188), .CLK(CLK), .Q(\keyTable[0][5] )
         );
  DFFPOSX1 \keyTable_reg[0][4]  ( .D(n1187), .CLK(CLK), .Q(\keyTable[0][4] )
         );
  DFFPOSX1 \keyTable_reg[0][3]  ( .D(n1186), .CLK(CLK), .Q(\keyTable[0][3] )
         );
  DFFPOSX1 \keyTable_reg[0][2]  ( .D(n1185), .CLK(CLK), .Q(\keyTable[0][2] )
         );
  DFFPOSX1 \keyTable_reg[0][1]  ( .D(n1184), .CLK(CLK), .Q(\keyTable[0][1] )
         );
  DFFPOSX1 \keyTable_reg[0][0]  ( .D(n1183), .CLK(CLK), .Q(\keyTable[0][0] )
         );
  DFFPOSX1 \keyTable_reg[1][7]  ( .D(n1182), .CLK(CLK), .Q(\keyTable[1][7] )
         );
  DFFPOSX1 \keyTable_reg[0][7]  ( .D(n1181), .CLK(CLK), .Q(\keyTable[0][7] )
         );
  DFFPOSX1 \prefillCounter_reg[7]  ( .D(n1139), .CLK(CLK), .Q(
        prefillCounter[7]) );
  DFFPOSX1 \prefillCounter_reg[1]  ( .D(n1140), .CLK(CLK), .Q(
        prefillCounter[1]) );
  DFFPOSX1 \prefillCounter_reg[2]  ( .D(n1141), .CLK(CLK), .Q(
        prefillCounter[2]) );
  DFFPOSX1 \prefillCounter_reg[3]  ( .D(n1142), .CLK(CLK), .Q(
        prefillCounter[3]) );
  DFFPOSX1 \prefillCounter_reg[4]  ( .D(n1143), .CLK(CLK), .Q(
        prefillCounter[4]) );
  DFFPOSX1 \prefillCounter_reg[5]  ( .D(n1144), .CLK(CLK), .Q(
        prefillCounter[5]) );
  DFFPOSX1 \prefillCounter_reg[6]  ( .D(n1145), .CLK(CLK), .Q(
        prefillCounter[6]) );
  DFFPOSX1 \temp_reg[7]  ( .D(n1180), .CLK(CLK), .Q(temp[7]) );
  DFFPOSX1 \temp_reg[0]  ( .D(n1173), .CLK(CLK), .Q(temp[0]) );
  DFFPOSX1 \temp_reg[1]  ( .D(n1174), .CLK(CLK), .Q(temp[1]) );
  DFFPOSX1 \temp_reg[2]  ( .D(n1175), .CLK(CLK), .Q(temp[2]) );
  DFFPOSX1 \temp_reg[3]  ( .D(n1176), .CLK(CLK), .Q(temp[3]) );
  DFFPOSX1 \temp_reg[4]  ( .D(n1177), .CLK(CLK), .Q(temp[4]) );
  DFFPOSX1 \temp_reg[5]  ( .D(n1178), .CLK(CLK), .Q(temp[5]) );
  DFFPOSX1 \temp_reg[6]  ( .D(n1179), .CLK(CLK), .Q(temp[6]) );
  DFFSR \si_reg[0]  ( .D(n1146), .CLK(CLK), .R(n241), .S(1'b1), .Q(si[0]) );
  DFFSR \si_reg[1]  ( .D(n1147), .CLK(CLK), .R(n240), .S(1'b1), .Q(si[1]) );
  DFFSR \si_reg[6]  ( .D(n1152), .CLK(CLK), .R(n240), .S(1'b1), .Q(si[6]) );
  DFFPOSX1 \delaydata_reg[7]  ( .D(n1110), .CLK(CLK), .Q(delaydata[7]) );
  DFFPOSX1 \delaydata_reg[0]  ( .D(n1117), .CLK(CLK), .Q(delaydata[0]) );
  DFFPOSX1 \delaydata_reg[1]  ( .D(n1116), .CLK(CLK), .Q(delaydata[1]) );
  DFFPOSX1 \delaydata_reg[2]  ( .D(n1115), .CLK(CLK), .Q(delaydata[2]) );
  DFFPOSX1 \delaydata_reg[3]  ( .D(n1114), .CLK(CLK), .Q(delaydata[3]) );
  DFFPOSX1 \delaydata_reg[4]  ( .D(n1113), .CLK(CLK), .Q(delaydata[4]) );
  DFFPOSX1 \delaydata_reg[5]  ( .D(n1112), .CLK(CLK), .Q(delaydata[5]) );
  DFFPOSX1 \delaydata_reg[6]  ( .D(n1111), .CLK(CLK), .Q(delaydata[6]) );
  DFFPOSX1 \intj_reg[7]  ( .D(n1169), .CLK(CLK), .Q(intj[7]) );
  DFFPOSX1 \intj_reg[0]  ( .D(n1162), .CLK(CLK), .Q(intj[0]) );
  DFFPOSX1 \intj_reg[1]  ( .D(n1163), .CLK(CLK), .Q(intj[1]) );
  DFFPOSX1 \intj_reg[2]  ( .D(n1164), .CLK(CLK), .Q(intj[2]) );
  DFFPOSX1 \intj_reg[3]  ( .D(n1165), .CLK(CLK), .Q(intj[3]) );
  DFFPOSX1 \intj_reg[4]  ( .D(n1166), .CLK(CLK), .Q(intj[4]) );
  DFFPOSX1 \intj_reg[5]  ( .D(n1167), .CLK(CLK), .Q(intj[5]) );
  DFFPOSX1 \intj_reg[6]  ( .D(n1168), .CLK(CLK), .Q(intj[6]) );
  DFFSR \sj_reg[3]  ( .D(n1158), .CLK(CLK), .R(n239), .S(1'b1), .Q(sj[3]) );
  DFFSR \sj_reg[2]  ( .D(n1159), .CLK(CLK), .R(n239), .S(1'b1), .Q(sj[2]) );
  DFFSR \sj_reg[1]  ( .D(n1160), .CLK(CLK), .R(n239), .S(1'b1), .Q(sj[1]) );
  DFFSR \sj_reg[0]  ( .D(n1161), .CLK(CLK), .R(n236), .S(1'b1), .Q(sj[0]) );
  DFFPOSX1 \keyi_reg[2]  ( .D(n1170), .CLK(CLK), .Q(keyi[2]) );
  DFFPOSX1 \keyi_reg[1]  ( .D(n1171), .CLK(CLK), .Q(keyi[1]) );
  DFFPOSX1 \keyi_reg[0]  ( .D(n1172), .CLK(CLK), .Q(keyi[0]) );
  DFFPOSX1 \inti_reg[7]  ( .D(n1125), .CLK(CLK), .Q(inti[7]) );
  DFFPOSX1 \inti_reg[0]  ( .D(n1118), .CLK(CLK), .Q(inti[0]) );
  DFFPOSX1 \inti_reg[1]  ( .D(n1119), .CLK(CLK), .Q(inti[1]) );
  DFFPOSX1 \inti_reg[2]  ( .D(n1120), .CLK(CLK), .Q(inti[2]) );
  DFFPOSX1 \inti_reg[3]  ( .D(n1121), .CLK(CLK), .Q(inti[3]) );
  DFFPOSX1 \inti_reg[4]  ( .D(n1122), .CLK(CLK), .Q(inti[4]) );
  DFFPOSX1 \inti_reg[5]  ( .D(n1123), .CLK(CLK), .Q(inti[5]) );
  DFFPOSX1 \inti_reg[6]  ( .D(n1124), .CLK(CLK), .Q(inti[6]) );
  DFFPOSX1 \PROCESSED_DATA_reg[0]  ( .D(n1258), .CLK(CLK), .Q(
        PROCESSED_DATA[0]) );
  DFFPOSX1 \PROCESSED_DATA_reg[1]  ( .D(n1259), .CLK(CLK), .Q(
        PROCESSED_DATA[1]) );
  DFFPOSX1 \PROCESSED_DATA_reg[2]  ( .D(n1260), .CLK(CLK), .Q(
        PROCESSED_DATA[2]) );
  DFFPOSX1 \PROCESSED_DATA_reg[3]  ( .D(n1261), .CLK(CLK), .Q(
        PROCESSED_DATA[3]) );
  DFFPOSX1 \PROCESSED_DATA_reg[4]  ( .D(n1262), .CLK(CLK), .Q(
        PROCESSED_DATA[4]) );
  DFFPOSX1 \PROCESSED_DATA_reg[5]  ( .D(n1263), .CLK(CLK), .Q(
        PROCESSED_DATA[5]) );
  DFFPOSX1 \PROCESSED_DATA_reg[6]  ( .D(n1264), .CLK(CLK), .Q(
        PROCESSED_DATA[6]) );
  DFFPOSX1 \PROCESSED_DATA_reg[7]  ( .D(n1265), .CLK(CLK), .Q(
        PROCESSED_DATA[7]) );
  DFFPOSX1 \faddr_reg[7]  ( .D(n1266), .CLK(CLK), .Q(faddr[7]) );
  DFFPOSX1 \ADDR_reg[7]  ( .D(n1267), .CLK(CLK), .Q(ADDR[7]) );
  DFFPOSX1 \faddr_reg[6]  ( .D(n1268), .CLK(CLK), .Q(faddr[6]) );
  DFFPOSX1 \ADDR_reg[6]  ( .D(n1269), .CLK(CLK), .Q(ADDR[6]) );
  DFFPOSX1 \faddr_reg[5]  ( .D(n1270), .CLK(CLK), .Q(faddr[5]) );
  DFFPOSX1 \ADDR_reg[5]  ( .D(n1271), .CLK(CLK), .Q(ADDR[5]) );
  DFFPOSX1 \faddr_reg[4]  ( .D(n1272), .CLK(CLK), .Q(faddr[4]) );
  DFFPOSX1 \ADDR_reg[4]  ( .D(n1273), .CLK(CLK), .Q(ADDR[4]) );
  DFFPOSX1 \faddr_reg[3]  ( .D(n1274), .CLK(CLK), .Q(faddr[3]) );
  DFFPOSX1 \ADDR_reg[3]  ( .D(n1275), .CLK(CLK), .Q(ADDR[3]) );
  DFFPOSX1 \faddr_reg[2]  ( .D(n1276), .CLK(CLK), .Q(faddr[2]) );
  DFFPOSX1 \ADDR_reg[2]  ( .D(n1277), .CLK(CLK), .Q(ADDR[2]) );
  DFFPOSX1 \faddr_reg[1]  ( .D(n1278), .CLK(CLK), .Q(faddr[1]) );
  DFFPOSX1 \ADDR_reg[1]  ( .D(n1279), .CLK(CLK), .Q(ADDR[1]) );
  DFFPOSX1 \faddr_reg[0]  ( .D(n1280), .CLK(CLK), .Q(faddr[0]) );
  DFFPOSX1 \ADDR_reg[0]  ( .D(n1281), .CLK(CLK), .Q(ADDR[0]) );
  DFFPOSX1 \fdata_reg[7]  ( .D(n1282), .CLK(CLK), .Q(fdata[7]) );
  DFFPOSX1 \fdata_reg[6]  ( .D(n1283), .CLK(CLK), .Q(fdata[6]) );
  DFFPOSX1 \fdata_reg[5]  ( .D(n1284), .CLK(CLK), .Q(fdata[5]) );
  DFFPOSX1 \fdata_reg[4]  ( .D(n1285), .CLK(CLK), .Q(fdata[4]) );
  DFFPOSX1 \fdata_reg[3]  ( .D(n1286), .CLK(CLK), .Q(fdata[3]) );
  DFFPOSX1 \fdata_reg[2]  ( .D(n1287), .CLK(CLK), .Q(fdata[2]) );
  DFFPOSX1 \fdata_reg[1]  ( .D(n1288), .CLK(CLK), .Q(fdata[1]) );
  DFFPOSX1 \fdata_reg[0]  ( .D(n1289), .CLK(CLK), .Q(fdata[0]) );
  DFFPOSX1 fw_enable_reg ( .D(n1290), .CLK(CLK), .Q(fw_enable) );
  DFFPOSX1 fr_enable_reg ( .D(n1291), .CLK(CLK), .Q(fr_enable) );
  DFFPOSX1 W_ENABLE_reg ( .D(n1292), .CLK(CLK), .Q(W_ENABLE) );
  DFFPOSX1 R_ENABLE_reg ( .D(n1293), .CLK(CLK), .Q(R_ENABLE) );
  DFFPOSX1 \DATA_reg[7]  ( .D(n1294), .CLK(CLK), .Q(DATA[7]) );
  DFFPOSX1 \DATA_reg[6]  ( .D(n1295), .CLK(CLK), .Q(DATA[6]) );
  DFFPOSX1 \DATA_reg[5]  ( .D(n1296), .CLK(CLK), .Q(DATA[5]) );
  DFFPOSX1 \DATA_reg[4]  ( .D(n1297), .CLK(CLK), .Q(DATA[4]) );
  DFFPOSX1 \DATA_reg[3]  ( .D(n1298), .CLK(CLK), .Q(DATA[3]) );
  DFFPOSX1 \DATA_reg[2]  ( .D(n1299), .CLK(CLK), .Q(DATA[2]) );
  DFFPOSX1 \DATA_reg[1]  ( .D(n1300), .CLK(CLK), .Q(DATA[1]) );
  DFFPOSX1 \DATA_reg[0]  ( .D(n1301), .CLK(CLK), .Q(DATA[0]) );
  NOR2X1 U110 ( .A(KEY_ERROR), .B(n1332), .Y(n1333) );
  OAI21X1 U111 ( .A(n1106), .B(n1331), .C(n1105), .Y(n1334) );
  NOR2X1 U123 ( .A(n1328), .B(n1106), .Y(n1330) );
  NAND3X1 U126 ( .A(n1327), .B(n1100), .C(n1326), .Y(nextState[1]) );
  NOR2X1 U130 ( .A(prefillCounter[2]), .B(prefillCounter[1]), .Y(n1324) );
  NAND3X1 U131 ( .A(n1323), .B(n1135), .C(n1322), .Y(n1325) );
  NOR2X1 U132 ( .A(prefillCounter[4]), .B(prefillCounter[3]), .Y(n1322) );
  NOR2X1 U133 ( .A(prefillCounter[7]), .B(prefillCounter[6]), .Y(n1323) );
  NAND3X1 U143 ( .A(n1109), .B(n1108), .C(BYTE_READY), .Y(n1329) );
  NAND2X1 U156 ( .A(OPCODE[0]), .B(n1108), .Y(n1331) );
  NAND2X1 U158 ( .A(BYTE_READY), .B(n1320), .Y(n1332) );
  OAI21X1 U159 ( .A(OPCODE[0]), .B(OPCODE[1]), .C(n1321), .Y(n1320) );
  NAND2X1 U160 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n1321) );
  NOR2X1 U669 ( .A(n1103), .B(n1104), .Y(n1319) );
  NOR2X1 U673 ( .A(n1101), .B(n1102), .Y(n1318) );
  AND2X2 U142 ( .A(n1331), .B(n1321), .Y(n1328) );
  KSA_0_DW01_inc_0 add_289 ( .A(si), .SUM({N431, N430, N429, N428, N427, N426, 
        N425, N424}) );
  KSA_0_DW01_inc_1 add_263 ( .A(prefillCounter), .SUM({N414, N413, N412, N411, 
        N410, N409, N408, N407}) );
  KSA_0_DW01_add_6 add_377 ( .A(temp), .B(extratemp), .CI(1'b0), .SUM({N527, 
        N526, N525, N524, N523, N522, N521, N520}) );
  KSA_0_DW01_add_7 add_337 ( .A(intj), .B(DATA_IN), .CI(1'b0), .SUM({N519, 
        N518, N517, N516, N515, N514, N513, N512}) );
  KSA_0_DW01_add_8 add_1_root_add_0_root_add_302_2 ( .A(DATA_IN), .B({sj[7:1], 
        n58}), .CI(1'b0), .SUM({N456, N455, N454, N453, N452, N451, N450, N449}) );
  KSA_0_DW01_add_9 add_0_root_add_0_root_add_302_2 ( .A({N472, N473, N474, 
        N475, N476, N477, N478, N479}), .B({N456, N455, N454, N453, N452, N451, 
        N450, N449}), .CI(1'b0), .SUM({N487, N486, N485, N484, N483, N482, 
        N481, N480}) );
  KSA_0_DW01_inc_3 r126 ( .A(inti), .SUM({N503, N502, N501, N500, N499, N498, 
        N497, N496}) );
  TBUFX1 \nfdata_tri[0]  ( .A(n1310), .EN(n77), .Y(nfdata[0]) );
  TBUFX1 \nfdata_tri[1]  ( .A(n1311), .EN(n77), .Y(nfdata[1]) );
  TBUFX1 \nfdata_tri[2]  ( .A(n1312), .EN(n77), .Y(nfdata[2]) );
  TBUFX1 \nfdata_tri[3]  ( .A(n1313), .EN(n77), .Y(nfdata[3]) );
  TBUFX1 \nfdata_tri[4]  ( .A(n1314), .EN(n77), .Y(nfdata[4]) );
  TBUFX1 \nfdata_tri[5]  ( .A(n1315), .EN(n77), .Y(nfdata[5]) );
  TBUFX1 \nfdata_tri[6]  ( .A(n1316), .EN(n77), .Y(nfdata[6]) );
  TBUFX1 \nfdata_tri[7]  ( .A(n1317), .EN(n77), .Y(nfdata[7]) );
  TBUFX1 \nfaddr_tri[4]  ( .A(n1306), .EN(n1099), .Y(nfaddr[4]) );
  TBUFX1 \nfaddr_tri[1]  ( .A(n1303), .EN(n1099), .Y(nfaddr[1]) );
  TBUFX1 \nfaddr_tri[2]  ( .A(n1304), .EN(n1099), .Y(nfaddr[2]) );
  TBUFX1 \nfaddr_tri[3]  ( .A(n1305), .EN(n1099), .Y(nfaddr[3]) );
  TBUFX1 \nfaddr_tri[0]  ( .A(n1302), .EN(n1099), .Y(nfaddr[0]) );
  TBUFX2 \nfaddr_tri[7]  ( .A(n1309), .EN(n1099), .Y(nfaddr[7]) );
  TBUFX1 \nfaddr_tri[6]  ( .A(n1308), .EN(n1099), .Y(nfaddr[6]) );
  TBUFX2 \nfaddr_tri[5]  ( .A(n1307), .EN(n1099), .Y(nfaddr[5]) );
  DFFSR \si_reg[7]  ( .D(n1153), .CLK(CLK), .R(n231), .S(1'b1), .Q(si[7]) );
  DFFSR \si_reg[3]  ( .D(n1149), .CLK(CLK), .R(n231), .S(1'b1), .Q(si[3]) );
  DFFSR \si_reg[2]  ( .D(n1148), .CLK(CLK), .R(n231), .S(1'b1), .Q(si[2]) );
  DFFSR \si_reg[5]  ( .D(n1151), .CLK(CLK), .R(n231), .S(1'b1), .Q(si[5]) );
  DFFSR \si_reg[4]  ( .D(n1150), .CLK(CLK), .R(n231), .S(1'b1), .Q(si[4]) );
  DFFSR \sj_reg[4]  ( .D(n1157), .CLK(CLK), .R(n231), .S(1'b1), .Q(sj[4]) );
  DFFSR \currentProcessedData_reg[6]  ( .D(nextProcessedData[6]), .CLK(CLK), 
        .R(n231), .S(1'b1), .Q(currentProcessedData[6]) );
  DFFSR \currentProcessedData_reg[4]  ( .D(nextProcessedData[4]), .CLK(CLK), 
        .R(n231), .S(1'b1), .Q(currentProcessedData[4]) );
  DFFSR \currentProcessedData_reg[1]  ( .D(nextProcessedData[1]), .CLK(CLK), 
        .R(n231), .S(1'b1), .Q(currentProcessedData[1]) );
  DFFSR \sj_reg[6]  ( .D(n1155), .CLK(CLK), .R(n231), .S(1'b1), .Q(sj[6]) );
  DFFSR \currentProcessedData_reg[7]  ( .D(nextProcessedData[7]), .CLK(CLK), 
        .R(n231), .S(1'b1), .Q(currentProcessedData[7]) );
  DFFSR \currentProcessedData_reg[5]  ( .D(nextProcessedData[5]), .CLK(CLK), 
        .R(n231), .S(1'b1), .Q(currentProcessedData[5]) );
  DFFSR \currentProcessedData_reg[3]  ( .D(nextProcessedData[3]), .CLK(CLK), 
        .R(n231), .S(1'b1), .Q(currentProcessedData[3]) );
  DFFSR \currentProcessedData_reg[2]  ( .D(nextProcessedData[2]), .CLK(CLK), 
        .R(n231), .S(1'b1), .Q(currentProcessedData[2]) );
  DFFSR \currentProcessedData_reg[0]  ( .D(nextProcessedData[0]), .CLK(CLK), 
        .R(n231), .S(1'b1), .Q(currentProcessedData[0]) );
  DFFSR \sj_reg[5]  ( .D(n1156), .CLK(CLK), .R(n231), .S(1'b1), .Q(sj[5]) );
  DFFSR \sj_reg[7]  ( .D(n1098), .CLK(CLK), .R(n231), .S(1'b1), .Q(sj[7]) );
  AND2X1 U3 ( .A(n1063), .B(n236), .Y(n3) );
  AND2X2 U4 ( .A(n175), .B(n144), .Y(n4) );
  INVX2 U7 ( .A(n701), .Y(n73) );
  AND2X2 U8 ( .A(n303), .B(n689), .Y(n5) );
  NAND2X1 U9 ( .A(n185), .B(n1088), .Y(n6) );
  AND2X2 U10 ( .A(n153), .B(n71), .Y(n7) );
  INVX1 U11 ( .A(n701), .Y(n452) );
  AND2X2 U12 ( .A(n1053), .B(n1051), .Y(n8) );
  INVX2 U13 ( .A(n225), .Y(n342) );
  INVX2 U14 ( .A(n265), .Y(n269) );
  OR2X1 U15 ( .A(n325), .B(n324), .Y(n9) );
  OR2X2 U16 ( .A(n361), .B(n360), .Y(n10) );
  NAND2X1 U17 ( .A(n33), .B(n36), .Y(n11) );
  AND2X1 U18 ( .A(n311), .B(n312), .Y(n12) );
  AND2X2 U19 ( .A(n65), .B(n68), .Y(n13) );
  NAND2X1 U37 ( .A(n153), .B(n71), .Y(n31) );
  INVX2 U38 ( .A(n214), .Y(n71) );
  BUFX4 U39 ( .A(n34), .Y(n32) );
  AND2X2 U40 ( .A(n208), .B(n144), .Y(n33) );
  NAND3X1 U41 ( .A(keyi[1]), .B(keyi[0]), .C(n520), .Y(n34) );
  INVX1 U42 ( .A(n169), .Y(n35) );
  BUFX4 U43 ( .A(n216), .Y(n169) );
  INVX2 U44 ( .A(n169), .Y(n117) );
  AND2X2 U45 ( .A(n213), .B(n299), .Y(n36) );
  INVX2 U46 ( .A(state[2]), .Y(n299) );
  NAND3X1 U47 ( .A(n54), .B(n267), .C(n84), .Y(n37) );
  INVX1 U48 ( .A(n171), .Y(n38) );
  NAND2X1 U49 ( .A(n214), .B(n299), .Y(n39) );
  XNOR2X1 U50 ( .A(n49), .B(n1069), .Y(n254) );
  NOR2X1 U51 ( .A(n229), .B(n1039), .Y(n40) );
  BUFX2 U52 ( .A(n486), .Y(n46) );
  INVX1 U53 ( .A(n215), .Y(n1087) );
  AND2X2 U54 ( .A(n149), .B(n252), .Y(n208) );
  INVX4 U55 ( .A(keyi[1]), .Y(n519) );
  INVX4 U56 ( .A(keyi[0]), .Y(n521) );
  INVX4 U57 ( .A(keyi[2]), .Y(n520) );
  BUFX4 U58 ( .A(n36), .Y(n41) );
  AND2X2 U59 ( .A(n229), .B(n244), .Y(n42) );
  INVX4 U60 ( .A(n83), .Y(n171) );
  INVX1 U61 ( .A(n420), .Y(n43) );
  INVX2 U62 ( .A(n43), .Y(n44) );
  BUFX4 U63 ( .A(n486), .Y(n45) );
  BUFX2 U64 ( .A(n175), .Y(n47) );
  INVX2 U65 ( .A(n299), .Y(n153) );
  BUFX2 U66 ( .A(n1063), .Y(n48) );
  BUFX4 U67 ( .A(state[4]), .Y(n49) );
  OAI21X1 U68 ( .A(n52), .B(n171), .C(n300), .Y(n50) );
  INVX1 U69 ( .A(n1073), .Y(n226) );
  INVX1 U70 ( .A(n66), .Y(n252) );
  BUFX2 U71 ( .A(n72), .Y(n51) );
  INVX2 U72 ( .A(n36), .Y(n52) );
  NAND2X1 U73 ( .A(n98), .B(n1020), .Y(n53) );
  INVX2 U74 ( .A(n97), .Y(n98) );
  NAND2X1 U75 ( .A(n40), .B(n41), .Y(n54) );
  INVX1 U76 ( .A(n178), .Y(n55) );
  INVX1 U77 ( .A(n55), .Y(n56) );
  INVX1 U78 ( .A(n692), .Y(n57) );
  BUFX2 U79 ( .A(state[1]), .Y(n149) );
  BUFX4 U80 ( .A(sj[0]), .Y(n58) );
  INVX1 U81 ( .A(n442), .Y(n1274) );
  INVX1 U82 ( .A(n441), .Y(n1275) );
  AND2X2 U83 ( .A(n639), .B(n59), .Y(n123) );
  NOR2X1 U84 ( .A(n180), .B(n166), .Y(n59) );
  AND2X2 U85 ( .A(n187), .B(n679), .Y(n60) );
  BUFX4 U86 ( .A(n1097), .Y(n61) );
  BUFX4 U87 ( .A(n1097), .Y(n62) );
  AND2X2 U88 ( .A(n210), .B(n1057), .Y(n147) );
  INVX1 U89 ( .A(n216), .Y(n656) );
  INVX2 U90 ( .A(n1053), .Y(n63) );
  INVX1 U91 ( .A(n60), .Y(n64) );
  INVX1 U92 ( .A(n64), .Y(n65) );
  INVX2 U93 ( .A(n211), .Y(n66) );
  INVX1 U94 ( .A(n211), .Y(n212) );
  NAND2X1 U95 ( .A(n154), .B(n41), .Y(n67) );
  NAND2X1 U96 ( .A(n154), .B(n41), .Y(n68) );
  INVX1 U97 ( .A(n310), .Y(n99) );
  BUFX2 U98 ( .A(n196), .Y(n69) );
  NOR2X1 U99 ( .A(n638), .B(n180), .Y(n70) );
  INVX2 U100 ( .A(n67), .Y(n89) );
  AND2X2 U101 ( .A(n271), .B(n270), .Y(n187) );
  INVX1 U102 ( .A(n458), .Y(n489) );
  INVX2 U103 ( .A(n39), .Y(n72) );
  INVX4 U104 ( .A(n86), .Y(n616) );
  INVX2 U105 ( .A(n211), .Y(n74) );
  INVX1 U106 ( .A(n54), .Y(n1053) );
  AND2X2 U107 ( .A(n271), .B(n270), .Y(n75) );
  BUFX4 U108 ( .A(n683), .Y(n76) );
  INVX1 U109 ( .A(n683), .Y(n228) );
  INVX2 U112 ( .A(n1061), .Y(n77) );
  INVX1 U113 ( .A(n171), .Y(n78) );
  NOR2X1 U114 ( .A(n364), .B(si[3]), .Y(n79) );
  INVX1 U115 ( .A(n79), .Y(n349) );
  NAND2X1 U116 ( .A(n109), .B(n314), .Y(n80) );
  NOR2X1 U117 ( .A(n80), .B(n81), .Y(n182) );
  OR2X2 U118 ( .A(n82), .B(n497), .Y(n81) );
  INVX1 U119 ( .A(n68), .Y(n82) );
  INVX2 U120 ( .A(n214), .Y(n1069) );
  AND2X2 U121 ( .A(n49), .B(n196), .Y(n83) );
  AND2X2 U122 ( .A(n210), .B(n1057), .Y(n84) );
  INVX1 U124 ( .A(n214), .Y(n164) );
  NOR2X1 U125 ( .A(n215), .B(n262), .Y(n85) );
  NOR2X1 U127 ( .A(n359), .B(n10), .Y(n1305) );
  MUX2X1 U128 ( .B(faddr[6]), .A(nfaddr[6]), .S(n237), .Y(n448) );
  AND2X2 U129 ( .A(n253), .B(n617), .Y(n86) );
  BUFX2 U134 ( .A(n221), .Y(n87) );
  INVX2 U135 ( .A(n157), .Y(n179) );
  INVX1 U136 ( .A(n118), .Y(n88) );
  NAND2X1 U137 ( .A(n11), .B(n3), .Y(n690) );
  MUX2X1 U138 ( .B(ADDR[6]), .A(nfaddr[6]), .S(n238), .Y(n447) );
  NAND2X1 U139 ( .A(n185), .B(n1088), .Y(n90) );
  INVX2 U140 ( .A(n104), .Y(n1094) );
  INVX1 U141 ( .A(n228), .Y(n91) );
  AND2X2 U144 ( .A(n79), .B(n1103), .Y(n92) );
  INVX1 U145 ( .A(n92), .Y(n330) );
  INVX1 U146 ( .A(n445), .Y(n1271) );
  INVX8 U147 ( .A(n76), .Y(n93) );
  INVX1 U148 ( .A(n448), .Y(n1268) );
  INVX1 U149 ( .A(n179), .Y(n94) );
  INVX1 U150 ( .A(n447), .Y(n1269) );
  AND2X2 U151 ( .A(n13), .B(n221), .Y(n223) );
  INVX1 U152 ( .A(n1020), .Y(n95) );
  INVX1 U153 ( .A(n95), .Y(n96) );
  NAND2X1 U154 ( .A(n150), .B(n60), .Y(n97) );
  NAND2X1 U155 ( .A(n98), .B(n1020), .Y(n773) );
  INVX1 U157 ( .A(n657), .Y(n496) );
  AND2X2 U161 ( .A(n100), .B(n99), .Y(n311) );
  NAND2X1 U162 ( .A(n656), .B(faddr[7]), .Y(n100) );
  NAND2X1 U163 ( .A(n109), .B(n314), .Y(n101) );
  INVX1 U164 ( .A(n151), .Y(n102) );
  NAND2X1 U165 ( .A(n679), .B(n75), .Y(n103) );
  AND2X2 U166 ( .A(n746), .B(n87), .Y(n104) );
  INVX1 U167 ( .A(n75), .Y(n105) );
  INVX1 U168 ( .A(n105), .Y(n106) );
  INVX1 U169 ( .A(n5), .Y(n225) );
  NOR2X1 U170 ( .A(n188), .B(n108), .Y(n107) );
  NAND2X1 U171 ( .A(n303), .B(n305), .Y(n108) );
  INVX1 U172 ( .A(n11), .Y(n1061) );
  BUFX2 U173 ( .A(n185), .Y(n109) );
  INVX1 U174 ( .A(si[0]), .Y(n1101) );
  BUFX2 U175 ( .A(n225), .Y(n110) );
  INVX2 U176 ( .A(n1076), .Y(n111) );
  INVX1 U177 ( .A(n182), .Y(n112) );
  INVX1 U178 ( .A(n112), .Y(n113) );
  AND2X2 U179 ( .A(n7), .B(n175), .Y(n114) );
  AND2X1 U180 ( .A(n7), .B(n208), .Y(n219) );
  INVX1 U181 ( .A(n228), .Y(n115) );
  INVX1 U182 ( .A(n153), .Y(n116) );
  NOR2X1 U183 ( .A(n118), .B(n119), .Y(n120) );
  NOR2X1 U184 ( .A(n120), .B(n103), .Y(n314) );
  INVX1 U185 ( .A(n33), .Y(n118) );
  INVX1 U186 ( .A(n164), .Y(n119) );
  BUFX2 U187 ( .A(n222), .Y(n121) );
  INVX1 U188 ( .A(n1039), .Y(n1040) );
  INVX1 U189 ( .A(n53), .Y(n746) );
  NOR2X1 U190 ( .A(n326), .B(n9), .Y(n1308) );
  AND2X2 U191 ( .A(n491), .B(n490), .Y(n122) );
  INVX1 U192 ( .A(n122), .Y(nextProcessedData[0]) );
  AND2X2 U193 ( .A(n12), .B(n313), .Y(n1309) );
  INVX1 U194 ( .A(n123), .Y(n1054) );
  AND2X2 U195 ( .A(n484), .B(n483), .Y(n125) );
  INVX1 U196 ( .A(n125), .Y(nextProcessedData[1]) );
  AND2X2 U197 ( .A(n480), .B(n479), .Y(n127) );
  INVX1 U198 ( .A(n127), .Y(nextProcessedData[2]) );
  AND2X2 U199 ( .A(n476), .B(n475), .Y(n129) );
  INVX1 U200 ( .A(n129), .Y(nextProcessedData[3]) );
  AND2X2 U201 ( .A(n472), .B(n471), .Y(n131) );
  INVX1 U202 ( .A(n131), .Y(nextProcessedData[4]) );
  AND2X2 U203 ( .A(n468), .B(n467), .Y(n132) );
  INVX1 U204 ( .A(n132), .Y(nextProcessedData[5]) );
  AND2X2 U205 ( .A(n464), .B(n463), .Y(n133) );
  INVX1 U206 ( .A(n133), .Y(nextProcessedData[6]) );
  AND2X2 U207 ( .A(n460), .B(n459), .Y(n134) );
  INVX1 U208 ( .A(n134), .Y(nextProcessedData[7]) );
  AND2X2 U209 ( .A(n1068), .B(n206), .Y(n135) );
  INVX1 U210 ( .A(n135), .Y(n596) );
  INVX1 U211 ( .A(n92), .Y(n136) );
  INVX1 U212 ( .A(n136), .Y(n137) );
  BUFX4 U213 ( .A(n184), .Y(n138) );
  BUFX4 U214 ( .A(n184), .Y(n139) );
  BUFX4 U215 ( .A(n184), .Y(n140) );
  BUFX4 U216 ( .A(n184), .Y(n141) );
  BUFX4 U217 ( .A(n184), .Y(n142) );
  BUFX4 U218 ( .A(n184), .Y(n143) );
  INVX2 U219 ( .A(n49), .Y(n144) );
  INVX1 U220 ( .A(n434), .Y(n1282) );
  INVX1 U221 ( .A(n433), .Y(n1283) );
  INVX1 U222 ( .A(n431), .Y(n1285) );
  INVX1 U223 ( .A(n430), .Y(n1286) );
  INVX1 U224 ( .A(n429), .Y(n1287) );
  INVX1 U225 ( .A(n428), .Y(n1288) );
  INVX1 U226 ( .A(n427), .Y(n1289) );
  INVX1 U227 ( .A(n410), .Y(n1294) );
  INVX1 U228 ( .A(n409), .Y(n1295) );
  INVX1 U229 ( .A(n407), .Y(n1297) );
  INVX1 U230 ( .A(n406), .Y(n1298) );
  INVX1 U231 ( .A(n405), .Y(n1299) );
  INVX1 U232 ( .A(n404), .Y(n1300) );
  INVX1 U233 ( .A(n403), .Y(n1301) );
  INVX1 U234 ( .A(n229), .Y(n145) );
  NOR2X1 U235 ( .A(n229), .B(n1039), .Y(n189) );
  BUFX2 U236 ( .A(n329), .Y(n146) );
  INVX1 U237 ( .A(n84), .Y(n1046) );
  AND2X2 U238 ( .A(n329), .B(n302), .Y(n148) );
  AND2X1 U239 ( .A(n146), .B(n302), .Y(n199) );
  BUFX2 U240 ( .A(state[1]), .Y(n230) );
  BUFX2 U241 ( .A(n701), .Y(n150) );
  INVX1 U242 ( .A(n450), .Y(n1266) );
  INVX1 U243 ( .A(n449), .Y(n1267) );
  INVX1 U244 ( .A(n160), .Y(n151) );
  NOR2X1 U245 ( .A(n229), .B(n152), .Y(n160) );
  NAND2X1 U246 ( .A(n74), .B(n243), .Y(n152) );
  INVX2 U247 ( .A(n230), .Y(n243) );
  AND2X2 U248 ( .A(n212), .B(n243), .Y(n196) );
  BUFX2 U249 ( .A(n190), .Y(n154) );
  AND2X2 U250 ( .A(n259), .B(n74), .Y(n156) );
  AND2X2 U251 ( .A(n451), .B(n458), .Y(n157) );
  INVX1 U252 ( .A(n94), .Y(n1134) );
  INVX1 U253 ( .A(n270), .Y(n1042) );
  INVX1 U254 ( .A(n156), .Y(n263) );
  BUFX2 U255 ( .A(n493), .Y(n161) );
  NAND3X1 U256 ( .A(n54), .B(n267), .C(n84), .Y(n162) );
  NAND2X1 U257 ( .A(n121), .B(n1072), .Y(n166) );
  INVX1 U258 ( .A(n101), .Y(n1099) );
  BUFX2 U259 ( .A(n114), .Y(n167) );
  NAND2X1 U260 ( .A(n85), .B(n107), .Y(n420) );
  INVX4 U261 ( .A(n188), .Y(n222) );
  AND2X2 U262 ( .A(n153), .B(n214), .Y(n192) );
  INVX2 U263 ( .A(n590), .Y(n170) );
  NOR2X1 U264 ( .A(n172), .B(n162), .Y(n216) );
  NAND2X1 U265 ( .A(n157), .B(n67), .Y(n172) );
  AND2X2 U266 ( .A(n149), .B(n252), .Y(n175) );
  INVX2 U267 ( .A(n253), .Y(n177) );
  INVX4 U268 ( .A(n223), .Y(n224) );
  NOR2X1 U269 ( .A(n1061), .B(n655), .Y(n660) );
  AND2X1 U270 ( .A(n96), .B(n1019), .Y(n181) );
  OR2X1 U271 ( .A(n568), .B(n569), .Y(n183) );
  AND2X1 U272 ( .A(keyi[2]), .B(keyi[1]), .Y(n200) );
  INVX2 U273 ( .A(n237), .Y(n234) );
  INVX2 U274 ( .A(n238), .Y(n233) );
  INVX2 U275 ( .A(n236), .Y(n235) );
  INVX2 U276 ( .A(n654), .Y(n1018) );
  BUFX2 U277 ( .A(n613), .Y(n201) );
  NOR2X1 U278 ( .A(n179), .B(n455), .Y(n178) );
  BUFX2 U279 ( .A(n231), .Y(n236) );
  BUFX2 U280 ( .A(n231), .Y(n237) );
  BUFX2 U281 ( .A(n231), .Y(n238) );
  BUFX2 U282 ( .A(n236), .Y(n239) );
  BUFX2 U283 ( .A(n237), .Y(n240) );
  BUFX2 U284 ( .A(n238), .Y(n241) );
  BUFX2 U285 ( .A(n231), .Y(n242) );
  OR2X2 U286 ( .A(n101), .B(n232), .Y(n180) );
  AND2X2 U287 ( .A(n221), .B(n774), .Y(n184) );
  AND2X2 U288 ( .A(n135), .B(n1044), .Y(n185) );
  AND2X2 U289 ( .A(n192), .B(n156), .Y(n188) );
  AND2X2 U290 ( .A(n197), .B(n144), .Y(n190) );
  INVX2 U291 ( .A(RST), .Y(n231) );
  AND2X2 U292 ( .A(n200), .B(n521), .Y(n191) );
  MUX2X1 U293 ( .B(n1101), .A(n521), .S(n193), .Y(n1172) );
  NAND2X1 U294 ( .A(n123), .B(n68), .Y(n193) );
  MUX2X1 U295 ( .B(n1102), .A(n519), .S(n194), .Y(n1171) );
  NAND2X1 U296 ( .A(n123), .B(n68), .Y(n194) );
  MUX2X1 U297 ( .B(n650), .A(n520), .S(n195), .Y(n1170) );
  NAND2X1 U298 ( .A(n123), .B(n68), .Y(n195) );
  NOR2X1 U299 ( .A(n149), .B(n212), .Y(n197) );
  AND2X2 U300 ( .A(n200), .B(keyi[0]), .Y(n198) );
  INVX1 U301 ( .A(n638), .Y(n639) );
  INVX1 U302 ( .A(n1057), .Y(n1082) );
  NAND2X1 U303 ( .A(n272), .B(n78), .Y(n202) );
  INVX1 U304 ( .A(n689), .Y(n294) );
  BUFX2 U305 ( .A(n1068), .Y(n203) );
  NAND2X1 U306 ( .A(n205), .B(n269), .Y(n206) );
  INVX1 U307 ( .A(n31), .Y(n205) );
  NAND2X1 U308 ( .A(n244), .B(n229), .Y(n207) );
  BUFX2 U309 ( .A(n149), .Y(n209) );
  INVX1 U310 ( .A(n227), .Y(n1074) );
  INVX4 U311 ( .A(n226), .Y(n227) );
  AND2X2 U312 ( .A(n1072), .B(n493), .Y(n210) );
  INVX1 U313 ( .A(n210), .Y(n1083) );
  INVX2 U314 ( .A(state[0]), .Y(n211) );
  INVX2 U315 ( .A(state[3]), .Y(n213) );
  INVX4 U316 ( .A(n213), .Y(n214) );
  AND2X2 U317 ( .A(n219), .B(n49), .Y(n215) );
  BUFX4 U318 ( .A(state[4]), .Y(n229) );
  AND2X1 U319 ( .A(n1087), .B(n150), .Y(n255) );
  INVX1 U320 ( .A(n114), .Y(n340) );
  INVX1 U321 ( .A(n1044), .Y(n253) );
  AND2X2 U322 ( .A(n617), .B(n111), .Y(n217) );
  AND2X2 U323 ( .A(n617), .B(n111), .Y(n218) );
  OR2X2 U324 ( .A(n1080), .B(n207), .Y(n1063) );
  INVX1 U325 ( .A(n31), .Y(n272) );
  INVX1 U326 ( .A(n1072), .Y(n1076) );
  INVX1 U327 ( .A(n1088), .Y(n590) );
  INVX1 U328 ( .A(n1080), .Y(n1041) );
  NAND2X1 U329 ( .A(n181), .B(n223), .Y(n1021) );
  NOR2X1 U330 ( .A(n657), .B(n183), .Y(n574) );
  INVX1 U331 ( .A(n689), .Y(n692) );
  NOR2X1 U332 ( .A(n638), .B(n180), .Y(n516) );
  BUFX2 U333 ( .A(n657), .Y(n220) );
  INVX2 U334 ( .A(n242), .Y(n232) );
  AND2X2 U335 ( .A(n178), .B(n268), .Y(n221) );
  INVX1 U336 ( .A(n87), .Y(n423) );
  INVX1 U337 ( .A(n1063), .Y(n295) );
  INVX4 U338 ( .A(n1021), .Y(n1036) );
  INVX8 U339 ( .A(n76), .Y(n684) );
  INVX2 U340 ( .A(si[1]), .Y(n1102) );
  INVX2 U341 ( .A(si[4]), .Y(n1103) );
  INVX2 U342 ( .A(si[5]), .Y(n1104) );
  INVX2 U343 ( .A(prefillCounter[5]), .Y(n1135) );
  NAND3X1 U344 ( .A(n197), .B(n145), .C(n192), .Y(n1072) );
  NOR2X1 U345 ( .A(n230), .B(n66), .Y(n244) );
  NAND2X1 U346 ( .A(n42), .B(n192), .Y(n493) );
  INVX2 U347 ( .A(n1329), .Y(n245) );
  NAND2X1 U348 ( .A(n1083), .B(n245), .Y(n250) );
  NAND2X1 U349 ( .A(n49), .B(n196), .Y(n264) );
  NAND2X1 U350 ( .A(n78), .B(n245), .Y(n247) );
  NAND3X1 U351 ( .A(n149), .B(n74), .C(n229), .Y(n265) );
  OAI21X1 U352 ( .A(n1328), .B(n1106), .C(n269), .Y(n246) );
  NAND2X1 U353 ( .A(n247), .B(n246), .Y(n248) );
  NAND2X1 U354 ( .A(n51), .B(n248), .Y(n249) );
  NAND2X1 U355 ( .A(n250), .B(n249), .Y(n251) );
  AOI22X1 U356 ( .A(n69), .B(n41), .C(n1105), .D(n251), .Y(n1327) );
  NAND2X1 U357 ( .A(n114), .B(n145), .Y(n1088) );
  NAND2X1 U358 ( .A(n149), .B(n74), .Y(n1039) );
  NAND2X1 U359 ( .A(n189), .B(n72), .Y(n270) );
  INVX2 U360 ( .A(permuteComplete), .Y(n1050) );
  NAND2X1 U361 ( .A(n192), .B(n33), .Y(n1044) );
  AOI21X1 U362 ( .A(n1042), .B(n1050), .C(n253), .Y(n256) );
  NAND3X1 U363 ( .A(n254), .B(n175), .C(n116), .Y(n701) );
  NAND3X1 U364 ( .A(n1088), .B(n256), .C(n255), .Y(n1065) );
  INVX2 U365 ( .A(n1065), .Y(n1100) );
  NOR2X1 U366 ( .A(prefillCounter[0]), .B(n1325), .Y(n257) );
  NAND3X1 U367 ( .A(n1324), .B(n1061), .C(n257), .Y(n258) );
  NAND3X1 U368 ( .A(n72), .B(n175), .C(n49), .Y(n458) );
  NAND2X1 U369 ( .A(n258), .B(n458), .Y(n261) );
  NAND2X1 U370 ( .A(n83), .B(n7), .Y(n679) );
  NOR2X1 U371 ( .A(n229), .B(n149), .Y(n259) );
  NAND2X1 U372 ( .A(n202), .B(n263), .Y(n260) );
  NOR2X1 U373 ( .A(n261), .B(n260), .Y(n1326) );
  NAND2X1 U374 ( .A(n42), .B(n72), .Y(n451) );
  NAND2X1 U375 ( .A(n42), .B(n36), .Y(n1068) );
  NAND2X1 U376 ( .A(n153), .B(n1069), .Y(n1080) );
  NAND2X1 U377 ( .A(n189), .B(n7), .Y(n300) );
  OAI21X1 U378 ( .A(n52), .B(n171), .C(n300), .Y(n262) );
  NOR2X1 U379 ( .A(n215), .B(n50), .Y(n454) );
  NAND2X1 U380 ( .A(n190), .B(n272), .Y(n303) );
  NAND2X1 U381 ( .A(n40), .B(n192), .Y(n305) );
  NOR2X1 U382 ( .A(n90), .B(n420), .Y(n268) );
  NAND2X1 U383 ( .A(n40), .B(n36), .Y(n634) );
  NAND2X1 U384 ( .A(n102), .B(n272), .Y(n267) );
  NAND2X1 U385 ( .A(n265), .B(n264), .Y(n266) );
  NAND2X1 U386 ( .A(n72), .B(n266), .Y(n1057) );
  NAND3X1 U387 ( .A(n634), .B(n267), .C(n147), .Y(n455) );
  AOI22X1 U388 ( .A(n160), .B(n72), .C(n269), .D(n36), .Y(n271) );
  NAND2X1 U389 ( .A(n679), .B(n187), .Y(n569) );
  NAND2X1 U390 ( .A(n190), .B(n72), .Y(n689) );
  NAND2X1 U391 ( .A(n294), .B(DATA_IN[7]), .Y(n274) );
  NAND2X1 U392 ( .A(n36), .B(n156), .Y(n654) );
  NAND2X1 U393 ( .A(prefillCounter[7]), .B(n1018), .Y(n309) );
  AOI22X1 U394 ( .A(extratemp[7]), .B(n295), .C(n73), .D(temp[7]), .Y(n273) );
  NAND3X1 U395 ( .A(n274), .B(n309), .C(n273), .Y(n275) );
  AOI21X1 U396 ( .A(fdata[7]), .B(n224), .C(n275), .Y(n1317) );
  NAND2X1 U397 ( .A(n294), .B(DATA_IN[6]), .Y(n277) );
  NAND2X1 U398 ( .A(prefillCounter[6]), .B(n1018), .Y(n320) );
  AOI22X1 U399 ( .A(extratemp[6]), .B(n295), .C(n73), .D(temp[6]), .Y(n276) );
  NAND3X1 U400 ( .A(n277), .B(n320), .C(n276), .Y(n278) );
  AOI21X1 U401 ( .A(fdata[6]), .B(n224), .C(n278), .Y(n1316) );
  NAND2X1 U402 ( .A(n294), .B(DATA_IN[5]), .Y(n280) );
  NAND2X1 U403 ( .A(n1018), .B(prefillCounter[5]), .Y(n327) );
  AOI22X1 U404 ( .A(extratemp[5]), .B(n295), .C(n73), .D(temp[5]), .Y(n279) );
  NAND3X1 U405 ( .A(n280), .B(n327), .C(n279), .Y(n281) );
  AOI21X1 U406 ( .A(n224), .B(fdata[5]), .C(n281), .Y(n1315) );
  NAND2X1 U407 ( .A(n294), .B(DATA_IN[4]), .Y(n283) );
  NAND2X1 U408 ( .A(prefillCounter[4]), .B(n1018), .Y(n338) );
  AOI22X1 U409 ( .A(extratemp[4]), .B(n295), .C(n73), .D(temp[4]), .Y(n282) );
  NAND3X1 U410 ( .A(n283), .B(n338), .C(n282), .Y(n284) );
  AOI21X1 U411 ( .A(fdata[4]), .B(n224), .C(n284), .Y(n1314) );
  NAND2X1 U412 ( .A(n294), .B(DATA_IN[3]), .Y(n286) );
  NAND2X1 U413 ( .A(prefillCounter[3]), .B(n1018), .Y(n355) );
  AOI22X1 U414 ( .A(extratemp[3]), .B(n295), .C(n73), .D(temp[3]), .Y(n285) );
  NAND3X1 U415 ( .A(n286), .B(n355), .C(n285), .Y(n287) );
  AOI21X1 U416 ( .A(fdata[3]), .B(n224), .C(n287), .Y(n1313) );
  NAND2X1 U417 ( .A(n294), .B(DATA_IN[2]), .Y(n289) );
  NAND2X1 U418 ( .A(prefillCounter[2]), .B(n1018), .Y(n369) );
  AOI22X1 U419 ( .A(extratemp[2]), .B(n295), .C(n73), .D(temp[2]), .Y(n288) );
  NAND3X1 U420 ( .A(n289), .B(n369), .C(n288), .Y(n290) );
  AOI21X1 U421 ( .A(fdata[2]), .B(n224), .C(n290), .Y(n1312) );
  NAND2X1 U422 ( .A(n294), .B(DATA_IN[1]), .Y(n292) );
  NAND2X1 U423 ( .A(prefillCounter[1]), .B(n1018), .Y(n383) );
  AOI22X1 U424 ( .A(extratemp[1]), .B(n295), .C(n73), .D(temp[1]), .Y(n291) );
  NAND3X1 U425 ( .A(n292), .B(n383), .C(n291), .Y(n293) );
  AOI21X1 U426 ( .A(fdata[1]), .B(n224), .C(n293), .Y(n1311) );
  NAND2X1 U427 ( .A(n294), .B(DATA_IN[0]), .Y(n297) );
  NAND2X1 U428 ( .A(prefillCounter[0]), .B(n1018), .Y(n395) );
  AOI22X1 U429 ( .A(extratemp[0]), .B(n295), .C(n73), .D(temp[0]), .Y(n296) );
  NAND3X1 U430 ( .A(n297), .B(n395), .C(n296), .Y(n298) );
  AOI21X1 U431 ( .A(n224), .B(fdata[0]), .C(n298), .Y(n1310) );
  NAND2X1 U432 ( .A(n4), .B(n116), .Y(n411) );
  NAND2X1 U433 ( .A(n411), .B(n300), .Y(n390) );
  OR2X2 U434 ( .A(si[1]), .B(si[0]), .Y(n378) );
  INVX2 U435 ( .A(n378), .Y(n301) );
  INVX2 U436 ( .A(si[2]), .Y(n650) );
  NAND2X1 U437 ( .A(n301), .B(n650), .Y(n364) );
  INVX2 U438 ( .A(si[3]), .Y(n648) );
  NAND2X1 U439 ( .A(n92), .B(n1104), .Y(n315) );
  INVX2 U440 ( .A(n315), .Y(n329) );
  INVX2 U441 ( .A(si[6]), .Y(n302) );
  XOR2X1 U442 ( .A(n148), .B(si[7]), .Y(n304) );
  AOI22X1 U443 ( .A(sj[7]), .B(n390), .C(n304), .D(n110), .Y(n313) );
  INVX2 U444 ( .A(n222), .Y(n497) );
  NAND2X1 U445 ( .A(n305), .B(n1063), .Y(n1073) );
  AOI22X1 U446 ( .A(N503), .B(n497), .C(intj[7]), .D(n227), .Y(n312) );
  NAND2X1 U447 ( .A(temp[7]), .B(n167), .Y(n308) );
  OAI21X1 U448 ( .A(n47), .B(n38), .C(n41), .Y(n306) );
  INVX2 U449 ( .A(n306), .Y(n397) );
  NAND2X1 U450 ( .A(n397), .B(inti[7]), .Y(n307) );
  NAND3X1 U451 ( .A(n309), .B(n308), .C(n307), .Y(n310) );
  NAND2X1 U452 ( .A(sj[6]), .B(n390), .Y(n319) );
  AND2X2 U453 ( .A(si[6]), .B(n315), .Y(n316) );
  OAI21X1 U454 ( .A(n199), .B(n316), .C(n110), .Y(n318) );
  AOI22X1 U455 ( .A(intj[6]), .B(n227), .C(N502), .D(n497), .Y(n317) );
  NAND3X1 U456 ( .A(n319), .B(n318), .C(n317), .Y(n326) );
  NAND2X1 U457 ( .A(temp[6]), .B(n167), .Y(n321) );
  NAND2X1 U458 ( .A(n321), .B(n320), .Y(n325) );
  INVX2 U459 ( .A(faddr[6]), .Y(n323) );
  NAND2X1 U460 ( .A(n397), .B(inti[6]), .Y(n322) );
  OAI21X1 U461 ( .A(n169), .B(n323), .C(n322), .Y(n324) );
  INVX2 U462 ( .A(temp[5]), .Y(n328) );
  OAI21X1 U463 ( .A(n340), .B(n328), .C(n327), .Y(n335) );
  AND2X2 U464 ( .A(sj[5]), .B(n390), .Y(n334) );
  AOI21X1 U465 ( .A(n330), .B(si[5]), .C(n146), .Y(n332) );
  AOI22X1 U466 ( .A(N501), .B(n497), .C(intj[5]), .D(n227), .Y(n331) );
  OAI21X1 U467 ( .A(n332), .B(n342), .C(n331), .Y(n333) );
  NOR3X1 U468 ( .A(n335), .B(n334), .C(n333), .Y(n337) );
  AOI22X1 U469 ( .A(n117), .B(faddr[5]), .C(n397), .D(inti[5]), .Y(n336) );
  AND2X2 U470 ( .A(n337), .B(n336), .Y(n1307) );
  INVX2 U471 ( .A(temp[4]), .Y(n339) );
  OAI21X1 U472 ( .A(n340), .B(n339), .C(n338), .Y(n346) );
  AND2X2 U473 ( .A(sj[4]), .B(n390), .Y(n345) );
  AOI21X1 U474 ( .A(n349), .B(si[4]), .C(n137), .Y(n343) );
  AOI22X1 U475 ( .A(N500), .B(n497), .C(intj[4]), .D(n227), .Y(n341) );
  OAI21X1 U476 ( .A(n343), .B(n342), .C(n341), .Y(n344) );
  NOR3X1 U477 ( .A(n346), .B(n345), .C(n344), .Y(n348) );
  AOI22X1 U478 ( .A(faddr[4]), .B(n117), .C(n397), .D(inti[4]), .Y(n347) );
  AND2X2 U479 ( .A(n348), .B(n347), .Y(n1306) );
  NAND2X1 U480 ( .A(sj[3]), .B(n390), .Y(n354) );
  NAND2X1 U481 ( .A(si[3]), .B(n364), .Y(n350) );
  NAND2X1 U482 ( .A(n350), .B(n349), .Y(n351) );
  NAND2X1 U483 ( .A(n351), .B(n225), .Y(n353) );
  AOI22X1 U484 ( .A(intj[3]), .B(n227), .C(N499), .D(n497), .Y(n352) );
  NAND3X1 U485 ( .A(n354), .B(n353), .C(n352), .Y(n361) );
  NAND2X1 U486 ( .A(temp[3]), .B(n167), .Y(n356) );
  NAND2X1 U487 ( .A(n356), .B(n355), .Y(n360) );
  INVX2 U488 ( .A(faddr[3]), .Y(n358) );
  NAND2X1 U489 ( .A(n397), .B(inti[3]), .Y(n357) );
  OAI21X1 U490 ( .A(n169), .B(n358), .C(n357), .Y(n359) );
  NAND2X1 U491 ( .A(n397), .B(inti[2]), .Y(n363) );
  NAND2X1 U492 ( .A(faddr[2]), .B(n35), .Y(n362) );
  NAND2X1 U493 ( .A(n363), .B(n362), .Y(n375) );
  NAND2X1 U494 ( .A(si[2]), .B(n378), .Y(n365) );
  NAND2X1 U495 ( .A(n365), .B(n364), .Y(n368) );
  INVX2 U496 ( .A(N498), .Y(n507) );
  NAND2X1 U497 ( .A(intj[2]), .B(n227), .Y(n366) );
  OAI21X1 U498 ( .A(n121), .B(n507), .C(n366), .Y(n367) );
  AOI21X1 U499 ( .A(n368), .B(n110), .C(n367), .Y(n373) );
  NAND2X1 U500 ( .A(sj[2]), .B(n390), .Y(n372) );
  INVX2 U501 ( .A(n369), .Y(n370) );
  AOI21X1 U502 ( .A(temp[2]), .B(n167), .C(n370), .Y(n371) );
  NAND3X1 U503 ( .A(n373), .B(n372), .C(n371), .Y(n374) );
  NOR2X1 U504 ( .A(n375), .B(n374), .Y(n1304) );
  NAND2X1 U505 ( .A(n397), .B(inti[1]), .Y(n377) );
  NAND2X1 U506 ( .A(faddr[1]), .B(n117), .Y(n376) );
  NAND2X1 U507 ( .A(n377), .B(n376), .Y(n389) );
  NAND2X1 U508 ( .A(si[0]), .B(si[1]), .Y(n379) );
  NAND2X1 U509 ( .A(n379), .B(n378), .Y(n382) );
  INVX2 U510 ( .A(N497), .Y(n509) );
  NAND2X1 U511 ( .A(intj[1]), .B(n227), .Y(n380) );
  OAI21X1 U512 ( .A(n121), .B(n509), .C(n380), .Y(n381) );
  AOI21X1 U513 ( .A(n382), .B(n110), .C(n381), .Y(n387) );
  NAND2X1 U514 ( .A(sj[1]), .B(n390), .Y(n386) );
  INVX2 U515 ( .A(n383), .Y(n384) );
  AOI21X1 U516 ( .A(temp[1]), .B(n167), .C(n384), .Y(n385) );
  NAND3X1 U517 ( .A(n387), .B(n386), .C(n385), .Y(n388) );
  NOR2X1 U518 ( .A(n389), .B(n388), .Y(n1303) );
  NAND2X1 U519 ( .A(n58), .B(n390), .Y(n394) );
  NAND2X1 U520 ( .A(n225), .B(n1101), .Y(n393) );
  INVX2 U521 ( .A(N496), .Y(n511) );
  NOR2X1 U522 ( .A(n222), .B(n511), .Y(n391) );
  AOI21X1 U523 ( .A(intj[0]), .B(n227), .C(n391), .Y(n392) );
  NAND3X1 U524 ( .A(n394), .B(n393), .C(n392), .Y(n402) );
  NAND2X1 U525 ( .A(temp[0]), .B(n167), .Y(n396) );
  NAND2X1 U526 ( .A(n396), .B(n395), .Y(n401) );
  INVX2 U527 ( .A(faddr[0]), .Y(n399) );
  NAND2X1 U528 ( .A(n397), .B(inti[0]), .Y(n398) );
  OAI21X1 U529 ( .A(n169), .B(n399), .C(n398), .Y(n400) );
  NOR3X1 U530 ( .A(n402), .B(n401), .C(n400), .Y(n1302) );
  MUX2X1 U531 ( .B(nfdata[0]), .A(DATA[0]), .S(n232), .Y(n403) );
  MUX2X1 U532 ( .B(nfdata[1]), .A(DATA[1]), .S(n234), .Y(n404) );
  MUX2X1 U533 ( .B(nfdata[2]), .A(DATA[2]), .S(n235), .Y(n405) );
  MUX2X1 U534 ( .B(nfdata[3]), .A(DATA[3]), .S(n235), .Y(n406) );
  MUX2X1 U535 ( .B(nfdata[4]), .A(DATA[4]), .S(n235), .Y(n407) );
  MUX2X1 U536 ( .B(nfdata[5]), .A(DATA[5]), .S(n235), .Y(n408) );
  INVX2 U537 ( .A(n408), .Y(n1296) );
  MUX2X1 U538 ( .B(nfdata[6]), .A(DATA[6]), .S(n234), .Y(n409) );
  MUX2X1 U539 ( .B(nfdata[7]), .A(DATA[7]), .S(n234), .Y(n410) );
  NOR2X1 U540 ( .A(n1018), .B(n103), .Y(n413) );
  AND2X2 U541 ( .A(n411), .B(n48), .Y(n412) );
  NAND3X1 U542 ( .A(n413), .B(n56), .C(n412), .Y(n419) );
  AOI21X1 U543 ( .A(fr_enable), .B(n419), .C(n44), .Y(n415) );
  INVX2 U544 ( .A(R_ENABLE), .Y(n414) );
  MUX2X1 U545 ( .B(n415), .A(n414), .S(n234), .Y(n1293) );
  AND2X2 U546 ( .A(n150), .B(n654), .Y(n416) );
  NAND3X1 U547 ( .A(n57), .B(n48), .C(n416), .Y(n424) );
  AOI21X1 U548 ( .A(fw_enable), .B(n423), .C(n424), .Y(n418) );
  INVX2 U549 ( .A(W_ENABLE), .Y(n417) );
  MUX2X1 U550 ( .B(n418), .A(n417), .S(n234), .Y(n1292) );
  OAI21X1 U551 ( .A(n235), .B(n419), .C(fr_enable), .Y(n422) );
  NAND2X1 U552 ( .A(n44), .B(n240), .Y(n421) );
  NAND2X1 U553 ( .A(n422), .B(n421), .Y(n1291) );
  OAI21X1 U554 ( .A(n235), .B(n423), .C(fw_enable), .Y(n426) );
  NAND2X1 U555 ( .A(n424), .B(n238), .Y(n425) );
  NAND2X1 U556 ( .A(n426), .B(n425), .Y(n1290) );
  MUX2X1 U557 ( .B(nfdata[0]), .A(fdata[0]), .S(n234), .Y(n427) );
  MUX2X1 U558 ( .B(nfdata[1]), .A(fdata[1]), .S(n234), .Y(n428) );
  MUX2X1 U559 ( .B(nfdata[2]), .A(fdata[2]), .S(n234), .Y(n429) );
  MUX2X1 U560 ( .B(nfdata[3]), .A(fdata[3]), .S(n234), .Y(n430) );
  MUX2X1 U561 ( .B(nfdata[4]), .A(fdata[4]), .S(n234), .Y(n431) );
  MUX2X1 U562 ( .B(nfdata[5]), .A(fdata[5]), .S(n234), .Y(n432) );
  INVX2 U563 ( .A(n432), .Y(n1284) );
  MUX2X1 U564 ( .B(nfdata[6]), .A(fdata[6]), .S(n234), .Y(n433) );
  MUX2X1 U565 ( .B(nfdata[7]), .A(fdata[7]), .S(n234), .Y(n434) );
  MUX2X1 U566 ( .B(nfaddr[0]), .A(ADDR[0]), .S(n233), .Y(n435) );
  INVX2 U567 ( .A(n435), .Y(n1281) );
  MUX2X1 U568 ( .B(nfaddr[0]), .A(faddr[0]), .S(n233), .Y(n436) );
  INVX2 U569 ( .A(n436), .Y(n1280) );
  MUX2X1 U570 ( .B(nfaddr[1]), .A(ADDR[1]), .S(n233), .Y(n437) );
  INVX2 U571 ( .A(n437), .Y(n1279) );
  MUX2X1 U572 ( .B(nfaddr[1]), .A(faddr[1]), .S(n233), .Y(n438) );
  INVX2 U573 ( .A(n438), .Y(n1278) );
  MUX2X1 U574 ( .B(nfaddr[2]), .A(ADDR[2]), .S(n233), .Y(n439) );
  INVX2 U575 ( .A(n439), .Y(n1277) );
  MUX2X1 U576 ( .B(nfaddr[2]), .A(faddr[2]), .S(n233), .Y(n440) );
  INVX2 U577 ( .A(n440), .Y(n1276) );
  MUX2X1 U578 ( .B(nfaddr[3]), .A(ADDR[3]), .S(n233), .Y(n441) );
  MUX2X1 U579 ( .B(nfaddr[3]), .A(faddr[3]), .S(n233), .Y(n442) );
  MUX2X1 U580 ( .B(nfaddr[4]), .A(ADDR[4]), .S(n233), .Y(n443) );
  INVX2 U581 ( .A(n443), .Y(n1273) );
  MUX2X1 U582 ( .B(nfaddr[4]), .A(faddr[4]), .S(n233), .Y(n444) );
  INVX2 U583 ( .A(n444), .Y(n1272) );
  MUX2X1 U584 ( .B(nfaddr[5]), .A(ADDR[5]), .S(n233), .Y(n445) );
  MUX2X1 U585 ( .B(nfaddr[5]), .A(faddr[5]), .S(n233), .Y(n446) );
  INVX2 U586 ( .A(n446), .Y(n1270) );
  MUX2X1 U587 ( .B(nfaddr[7]), .A(ADDR[7]), .S(n232), .Y(n449) );
  MUX2X1 U588 ( .B(nfaddr[7]), .A(faddr[7]), .S(n233), .Y(n450) );
  INVX2 U589 ( .A(n451), .Y(n488) );
  XOR2X1 U590 ( .A(delaydata[7]), .B(temp[7]), .Y(n457) );
  NOR2X1 U591 ( .A(n452), .B(n1073), .Y(n453) );
  NAND3X1 U592 ( .A(n5), .B(n454), .C(n453), .Y(n657) );
  NOR2X1 U593 ( .A(n37), .B(n220), .Y(n456) );
  NAND3X1 U594 ( .A(n654), .B(n182), .C(n456), .Y(n486) );
  AOI22X1 U595 ( .A(n488), .B(n457), .C(n45), .D(currentProcessedData[7]), .Y(
        n460) );
  NAND2X1 U596 ( .A(BYTE[7]), .B(n489), .Y(n459) );
  INVX2 U597 ( .A(PROCESSED_DATA[7]), .Y(n461) );
  MUX2X1 U598 ( .B(n134), .A(n461), .S(n232), .Y(n1265) );
  XOR2X1 U599 ( .A(delaydata[6]), .B(temp[6]), .Y(n462) );
  AOI22X1 U600 ( .A(n488), .B(n462), .C(n46), .D(currentProcessedData[6]), .Y(
        n464) );
  NAND2X1 U601 ( .A(BYTE[6]), .B(n489), .Y(n463) );
  INVX2 U602 ( .A(PROCESSED_DATA[6]), .Y(n465) );
  MUX2X1 U603 ( .B(n133), .A(n465), .S(n232), .Y(n1264) );
  XOR2X1 U604 ( .A(delaydata[5]), .B(temp[5]), .Y(n466) );
  AOI22X1 U605 ( .A(n488), .B(n466), .C(n45), .D(currentProcessedData[5]), .Y(
        n468) );
  NAND2X1 U606 ( .A(BYTE[5]), .B(n489), .Y(n467) );
  INVX2 U607 ( .A(PROCESSED_DATA[5]), .Y(n469) );
  MUX2X1 U608 ( .B(n132), .A(n469), .S(n232), .Y(n1263) );
  XOR2X1 U609 ( .A(delaydata[4]), .B(temp[4]), .Y(n470) );
  AOI22X1 U610 ( .A(n488), .B(n470), .C(n46), .D(currentProcessedData[4]), .Y(
        n472) );
  NAND2X1 U611 ( .A(BYTE[4]), .B(n489), .Y(n471) );
  INVX2 U612 ( .A(PROCESSED_DATA[4]), .Y(n473) );
  MUX2X1 U613 ( .B(n131), .A(n473), .S(n232), .Y(n1262) );
  XOR2X1 U614 ( .A(delaydata[3]), .B(temp[3]), .Y(n474) );
  AOI22X1 U615 ( .A(n488), .B(n474), .C(n45), .D(currentProcessedData[3]), .Y(
        n476) );
  NAND2X1 U616 ( .A(BYTE[3]), .B(n489), .Y(n475) );
  INVX2 U617 ( .A(PROCESSED_DATA[3]), .Y(n477) );
  MUX2X1 U618 ( .B(n129), .A(n477), .S(n232), .Y(n1261) );
  XOR2X1 U619 ( .A(delaydata[2]), .B(temp[2]), .Y(n478) );
  AOI22X1 U620 ( .A(n488), .B(n478), .C(n45), .D(currentProcessedData[2]), .Y(
        n480) );
  NAND2X1 U621 ( .A(BYTE[2]), .B(n489), .Y(n479) );
  INVX2 U622 ( .A(PROCESSED_DATA[2]), .Y(n481) );
  MUX2X1 U623 ( .B(n127), .A(n481), .S(n232), .Y(n1260) );
  XOR2X1 U624 ( .A(delaydata[1]), .B(temp[1]), .Y(n482) );
  AOI22X1 U625 ( .A(n488), .B(n482), .C(n46), .D(currentProcessedData[1]), .Y(
        n484) );
  NAND2X1 U626 ( .A(BYTE[1]), .B(n489), .Y(n483) );
  INVX2 U627 ( .A(PROCESSED_DATA[1]), .Y(n485) );
  MUX2X1 U628 ( .B(n125), .A(n485), .S(n232), .Y(n1259) );
  XOR2X1 U629 ( .A(delaydata[0]), .B(temp[0]), .Y(n487) );
  AOI22X1 U630 ( .A(n488), .B(n487), .C(n45), .D(currentProcessedData[0]), .Y(
        n491) );
  NAND2X1 U631 ( .A(BYTE[0]), .B(n489), .Y(n490) );
  INVX2 U632 ( .A(PROCESSED_DATA[0]), .Y(n492) );
  MUX2X1 U633 ( .B(n122), .A(n492), .S(n232), .Y(n1258) );
  NAND2X1 U634 ( .A(n102), .B(n164), .Y(n570) );
  NAND2X1 U635 ( .A(n161), .B(n1057), .Y(n1071) );
  INVX2 U636 ( .A(n1071), .Y(n494) );
  NAND2X1 U637 ( .A(n494), .B(n157), .Y(n571) );
  INVX2 U638 ( .A(n571), .Y(n495) );
  NAND3X1 U639 ( .A(n495), .B(n570), .C(n496), .Y(n638) );
  NAND2X1 U640 ( .A(n497), .B(n516), .Y(n515) );
  INVX2 U641 ( .A(N502), .Y(n499) );
  NAND3X1 U642 ( .A(n68), .B(n63), .C(n70), .Y(n512) );
  NAND2X1 U643 ( .A(inti[6]), .B(n512), .Y(n498) );
  OAI21X1 U644 ( .A(n515), .B(n499), .C(n498), .Y(n1124) );
  INVX2 U645 ( .A(N501), .Y(n501) );
  NAND2X1 U646 ( .A(inti[5]), .B(n512), .Y(n500) );
  OAI21X1 U647 ( .A(n515), .B(n501), .C(n500), .Y(n1123) );
  INVX2 U648 ( .A(N500), .Y(n503) );
  NAND2X1 U649 ( .A(inti[4]), .B(n512), .Y(n502) );
  OAI21X1 U650 ( .A(n515), .B(n503), .C(n502), .Y(n1122) );
  INVX2 U651 ( .A(N499), .Y(n505) );
  NAND2X1 U652 ( .A(inti[3]), .B(n512), .Y(n504) );
  OAI21X1 U653 ( .A(n515), .B(n505), .C(n504), .Y(n1121) );
  NAND2X1 U654 ( .A(inti[2]), .B(n512), .Y(n506) );
  OAI21X1 U655 ( .A(n515), .B(n507), .C(n506), .Y(n1120) );
  NAND2X1 U656 ( .A(inti[1]), .B(n512), .Y(n508) );
  OAI21X1 U657 ( .A(n515), .B(n509), .C(n508), .Y(n1119) );
  NAND2X1 U658 ( .A(inti[0]), .B(n512), .Y(n510) );
  OAI21X1 U659 ( .A(n515), .B(n511), .C(n510), .Y(n1118) );
  INVX2 U660 ( .A(N503), .Y(n514) );
  NAND2X1 U661 ( .A(inti[7]), .B(n512), .Y(n513) );
  OAI21X1 U662 ( .A(n515), .B(n514), .C(n513), .Y(n1125) );
  NAND3X1 U663 ( .A(keyi[2]), .B(n519), .C(n521), .Y(n517) );
  INVX2 U664 ( .A(n517), .Y(n559) );
  NAND3X1 U665 ( .A(keyi[2]), .B(keyi[0]), .C(n519), .Y(n518) );
  INVX2 U666 ( .A(n518), .Y(n558) );
  AOI22X1 U667 ( .A(\keyTable[4][7] ), .B(n559), .C(\keyTable[5][7] ), .D(n558), .Y(n527) );
  AOI22X1 U668 ( .A(\keyTable[6][7] ), .B(n191), .C(\keyTable[7][7] ), .D(n198), .Y(n526) );
  INVX2 U670 ( .A(\keyTable[3][7] ), .Y(n939) );
  NAND3X1 U671 ( .A(keyi[1]), .B(n520), .C(n521), .Y(n560) );
  INVX2 U672 ( .A(\keyTable[2][7] ), .Y(n923) );
  OAI22X1 U674 ( .A(n32), .B(n939), .C(n560), .D(n923), .Y(n524) );
  NAND3X1 U675 ( .A(keyi[0]), .B(n520), .C(n519), .Y(n562) );
  INVX2 U676 ( .A(\keyTable[1][7] ), .Y(n786) );
  NOR2X1 U677 ( .A(keyi[2]), .B(keyi[1]), .Y(n522) );
  NAND2X1 U678 ( .A(n522), .B(n521), .Y(n561) );
  INVX2 U679 ( .A(\keyTable[0][7] ), .Y(n784) );
  OAI22X1 U680 ( .A(n562), .B(n786), .C(n561), .D(n784), .Y(n523) );
  NOR2X1 U681 ( .A(n524), .B(n523), .Y(n525) );
  NAND3X1 U682 ( .A(n527), .B(n526), .C(n525), .Y(N472) );
  AOI22X1 U683 ( .A(\keyTable[4][6] ), .B(n559), .C(\keyTable[5][6] ), .D(n558), .Y(n532) );
  AOI22X1 U684 ( .A(\keyTable[6][6] ), .B(n191), .C(\keyTable[7][6] ), .D(n198), .Y(n531) );
  INVX2 U685 ( .A(\keyTable[3][6] ), .Y(n941) );
  INVX2 U686 ( .A(\keyTable[2][6] ), .Y(n925) );
  OAI22X1 U687 ( .A(n32), .B(n941), .C(n560), .D(n925), .Y(n529) );
  INVX2 U688 ( .A(\keyTable[1][6] ), .Y(n885) );
  INVX2 U689 ( .A(\keyTable[0][6] ), .Y(n883) );
  OAI22X1 U690 ( .A(n562), .B(n885), .C(n561), .D(n883), .Y(n528) );
  NOR2X1 U691 ( .A(n529), .B(n528), .Y(n530) );
  NAND3X1 U692 ( .A(n532), .B(n531), .C(n530), .Y(N473) );
  AOI22X1 U693 ( .A(\keyTable[4][5] ), .B(n559), .C(\keyTable[5][5] ), .D(n558), .Y(n537) );
  AOI22X1 U694 ( .A(\keyTable[6][5] ), .B(n191), .C(\keyTable[7][5] ), .D(n198), .Y(n536) );
  INVX2 U695 ( .A(\keyTable[3][5] ), .Y(n943) );
  INVX2 U696 ( .A(\keyTable[2][5] ), .Y(n927) );
  OAI22X1 U697 ( .A(n32), .B(n943), .C(n560), .D(n927), .Y(n534) );
  INVX2 U698 ( .A(\keyTable[1][5] ), .Y(n887) );
  INVX2 U699 ( .A(\keyTable[0][5] ), .Y(n870) );
  OAI22X1 U700 ( .A(n562), .B(n887), .C(n561), .D(n870), .Y(n533) );
  NOR2X1 U701 ( .A(n534), .B(n533), .Y(n535) );
  NAND3X1 U702 ( .A(n537), .B(n536), .C(n535), .Y(N474) );
  AOI22X1 U703 ( .A(\keyTable[4][4] ), .B(n559), .C(\keyTable[5][4] ), .D(n558), .Y(n542) );
  AOI22X1 U704 ( .A(\keyTable[6][4] ), .B(n191), .C(\keyTable[7][4] ), .D(n198), .Y(n541) );
  INVX2 U705 ( .A(\keyTable[3][4] ), .Y(n945) );
  INVX2 U706 ( .A(\keyTable[2][4] ), .Y(n929) );
  OAI22X1 U707 ( .A(n32), .B(n945), .C(n560), .D(n929), .Y(n539) );
  INVX2 U708 ( .A(\keyTable[1][4] ), .Y(n889) );
  INVX2 U709 ( .A(\keyTable[0][4] ), .Y(n868) );
  OAI22X1 U710 ( .A(n562), .B(n889), .C(n561), .D(n868), .Y(n538) );
  NOR2X1 U711 ( .A(n539), .B(n538), .Y(n540) );
  NAND3X1 U712 ( .A(n542), .B(n541), .C(n540), .Y(N475) );
  AOI22X1 U713 ( .A(\keyTable[4][3] ), .B(n559), .C(\keyTable[5][3] ), .D(n558), .Y(n547) );
  AOI22X1 U714 ( .A(\keyTable[6][3] ), .B(n191), .C(\keyTable[7][3] ), .D(n198), .Y(n546) );
  INVX2 U715 ( .A(\keyTable[3][3] ), .Y(n947) );
  INVX2 U716 ( .A(\keyTable[2][3] ), .Y(n931) );
  OAI22X1 U717 ( .A(n32), .B(n947), .C(n560), .D(n931), .Y(n544) );
  INVX2 U718 ( .A(\keyTable[1][3] ), .Y(n898) );
  INVX2 U719 ( .A(\keyTable[0][3] ), .Y(n866) );
  OAI22X1 U720 ( .A(n562), .B(n898), .C(n561), .D(n866), .Y(n543) );
  NOR2X1 U721 ( .A(n544), .B(n543), .Y(n545) );
  NAND3X1 U722 ( .A(n547), .B(n546), .C(n545), .Y(N476) );
  AOI22X1 U723 ( .A(\keyTable[4][2] ), .B(n559), .C(\keyTable[5][2] ), .D(n558), .Y(n552) );
  AOI22X1 U724 ( .A(\keyTable[6][2] ), .B(n191), .C(\keyTable[7][2] ), .D(n198), .Y(n551) );
  INVX2 U725 ( .A(\keyTable[3][2] ), .Y(n949) );
  INVX2 U726 ( .A(\keyTable[2][2] ), .Y(n933) );
  OAI22X1 U727 ( .A(n32), .B(n949), .C(n560), .D(n933), .Y(n549) );
  INVX2 U728 ( .A(\keyTable[1][2] ), .Y(n917) );
  INVX2 U729 ( .A(\keyTable[0][2] ), .Y(n864) );
  OAI22X1 U730 ( .A(n562), .B(n917), .C(n561), .D(n864), .Y(n548) );
  NOR2X1 U731 ( .A(n549), .B(n548), .Y(n550) );
  NAND3X1 U732 ( .A(n552), .B(n551), .C(n550), .Y(N477) );
  AOI22X1 U733 ( .A(\keyTable[4][1] ), .B(n559), .C(\keyTable[5][1] ), .D(n558), .Y(n557) );
  AOI22X1 U734 ( .A(\keyTable[6][1] ), .B(n191), .C(\keyTable[7][1] ), .D(n198), .Y(n556) );
  INVX2 U735 ( .A(\keyTable[3][1] ), .Y(n951) );
  INVX2 U736 ( .A(\keyTable[2][1] ), .Y(n935) );
  OAI22X1 U737 ( .A(n32), .B(n951), .C(n560), .D(n935), .Y(n554) );
  INVX2 U738 ( .A(\keyTable[1][1] ), .Y(n919) );
  INVX2 U739 ( .A(\keyTable[0][1] ), .Y(n790) );
  OAI22X1 U740 ( .A(n562), .B(n919), .C(n561), .D(n790), .Y(n553) );
  NOR2X1 U741 ( .A(n554), .B(n553), .Y(n555) );
  NAND3X1 U742 ( .A(n557), .B(n556), .C(n555), .Y(N478) );
  AOI22X1 U743 ( .A(\keyTable[4][0] ), .B(n559), .C(\keyTable[5][0] ), .D(n558), .Y(n567) );
  AOI22X1 U744 ( .A(\keyTable[6][0] ), .B(n191), .C(\keyTable[7][0] ), .D(n198), .Y(n566) );
  INVX2 U745 ( .A(\keyTable[3][0] ), .Y(n953) );
  INVX2 U746 ( .A(\keyTable[2][0] ), .Y(n937) );
  OAI22X1 U747 ( .A(n32), .B(n953), .C(n560), .D(n937), .Y(n564) );
  INVX2 U748 ( .A(\keyTable[1][0] ), .Y(n921) );
  INVX2 U749 ( .A(\keyTable[0][0] ), .Y(n788) );
  OAI22X1 U750 ( .A(n562), .B(n921), .C(n561), .D(n788), .Y(n563) );
  NOR2X1 U751 ( .A(n564), .B(n563), .Y(n565) );
  NAND3X1 U752 ( .A(n567), .B(n566), .C(n565), .Y(N479) );
  NAND3X1 U753 ( .A(n634), .B(n11), .C(n222), .Y(n568) );
  INVX2 U754 ( .A(n570), .Y(n572) );
  NOR3X1 U755 ( .A(n572), .B(n89), .C(n571), .Y(n573) );
  AND2X2 U756 ( .A(n574), .B(n573), .Y(n597) );
  NAND2X1 U757 ( .A(n597), .B(n109), .Y(n593) );
  INVX2 U758 ( .A(n593), .Y(n579) );
  INVX2 U759 ( .A(n58), .Y(n576) );
  NAND2X1 U760 ( .A(N480), .B(n590), .Y(n575) );
  OAI21X1 U761 ( .A(n579), .B(n576), .C(n575), .Y(n1161) );
  INVX2 U762 ( .A(sj[1]), .Y(n578) );
  NAND2X1 U763 ( .A(N481), .B(n590), .Y(n577) );
  OAI21X1 U764 ( .A(n579), .B(n578), .C(n577), .Y(n1160) );
  NAND2X1 U765 ( .A(sj[2]), .B(n593), .Y(n581) );
  NAND2X1 U766 ( .A(N482), .B(n590), .Y(n580) );
  NAND2X1 U767 ( .A(n581), .B(n580), .Y(n1159) );
  NAND2X1 U768 ( .A(sj[3]), .B(n593), .Y(n583) );
  NAND2X1 U769 ( .A(N483), .B(n590), .Y(n582) );
  NAND2X1 U770 ( .A(n583), .B(n582), .Y(n1158) );
  NAND2X1 U771 ( .A(sj[4]), .B(n593), .Y(n585) );
  NAND2X1 U772 ( .A(N484), .B(n590), .Y(n584) );
  NAND2X1 U773 ( .A(n585), .B(n584), .Y(n1157) );
  NAND2X1 U774 ( .A(sj[5]), .B(n593), .Y(n587) );
  NAND2X1 U775 ( .A(N485), .B(n590), .Y(n586) );
  NAND2X1 U776 ( .A(n587), .B(n586), .Y(n1156) );
  NAND2X1 U777 ( .A(sj[6]), .B(n593), .Y(n592) );
  NAND2X1 U778 ( .A(N486), .B(n590), .Y(n591) );
  NAND2X1 U779 ( .A(n592), .B(n591), .Y(n1155) );
  NAND2X1 U780 ( .A(sj[7]), .B(n593), .Y(n595) );
  INVX2 U781 ( .A(N487), .Y(n594) );
  AOI22X1 U782 ( .A(n595), .B(n170), .C(n595), .D(n594), .Y(n1098) );
  NOR2X1 U783 ( .A(n235), .B(n596), .Y(n598) );
  NAND3X1 U784 ( .A(n598), .B(n1088), .C(n597), .Y(n613) );
  INVX2 U785 ( .A(n613), .Y(n617) );
  INVX2 U786 ( .A(N518), .Y(n600) );
  NAND2X1 U787 ( .A(intj[6]), .B(n201), .Y(n599) );
  OAI21X1 U788 ( .A(n616), .B(n600), .C(n599), .Y(n1168) );
  INVX2 U789 ( .A(N517), .Y(n602) );
  NAND2X1 U790 ( .A(intj[5]), .B(n201), .Y(n601) );
  OAI21X1 U791 ( .A(n616), .B(n602), .C(n601), .Y(n1167) );
  INVX2 U792 ( .A(N516), .Y(n604) );
  NAND2X1 U793 ( .A(intj[4]), .B(n201), .Y(n603) );
  OAI21X1 U794 ( .A(n616), .B(n604), .C(n603), .Y(n1166) );
  INVX2 U795 ( .A(N515), .Y(n606) );
  NAND2X1 U796 ( .A(intj[3]), .B(n201), .Y(n605) );
  OAI21X1 U797 ( .A(n616), .B(n606), .C(n605), .Y(n1165) );
  INVX2 U798 ( .A(N514), .Y(n608) );
  NAND2X1 U799 ( .A(intj[2]), .B(n201), .Y(n607) );
  OAI21X1 U800 ( .A(n616), .B(n608), .C(n607), .Y(n1164) );
  INVX2 U801 ( .A(N513), .Y(n610) );
  NAND2X1 U802 ( .A(intj[1]), .B(n201), .Y(n609) );
  OAI21X1 U803 ( .A(n616), .B(n610), .C(n609), .Y(n1163) );
  INVX2 U804 ( .A(N512), .Y(n612) );
  NAND2X1 U805 ( .A(intj[0]), .B(n201), .Y(n611) );
  OAI21X1 U806 ( .A(n616), .B(n612), .C(n611), .Y(n1162) );
  INVX2 U807 ( .A(N519), .Y(n615) );
  NAND2X1 U808 ( .A(intj[7]), .B(n201), .Y(n614) );
  OAI21X1 U809 ( .A(n616), .B(n615), .C(n614), .Y(n1169) );
  INVX2 U810 ( .A(delaydata[6]), .Y(n619) );
  INVX2 U811 ( .A(BYTE[6]), .Y(n618) );
  MUX2X1 U812 ( .B(n619), .A(n618), .S(n218), .Y(n1111) );
  INVX2 U813 ( .A(delaydata[5]), .Y(n621) );
  INVX2 U814 ( .A(BYTE[5]), .Y(n620) );
  MUX2X1 U815 ( .B(n621), .A(n620), .S(n217), .Y(n1112) );
  INVX2 U816 ( .A(delaydata[4]), .Y(n623) );
  INVX2 U817 ( .A(BYTE[4]), .Y(n622) );
  MUX2X1 U818 ( .B(n623), .A(n622), .S(n218), .Y(n1113) );
  INVX2 U819 ( .A(delaydata[3]), .Y(n625) );
  INVX2 U820 ( .A(BYTE[3]), .Y(n624) );
  MUX2X1 U821 ( .B(n625), .A(n624), .S(n217), .Y(n1114) );
  INVX2 U822 ( .A(delaydata[2]), .Y(n627) );
  INVX2 U823 ( .A(BYTE[2]), .Y(n626) );
  MUX2X1 U824 ( .B(n627), .A(n626), .S(n218), .Y(n1115) );
  INVX2 U825 ( .A(delaydata[1]), .Y(n629) );
  INVX2 U826 ( .A(BYTE[1]), .Y(n628) );
  MUX2X1 U827 ( .B(n629), .A(n628), .S(n217), .Y(n1116) );
  INVX2 U828 ( .A(delaydata[0]), .Y(n631) );
  INVX2 U829 ( .A(BYTE[0]), .Y(n630) );
  MUX2X1 U830 ( .B(n631), .A(n630), .S(n218), .Y(n1117) );
  INVX2 U831 ( .A(delaydata[7]), .Y(n633) );
  INVX2 U832 ( .A(BYTE[7]), .Y(n632) );
  MUX2X1 U833 ( .B(n633), .A(n632), .S(n217), .Y(n1110) );
  NAND3X1 U834 ( .A(si[3]), .B(si[2]), .C(si[6]), .Y(n636) );
  NAND2X1 U835 ( .A(n1319), .B(si[7]), .Y(n635) );
  NOR2X1 U836 ( .A(n636), .B(n635), .Y(n637) );
  NAND2X1 U837 ( .A(n637), .B(n1318), .Y(n1051) );
  NAND2X1 U838 ( .A(N431), .B(n8), .Y(n641) );
  NAND2X1 U839 ( .A(n113), .B(n639), .Y(n644) );
  NAND2X1 U840 ( .A(si[7]), .B(n644), .Y(n640) );
  NAND2X1 U841 ( .A(n641), .B(n640), .Y(n1153) );
  NAND2X1 U842 ( .A(N430), .B(n8), .Y(n643) );
  NAND2X1 U843 ( .A(si[6]), .B(n644), .Y(n642) );
  NAND2X1 U844 ( .A(n643), .B(n642), .Y(n1152) );
  INVX2 U845 ( .A(n644), .Y(n653) );
  NAND2X1 U846 ( .A(N429), .B(n8), .Y(n645) );
  OAI21X1 U847 ( .A(n1104), .B(n653), .C(n645), .Y(n1151) );
  NAND2X1 U848 ( .A(N428), .B(n8), .Y(n646) );
  OAI21X1 U849 ( .A(n1103), .B(n653), .C(n646), .Y(n1150) );
  NAND2X1 U850 ( .A(N427), .B(n8), .Y(n647) );
  OAI21X1 U851 ( .A(n653), .B(n648), .C(n647), .Y(n1149) );
  NAND2X1 U852 ( .A(N426), .B(n8), .Y(n649) );
  OAI21X1 U853 ( .A(n653), .B(n650), .C(n649), .Y(n1148) );
  NAND2X1 U854 ( .A(N425), .B(n8), .Y(n651) );
  OAI21X1 U855 ( .A(n1102), .B(n653), .C(n651), .Y(n1147) );
  NAND2X1 U856 ( .A(N424), .B(n8), .Y(n652) );
  OAI21X1 U857 ( .A(n1101), .B(n653), .C(n652), .Y(n1146) );
  NAND2X1 U858 ( .A(n222), .B(n654), .Y(n655) );
  NAND2X1 U859 ( .A(n106), .B(n237), .Y(n658) );
  NOR3X1 U860 ( .A(n658), .B(n220), .C(n656), .Y(n659) );
  NAND2X1 U861 ( .A(n660), .B(n659), .Y(n683) );
  NAND2X1 U862 ( .A(temp[6]), .B(n115), .Y(n663) );
  NAND3X1 U863 ( .A(DATA_IN[6]), .B(n6), .C(n684), .Y(n662) );
  INVX2 U864 ( .A(n202), .Y(n685) );
  NAND3X1 U865 ( .A(N526), .B(n685), .C(n684), .Y(n661) );
  NAND3X1 U866 ( .A(n663), .B(n662), .C(n661), .Y(n1179) );
  NAND2X1 U867 ( .A(temp[5]), .B(n115), .Y(n666) );
  NAND3X1 U868 ( .A(DATA_IN[5]), .B(n6), .C(n684), .Y(n665) );
  NAND3X1 U869 ( .A(N525), .B(n685), .C(n93), .Y(n664) );
  NAND3X1 U870 ( .A(n666), .B(n665), .C(n664), .Y(n1178) );
  NAND2X1 U871 ( .A(temp[4]), .B(n91), .Y(n669) );
  NAND3X1 U872 ( .A(DATA_IN[4]), .B(n6), .C(n93), .Y(n668) );
  NAND3X1 U873 ( .A(N524), .B(n685), .C(n684), .Y(n667) );
  NAND3X1 U874 ( .A(n669), .B(n668), .C(n667), .Y(n1177) );
  NAND2X1 U875 ( .A(temp[3]), .B(n91), .Y(n672) );
  NAND3X1 U876 ( .A(DATA_IN[3]), .B(n6), .C(n93), .Y(n671) );
  NAND3X1 U877 ( .A(N523), .B(n685), .C(n93), .Y(n670) );
  NAND3X1 U878 ( .A(n672), .B(n671), .C(n670), .Y(n1176) );
  NAND2X1 U879 ( .A(temp[2]), .B(n115), .Y(n675) );
  NAND3X1 U880 ( .A(DATA_IN[2]), .B(n6), .C(n684), .Y(n674) );
  NAND3X1 U881 ( .A(N522), .B(n685), .C(n93), .Y(n673) );
  NAND3X1 U882 ( .A(n675), .B(n674), .C(n673), .Y(n1175) );
  NAND2X1 U883 ( .A(temp[1]), .B(n91), .Y(n678) );
  NAND3X1 U884 ( .A(DATA_IN[1]), .B(n6), .C(n93), .Y(n677) );
  NAND3X1 U885 ( .A(N521), .B(n685), .C(n684), .Y(n676) );
  NAND3X1 U886 ( .A(n678), .B(n677), .C(n676), .Y(n1174) );
  NAND2X1 U887 ( .A(temp[0]), .B(n76), .Y(n682) );
  NAND3X1 U888 ( .A(DATA_IN[0]), .B(n6), .C(n684), .Y(n681) );
  NAND3X1 U889 ( .A(N520), .B(n685), .C(n93), .Y(n680) );
  NAND3X1 U890 ( .A(n682), .B(n681), .C(n680), .Y(n1173) );
  NAND2X1 U891 ( .A(temp[7]), .B(n115), .Y(n688) );
  NAND3X1 U892 ( .A(DATA_IN[7]), .B(n6), .C(n93), .Y(n687) );
  NAND3X1 U893 ( .A(N527), .B(n685), .C(n684), .Y(n686) );
  NAND3X1 U894 ( .A(n688), .B(n687), .C(n686), .Y(n1180) );
  NOR2X1 U895 ( .A(n692), .B(n690), .Y(n1020) );
  NAND2X1 U896 ( .A(n104), .B(n1018), .Y(n1097) );
  INVX2 U897 ( .A(N413), .Y(n750) );
  NAND2X1 U898 ( .A(prefillCounter[6]), .B(n1094), .Y(n748) );
  OAI21X1 U899 ( .A(n61), .B(n750), .C(n748), .Y(n1145) );
  INVX2 U900 ( .A(N412), .Y(n754) );
  NAND2X1 U901 ( .A(n1094), .B(prefillCounter[5]), .Y(n752) );
  OAI21X1 U902 ( .A(n61), .B(n754), .C(n752), .Y(n1144) );
  INVX2 U903 ( .A(N411), .Y(n758) );
  NAND2X1 U904 ( .A(prefillCounter[4]), .B(n1094), .Y(n756) );
  OAI21X1 U905 ( .A(n62), .B(n758), .C(n756), .Y(n1143) );
  INVX2 U906 ( .A(N410), .Y(n765) );
  NAND2X1 U907 ( .A(prefillCounter[3]), .B(n1094), .Y(n760) );
  OAI21X1 U908 ( .A(n62), .B(n765), .C(n760), .Y(n1142) );
  INVX2 U909 ( .A(N409), .Y(n767) );
  NAND2X1 U914 ( .A(prefillCounter[2]), .B(n1094), .Y(n766) );
  OAI21X1 U915 ( .A(n62), .B(n767), .C(n766), .Y(n1141) );
  INVX2 U916 ( .A(N408), .Y(n769) );
  NAND2X1 U917 ( .A(prefillCounter[1]), .B(n1094), .Y(n768) );
  OAI21X1 U918 ( .A(n62), .B(n769), .C(n768), .Y(n1140) );
  INVX2 U920 ( .A(N414), .Y(n772) );
  NAND2X1 U921 ( .A(prefillCounter[7]), .B(n1094), .Y(n771) );
  OAI21X1 U922 ( .A(n61), .B(n772), .C(n771), .Y(n1139) );
  INVX2 U923 ( .A(KEY[7]), .Y(n783) );
  NOR2X1 U932 ( .A(n89), .B(n773), .Y(n774) );
  MUX2X1 U933 ( .B(n784), .A(n783), .S(n138), .Y(n1181) );
  INVX2 U934 ( .A(KEY[15]), .Y(n785) );
  MUX2X1 U935 ( .B(n786), .A(n785), .S(n141), .Y(n1182) );
  INVX2 U936 ( .A(KEY[0]), .Y(n787) );
  MUX2X1 U937 ( .B(n788), .A(n787), .S(n138), .Y(n1183) );
  INVX2 U938 ( .A(KEY[1]), .Y(n789) );
  MUX2X1 U939 ( .B(n790), .A(n789), .S(n138), .Y(n1184) );
  INVX2 U940 ( .A(KEY[2]), .Y(n791) );
  MUX2X1 U941 ( .B(n864), .A(n791), .S(n143), .Y(n1185) );
  INVX2 U942 ( .A(KEY[3]), .Y(n865) );
  MUX2X1 U943 ( .B(n866), .A(n865), .S(n138), .Y(n1186) );
  INVX2 U944 ( .A(KEY[4]), .Y(n867) );
  MUX2X1 U945 ( .B(n868), .A(n867), .S(n142), .Y(n1187) );
  INVX2 U946 ( .A(KEY[5]), .Y(n869) );
  MUX2X1 U947 ( .B(n870), .A(n869), .S(n142), .Y(n1188) );
  INVX2 U948 ( .A(KEY[6]), .Y(n871) );
  MUX2X1 U949 ( .B(n883), .A(n871), .S(n140), .Y(n1189) );
  INVX2 U950 ( .A(KEY[14]), .Y(n884) );
  MUX2X1 U951 ( .B(n885), .A(n884), .S(n143), .Y(n1190) );
  INVX2 U952 ( .A(KEY[13]), .Y(n886) );
  MUX2X1 U953 ( .B(n887), .A(n886), .S(n139), .Y(n1191) );
  INVX2 U954 ( .A(KEY[12]), .Y(n888) );
  MUX2X1 U955 ( .B(n889), .A(n888), .S(n139), .Y(n1192) );
  INVX2 U956 ( .A(KEY[11]), .Y(n890) );
  MUX2X1 U957 ( .B(n898), .A(n890), .S(n139), .Y(n1193) );
  INVX2 U958 ( .A(KEY[10]), .Y(n916) );
  MUX2X1 U959 ( .B(n917), .A(n916), .S(n140), .Y(n1194) );
  INVX2 U960 ( .A(KEY[9]), .Y(n918) );
  MUX2X1 U961 ( .B(n919), .A(n918), .S(n142), .Y(n1195) );
  INVX2 U962 ( .A(KEY[8]), .Y(n920) );
  MUX2X1 U963 ( .B(n921), .A(n920), .S(n140), .Y(n1196) );
  INVX2 U964 ( .A(KEY[23]), .Y(n922) );
  MUX2X1 U965 ( .B(n923), .A(n922), .S(n138), .Y(n1197) );
  INVX2 U966 ( .A(KEY[22]), .Y(n924) );
  MUX2X1 U967 ( .B(n925), .A(n924), .S(n138), .Y(n1198) );
  INVX2 U968 ( .A(KEY[21]), .Y(n926) );
  MUX2X1 U969 ( .B(n927), .A(n926), .S(n138), .Y(n1199) );
  INVX2 U970 ( .A(KEY[20]), .Y(n928) );
  MUX2X1 U971 ( .B(n929), .A(n928), .S(n138), .Y(n1200) );
  INVX2 U972 ( .A(KEY[19]), .Y(n930) );
  MUX2X1 U973 ( .B(n931), .A(n930), .S(n138), .Y(n1201) );
  INVX2 U974 ( .A(KEY[18]), .Y(n932) );
  MUX2X1 U975 ( .B(n933), .A(n932), .S(n141), .Y(n1202) );
  INVX2 U976 ( .A(KEY[17]), .Y(n934) );
  MUX2X1 U977 ( .B(n935), .A(n934), .S(n139), .Y(n1203) );
  INVX2 U978 ( .A(KEY[16]), .Y(n936) );
  MUX2X1 U979 ( .B(n937), .A(n936), .S(n138), .Y(n1204) );
  INVX2 U980 ( .A(KEY[31]), .Y(n938) );
  MUX2X1 U981 ( .B(n939), .A(n938), .S(n139), .Y(n1205) );
  INVX2 U982 ( .A(KEY[30]), .Y(n940) );
  MUX2X1 U983 ( .B(n941), .A(n940), .S(n143), .Y(n1206) );
  INVX2 U984 ( .A(KEY[29]), .Y(n942) );
  MUX2X1 U985 ( .B(n943), .A(n942), .S(n141), .Y(n1207) );
  INVX2 U986 ( .A(KEY[28]), .Y(n944) );
  MUX2X1 U987 ( .B(n945), .A(n944), .S(n143), .Y(n1208) );
  INVX2 U988 ( .A(KEY[27]), .Y(n946) );
  MUX2X1 U989 ( .B(n947), .A(n946), .S(n141), .Y(n1209) );
  INVX2 U990 ( .A(KEY[26]), .Y(n948) );
  MUX2X1 U991 ( .B(n949), .A(n948), .S(n140), .Y(n1210) );
  INVX2 U992 ( .A(KEY[25]), .Y(n950) );
  MUX2X1 U993 ( .B(n951), .A(n950), .S(n143), .Y(n1211) );
  INVX2 U994 ( .A(KEY[24]), .Y(n952) );
  MUX2X1 U995 ( .B(n953), .A(n952), .S(n142), .Y(n1212) );
  INVX2 U996 ( .A(\keyTable[4][7] ), .Y(n955) );
  INVX2 U997 ( .A(KEY[39]), .Y(n954) );
  MUX2X1 U998 ( .B(n955), .A(n954), .S(n142), .Y(n1213) );
  INVX2 U999 ( .A(\keyTable[4][6] ), .Y(n957) );
  INVX2 U1000 ( .A(KEY[38]), .Y(n956) );
  MUX2X1 U1001 ( .B(n957), .A(n956), .S(n140), .Y(n1214) );
  INVX2 U1002 ( .A(\keyTable[4][5] ), .Y(n959) );
  INVX2 U1003 ( .A(KEY[37]), .Y(n958) );
  MUX2X1 U1004 ( .B(n959), .A(n958), .S(n142), .Y(n1215) );
  INVX2 U1005 ( .A(\keyTable[4][4] ), .Y(n961) );
  INVX2 U1006 ( .A(KEY[36]), .Y(n960) );
  MUX2X1 U1007 ( .B(n961), .A(n960), .S(n140), .Y(n1216) );
  INVX2 U1008 ( .A(\keyTable[4][3] ), .Y(n963) );
  INVX2 U1009 ( .A(KEY[35]), .Y(n962) );
  MUX2X1 U1010 ( .B(n963), .A(n962), .S(n139), .Y(n1217) );
  INVX2 U1011 ( .A(\keyTable[4][2] ), .Y(n965) );
  INVX2 U1012 ( .A(KEY[34]), .Y(n964) );
  MUX2X1 U1013 ( .B(n965), .A(n964), .S(n143), .Y(n1218) );
  INVX2 U1014 ( .A(\keyTable[4][1] ), .Y(n967) );
  INVX2 U1015 ( .A(KEY[33]), .Y(n966) );
  MUX2X1 U1016 ( .B(n967), .A(n966), .S(n142), .Y(n1219) );
  INVX2 U1017 ( .A(\keyTable[4][0] ), .Y(n969) );
  INVX2 U1018 ( .A(KEY[32]), .Y(n968) );
  MUX2X1 U1019 ( .B(n969), .A(n968), .S(n141), .Y(n1220) );
  INVX2 U1020 ( .A(\keyTable[5][7] ), .Y(n971) );
  INVX2 U1021 ( .A(KEY[47]), .Y(n970) );
  MUX2X1 U1022 ( .B(n971), .A(n970), .S(n139), .Y(n1221) );
  INVX2 U1023 ( .A(\keyTable[5][6] ), .Y(n973) );
  INVX2 U1024 ( .A(KEY[46]), .Y(n972) );
  MUX2X1 U1025 ( .B(n973), .A(n972), .S(n141), .Y(n1222) );
  INVX2 U1026 ( .A(\keyTable[5][5] ), .Y(n975) );
  INVX2 U1027 ( .A(KEY[45]), .Y(n974) );
  MUX2X1 U1028 ( .B(n975), .A(n974), .S(n141), .Y(n1223) );
  INVX2 U1029 ( .A(\keyTable[5][4] ), .Y(n977) );
  INVX2 U1030 ( .A(KEY[44]), .Y(n976) );
  MUX2X1 U1031 ( .B(n977), .A(n976), .S(n139), .Y(n1224) );
  INVX2 U1032 ( .A(\keyTable[5][3] ), .Y(n979) );
  INVX2 U1033 ( .A(KEY[43]), .Y(n978) );
  MUX2X1 U1034 ( .B(n979), .A(n978), .S(n141), .Y(n1225) );
  INVX2 U1035 ( .A(\keyTable[5][2] ), .Y(n981) );
  INVX2 U1036 ( .A(KEY[42]), .Y(n980) );
  MUX2X1 U1037 ( .B(n981), .A(n980), .S(n141), .Y(n1226) );
  INVX2 U1038 ( .A(\keyTable[5][1] ), .Y(n983) );
  INVX2 U1039 ( .A(KEY[41]), .Y(n982) );
  MUX2X1 U1040 ( .B(n983), .A(n982), .S(n141), .Y(n1227) );
  INVX2 U1041 ( .A(\keyTable[5][0] ), .Y(n985) );
  INVX2 U1042 ( .A(KEY[40]), .Y(n984) );
  MUX2X1 U1043 ( .B(n985), .A(n984), .S(n143), .Y(n1228) );
  INVX2 U1044 ( .A(\keyTable[6][7] ), .Y(n987) );
  INVX2 U1045 ( .A(KEY[55]), .Y(n986) );
  MUX2X1 U1046 ( .B(n987), .A(n986), .S(n140), .Y(n1229) );
  INVX2 U1047 ( .A(\keyTable[6][6] ), .Y(n989) );
  INVX2 U1048 ( .A(KEY[54]), .Y(n988) );
  MUX2X1 U1049 ( .B(n989), .A(n988), .S(n143), .Y(n1230) );
  INVX2 U1050 ( .A(\keyTable[6][5] ), .Y(n991) );
  INVX2 U1051 ( .A(KEY[53]), .Y(n990) );
  MUX2X1 U1052 ( .B(n991), .A(n990), .S(n141), .Y(n1231) );
  INVX2 U1053 ( .A(\keyTable[6][4] ), .Y(n993) );
  INVX2 U1054 ( .A(KEY[52]), .Y(n992) );
  MUX2X1 U1055 ( .B(n993), .A(n992), .S(n139), .Y(n1232) );
  INVX2 U1056 ( .A(\keyTable[6][3] ), .Y(n995) );
  INVX2 U1057 ( .A(KEY[51]), .Y(n994) );
  MUX2X1 U1058 ( .B(n995), .A(n994), .S(n143), .Y(n1233) );
  INVX2 U1059 ( .A(\keyTable[6][2] ), .Y(n997) );
  INVX2 U1060 ( .A(KEY[50]), .Y(n996) );
  MUX2X1 U1061 ( .B(n997), .A(n996), .S(n142), .Y(n1234) );
  INVX2 U1062 ( .A(\keyTable[6][1] ), .Y(n999) );
  INVX2 U1063 ( .A(KEY[49]), .Y(n998) );
  MUX2X1 U1064 ( .B(n999), .A(n998), .S(n140), .Y(n1235) );
  INVX2 U1065 ( .A(\keyTable[6][0] ), .Y(n1001) );
  INVX2 U1066 ( .A(KEY[48]), .Y(n1000) );
  MUX2X1 U1067 ( .B(n1001), .A(n1000), .S(n140), .Y(n1236) );
  INVX2 U1068 ( .A(\keyTable[7][7] ), .Y(n1003) );
  INVX2 U1069 ( .A(KEY[63]), .Y(n1002) );
  MUX2X1 U1070 ( .B(n1003), .A(n1002), .S(n140), .Y(n1237) );
  INVX2 U1071 ( .A(\keyTable[7][6] ), .Y(n1005) );
  INVX2 U1072 ( .A(KEY[62]), .Y(n1004) );
  MUX2X1 U1073 ( .B(n1005), .A(n1004), .S(n139), .Y(n1238) );
  INVX2 U1074 ( .A(\keyTable[7][5] ), .Y(n1007) );
  INVX2 U1075 ( .A(KEY[61]), .Y(n1006) );
  MUX2X1 U1076 ( .B(n1007), .A(n1006), .S(n142), .Y(n1239) );
  INVX2 U1077 ( .A(\keyTable[7][4] ), .Y(n1009) );
  INVX2 U1078 ( .A(KEY[60]), .Y(n1008) );
  MUX2X1 U1079 ( .B(n1009), .A(n1008), .S(n143), .Y(n1240) );
  INVX2 U1080 ( .A(\keyTable[7][3] ), .Y(n1011) );
  INVX2 U1081 ( .A(KEY[59]), .Y(n1010) );
  MUX2X1 U1082 ( .B(n1011), .A(n1010), .S(n143), .Y(n1241) );
  INVX2 U1083 ( .A(\keyTable[7][2] ), .Y(n1013) );
  INVX2 U1084 ( .A(KEY[58]), .Y(n1012) );
  MUX2X1 U1085 ( .B(n1013), .A(n1012), .S(n139), .Y(n1242) );
  INVX2 U1086 ( .A(\keyTable[7][1] ), .Y(n1015) );
  INVX2 U1087 ( .A(KEY[57]), .Y(n1014) );
  MUX2X1 U1088 ( .B(n1015), .A(n1014), .S(n140), .Y(n1243) );
  INVX2 U1089 ( .A(\keyTable[7][0] ), .Y(n1017) );
  INVX2 U1090 ( .A(KEY[56]), .Y(n1016) );
  MUX2X1 U1091 ( .B(n1017), .A(n1016), .S(n142), .Y(n1244) );
  INVX2 U1092 ( .A(extratemp[0]), .Y(n1023) );
  INVX2 U1093 ( .A(DATA_IN[0]), .Y(n1022) );
  AOI21X1 U1094 ( .A(n88), .B(n51), .C(n1018), .Y(n1019) );
  MUX2X1 U1095 ( .B(n1023), .A(n1022), .S(n1036), .Y(n1126) );
  INVX2 U1096 ( .A(extratemp[1]), .Y(n1025) );
  INVX2 U1097 ( .A(DATA_IN[1]), .Y(n1024) );
  MUX2X1 U1098 ( .B(n1025), .A(n1024), .S(n1036), .Y(n1127) );
  INVX2 U1099 ( .A(extratemp[2]), .Y(n1027) );
  INVX2 U1100 ( .A(DATA_IN[2]), .Y(n1026) );
  MUX2X1 U1101 ( .B(n1027), .A(n1026), .S(n1036), .Y(n1128) );
  INVX2 U1102 ( .A(extratemp[3]), .Y(n1029) );
  INVX2 U1103 ( .A(DATA_IN[3]), .Y(n1028) );
  MUX2X1 U1104 ( .B(n1029), .A(n1028), .S(n1036), .Y(n1129) );
  INVX2 U1105 ( .A(extratemp[4]), .Y(n1031) );
  INVX2 U1106 ( .A(DATA_IN[4]), .Y(n1030) );
  MUX2X1 U1107 ( .B(n1031), .A(n1030), .S(n1036), .Y(n1130) );
  INVX2 U1108 ( .A(extratemp[5]), .Y(n1033) );
  INVX2 U1109 ( .A(DATA_IN[5]), .Y(n1032) );
  MUX2X1 U1110 ( .B(n1033), .A(n1032), .S(n1036), .Y(n1131) );
  INVX2 U1111 ( .A(extratemp[6]), .Y(n1035) );
  INVX2 U1112 ( .A(DATA_IN[6]), .Y(n1034) );
  MUX2X1 U1113 ( .B(n1035), .A(n1034), .S(n1036), .Y(n1132) );
  INVX2 U1114 ( .A(extratemp[7]), .Y(n1038) );
  INVX2 U1115 ( .A(DATA_IN[7]), .Y(n1037) );
  MUX2X1 U1116 ( .B(n1038), .A(n1037), .S(n1036), .Y(n1133) );
  AOI21X1 U1117 ( .A(n1041), .B(n1040), .C(n1134), .Y(n1049) );
  NAND2X1 U1118 ( .A(permuteComplete), .B(n1042), .Y(n1043) );
  NAND3X1 U1119 ( .A(n177), .B(n121), .C(n1043), .Y(n1089) );
  INVX2 U1120 ( .A(n1089), .Y(n1048) );
  OAI21X1 U1121 ( .A(n49), .B(n209), .C(n118), .Y(n1045) );
  AOI22X1 U1122 ( .A(n1105), .B(n1046), .C(n51), .D(n1045), .Y(n1047) );
  NAND3X1 U1123 ( .A(n1049), .B(n1048), .C(n1047), .Y(nextState[3]) );
  OAI21X1 U1124 ( .A(n1054), .B(n1051), .C(n1050), .Y(n1052) );
  NAND2X1 U1125 ( .A(n1053), .B(n1052), .Y(n1056) );
  NAND2X1 U1126 ( .A(permuteComplete), .B(n1054), .Y(n1055) );
  NAND2X1 U1127 ( .A(n1056), .B(n1055), .Y(n1154) );
  NAND3X1 U1128 ( .A(n1107), .B(BYTE_READY), .C(n1083), .Y(n1060) );
  NAND2X1 U1129 ( .A(n1332), .B(n1082), .Y(n1059) );
  NAND2X1 U1130 ( .A(n154), .B(n164), .Y(n1058) );
  NAND3X1 U1131 ( .A(n1060), .B(n1059), .C(n1058), .Y(n1062) );
  AOI21X1 U1132 ( .A(n1062), .B(n1105), .C(n1061), .Y(n1067) );
  NAND2X1 U1133 ( .A(n342), .B(n48), .Y(n1064) );
  NOR3X1 U1134 ( .A(n1065), .B(n1064), .C(n1134), .Y(n1066) );
  NAND3X1 U1135 ( .A(n203), .B(n1067), .C(n1066), .Y(nextState[0]) );
  NAND2X1 U1136 ( .A(n49), .B(n164), .Y(n1079) );
  INVX2 U1137 ( .A(n1334), .Y(n1070) );
  NAND2X1 U1138 ( .A(n1071), .B(n1070), .Y(n1078) );
  NAND2X1 U1139 ( .A(n1074), .B(n94), .Y(n1075) );
  AOI21X1 U1140 ( .A(n1333), .B(n1076), .C(n1075), .Y(n1077) );
  NAND3X1 U1141 ( .A(n1079), .B(n1078), .C(n1077), .Y(nextState[4]) );
  AND2X2 U1142 ( .A(n41), .B(n74), .Y(n1081) );
  MUX2X1 U1143 ( .B(n1041), .A(n1081), .S(n209), .Y(n1093) );
  NAND2X1 U1144 ( .A(n1330), .B(n1082), .Y(n1085) );
  NAND2X1 U1145 ( .A(n1329), .B(n1083), .Y(n1084) );
  NAND2X1 U1146 ( .A(n1085), .B(n1084), .Y(n1086) );
  NAND2X1 U1147 ( .A(n1086), .B(n1105), .Y(n1092) );
  NAND2X1 U1148 ( .A(n170), .B(n1087), .Y(n1090) );
  NOR2X1 U1149 ( .A(n1090), .B(n1089), .Y(n1091) );
  NAND3X1 U1150 ( .A(n1093), .B(n1092), .C(n1091), .Y(nextState[2]) );
  INVX2 U1151 ( .A(N407), .Y(n1096) );
  NAND2X1 U1152 ( .A(prefillCounter[0]), .B(n1094), .Y(n1095) );
  OAI21X1 U1153 ( .A(n61), .B(n1096), .C(n1095), .Y(n1138) );
  INVX2 U1154 ( .A(KEY_ERROR), .Y(n1105) );
  INVX2 U1155 ( .A(BYTE_READY), .Y(n1106) );
  INVX2 U1156 ( .A(n1331), .Y(n1107) );
  INVX2 U1157 ( .A(OPCODE[1]), .Y(n1108) );
  INVX2 U1158 ( .A(OPCODE[0]), .Y(n1109) );
endmodule


module uart_edge_detector_0 ( CLK, RST, SERIAL_IN, START_BIT );
  input CLK, RST, SERIAL_IN;
  output START_BIT;
  wire   Q_int, Q_int2, n2, n4;

  DFFSR Q_int_reg ( .D(SERIAL_IN), .CLK(CLK), .R(n2), .S(1'b1), .Q(Q_int) );
  DFFSR Q_int2_reg ( .D(Q_int), .CLK(CLK), .R(n2), .S(1'b1), .Q(Q_int2) );
  NOR2X1 U7 ( .A(Q_int), .B(n4), .Y(START_BIT) );
  INVX2 U4 ( .A(RST), .Y(n2) );
  INVX2 U6 ( .A(Q_int2), .Y(n4) );
endmodule


module uart_error_0 ( RST, CLK, RBUF_FULL, CHK_ERROR, OE );
  input RST, CLK, RBUF_FULL, CHK_ERROR;
  output OE;
  wire   OE_prime, n1;

  DFFSR OE_reg ( .D(OE_prime), .CLK(CLK), .R(n1), .S(1'b1), .Q(OE) );
  AND2X2 U5 ( .A(RBUF_FULL), .B(CHK_ERROR), .Y(OE_prime) );
  INVX2 U3 ( .A(RST), .Y(n1) );
endmodule


module uart_rcu_0 ( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT, RBUF_LOAD, 
        TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR );
  input CLK, RST, START_BIT, STOP_RCVING, SB_DETECT;
  output RBUF_LOAD, TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR;
  wire   timerRunning, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N99, \add_46/carry[6] , \add_46/carry[5] ,
         \add_46/carry[4] , \add_46/carry[3] , n3, n4, n5, n6, n7, n25, n32,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115;
  wire   [2:0] state;
  wire   [7:0] count;
  wire   [7:0] nextCount;
  wire   [2:0] nextState;

  DFFSR \count_reg[0]  ( .D(nextCount[0]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[0]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(n43), .CLK(CLK), .R(n4), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[0]) );
  DFFSR SBC_CLR_reg ( .D(n85), .CLK(CLK), .R(n4), .S(1'b1), .Q(SBC_CLR) );
  DFFSR TIMER_TRIG_reg ( .D(n84), .CLK(CLK), .R(n4), .S(1'b1), .Q(TIMER_TRIG)
         );
  DFFSR RBUF_LOAD_reg ( .D(n83), .CLK(CLK), .R(n4), .S(1'b1), .Q(RBUF_LOAD) );
  DFFSR timerRunning_reg ( .D(n89), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        timerRunning) );
  DFFSR \nextCount_reg[1]  ( .D(N32), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        nextCount[1]) );
  DFFSR \count_reg[1]  ( .D(nextCount[1]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        count[1]) );
  DFFSR \nextCount_reg[0]  ( .D(N31), .CLK(CLK), .R(1'b1), .S(n5), .Q(
        nextCount[0]) );
  DFFSR \nextCount_reg[2]  ( .D(N33), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        nextCount[2]) );
  DFFSR \count_reg[2]  ( .D(nextCount[2]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[2]) );
  DFFSR \nextCount_reg[3]  ( .D(N34), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[3]) );
  DFFSR \count_reg[3]  ( .D(nextCount[3]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[3]) );
  DFFSR \nextCount_reg[4]  ( .D(N35), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[4]) );
  DFFSR \count_reg[4]  ( .D(nextCount[4]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[4]) );
  DFFSR \nextCount_reg[5]  ( .D(N36), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[5]) );
  DFFSR \count_reg[5]  ( .D(nextCount[5]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[5]) );
  DFFSR \nextCount_reg[6]  ( .D(N37), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[6]) );
  DFFSR \count_reg[6]  ( .D(nextCount[6]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[6]) );
  DFFSR \nextCount_reg[7]  ( .D(N38), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        nextCount[7]) );
  DFFSR \count_reg[7]  ( .D(nextCount[7]), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        count[7]) );
  DFFSR SBC_EN_reg ( .D(n87), .CLK(CLK), .R(n4), .S(1'b1), .Q(SBC_EN) );
  AND2X2 U33 ( .A(N30), .B(timerRunning), .Y(N38) );
  AND2X2 U34 ( .A(N29), .B(timerRunning), .Y(N37) );
  AND2X2 U35 ( .A(N28), .B(timerRunning), .Y(N36) );
  AND2X2 U36 ( .A(N27), .B(timerRunning), .Y(N35) );
  AND2X2 U37 ( .A(N26), .B(timerRunning), .Y(N34) );
  AND2X2 U38 ( .A(N25), .B(timerRunning), .Y(N33) );
  AND2X2 U39 ( .A(N24), .B(timerRunning), .Y(N32) );
  OAI21X1 U54 ( .A(n114), .B(n45), .C(n113), .Y(n115) );
  OAI21X1 U55 ( .A(n46), .B(n44), .C(n45), .Y(n113) );
  NAND2X1 U56 ( .A(n112), .B(n111), .Y(n89) );
  OAI21X1 U57 ( .A(n110), .B(n109), .C(timerRunning), .Y(n111) );
  NAND2X1 U58 ( .A(n108), .B(n107), .Y(n109) );
  NAND2X1 U59 ( .A(n106), .B(n107), .Y(n88) );
  NAND3X1 U60 ( .A(n37), .B(n112), .C(CHK_ERROR), .Y(n106) );
  OAI21X1 U61 ( .A(n105), .B(n82), .C(n104), .Y(n87) );
  NAND2X1 U62 ( .A(n107), .B(n103), .Y(n105) );
  NAND2X1 U63 ( .A(n102), .B(n40), .Y(n107) );
  NAND3X1 U64 ( .A(n101), .B(n100), .C(n99), .Y(n86) );
  NAND3X1 U65 ( .A(n36), .B(n112), .C(SET_RBUF_FULL), .Y(n99) );
  NAND2X1 U66 ( .A(n103), .B(n100), .Y(n110) );
  NAND3X1 U67 ( .A(nextState[0]), .B(nextState[1]), .C(n102), .Y(n100) );
  NAND3X1 U68 ( .A(n38), .B(n40), .C(n102), .Y(n101) );
  OAI21X1 U69 ( .A(n98), .B(n47), .C(n112), .Y(n85) );
  OAI21X1 U70 ( .A(n98), .B(n81), .C(n112), .Y(n84) );
  NAND2X1 U71 ( .A(n103), .B(n104), .Y(n98) );
  NAND3X1 U72 ( .A(nextState[1]), .B(n38), .C(n41), .Y(n104) );
  NAND2X1 U73 ( .A(n97), .B(n108), .Y(n83) );
  NAND3X1 U74 ( .A(nextState[1]), .B(n38), .C(n102), .Y(n108) );
  NAND3X1 U75 ( .A(n103), .B(n112), .C(RBUF_LOAD), .Y(n97) );
  NAND3X1 U76 ( .A(nextState[0]), .B(n40), .C(n41), .Y(n112) );
  NAND3X1 U77 ( .A(n38), .B(n40), .C(n41), .Y(n103) );
  OAI21X1 U78 ( .A(n42), .B(n45), .C(n96), .Y(n102) );
  NAND3X1 U79 ( .A(state[0]), .B(n45), .C(state[1]), .Y(n96) );
  NAND2X1 U80 ( .A(n95), .B(n94), .Y(n114) );
  OAI21X1 U81 ( .A(n93), .B(n94), .C(n95), .Y(nextState[1]) );
  NOR2X1 U82 ( .A(N99), .B(state[2]), .Y(n93) );
  OAI21X1 U83 ( .A(state[2]), .B(n92), .C(n95), .Y(nextState[0]) );
  NAND2X1 U84 ( .A(state[1]), .B(n46), .Y(n95) );
  AOI21X1 U85 ( .A(START_BIT), .B(n46), .C(n91), .Y(n92) );
  OAI21X1 U86 ( .A(N99), .B(n94), .C(n90), .Y(n91) );
  NAND2X1 U87 ( .A(SB_DETECT), .B(state[1]), .Y(n90) );
  NAND2X1 U88 ( .A(state[0]), .B(n44), .Y(n94) );
  NAND2X1 U89 ( .A(n39), .B(timerRunning), .Y(N31) );
  DFFSR SET_RBUF_FULL_reg ( .D(n86), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        SET_RBUF_FULL) );
  DFFSR CHK_ERROR_reg ( .D(n88), .CLK(CLK), .R(n4), .S(1'b1), .Q(CHK_ERROR) );
  INVX2 U7 ( .A(RST), .Y(n4) );
  INVX2 U8 ( .A(RST), .Y(n5) );
  XNOR2X1 U24 ( .A(count[7]), .B(n3), .Y(N30) );
  NAND2X1 U31 ( .A(count[6]), .B(\add_46/carry[6] ), .Y(n3) );
  XOR2X1 U40 ( .A(\add_46/carry[6] ), .B(count[6]), .Y(N29) );
  AND2X1 U41 ( .A(count[5]), .B(\add_46/carry[5] ), .Y(\add_46/carry[6] ) );
  XOR2X1 U42 ( .A(\add_46/carry[5] ), .B(count[5]), .Y(N28) );
  AND2X1 U43 ( .A(count[4]), .B(\add_46/carry[4] ), .Y(\add_46/carry[5] ) );
  XOR2X1 U44 ( .A(\add_46/carry[4] ), .B(count[4]), .Y(N27) );
  AND2X1 U45 ( .A(count[3]), .B(\add_46/carry[3] ), .Y(\add_46/carry[4] ) );
  XOR2X1 U46 ( .A(\add_46/carry[3] ), .B(count[3]), .Y(N26) );
  AND2X1 U47 ( .A(count[2]), .B(count[1]), .Y(\add_46/carry[3] ) );
  XOR2X1 U48 ( .A(count[1]), .B(count[2]), .Y(N25) );
  INVX2 U49 ( .A(count[1]), .Y(N24) );
  OAI21X1 U50 ( .A(count[0]), .B(count[1]), .C(count[2]), .Y(n6) );
  NOR2X1 U51 ( .A(n35), .B(n6), .Y(n7) );
  OAI21X1 U52 ( .A(n7), .B(count[4]), .C(count[6]), .Y(n25) );
  OAI21X1 U53 ( .A(n34), .B(n25), .C(n32), .Y(N99) );
  INVX2 U90 ( .A(count[7]), .Y(n32) );
  INVX2 U91 ( .A(count[5]), .Y(n34) );
  INVX2 U92 ( .A(count[3]), .Y(n35) );
  INVX2 U93 ( .A(n110), .Y(n36) );
  INVX2 U94 ( .A(n105), .Y(n37) );
  INVX2 U95 ( .A(nextState[0]), .Y(n38) );
  INVX2 U96 ( .A(count[0]), .Y(n39) );
  INVX2 U97 ( .A(nextState[1]), .Y(n40) );
  INVX2 U98 ( .A(n102), .Y(n41) );
  INVX2 U99 ( .A(n114), .Y(n42) );
  INVX2 U100 ( .A(n115), .Y(n43) );
  INVX2 U101 ( .A(state[1]), .Y(n44) );
  INVX2 U102 ( .A(state[2]), .Y(n45) );
  INVX2 U103 ( .A(state[0]), .Y(n46) );
  INVX2 U104 ( .A(SBC_CLR), .Y(n47) );
  INVX2 U105 ( .A(TIMER_TRIG), .Y(n81) );
  INVX2 U106 ( .A(SBC_EN), .Y(n82) );
endmodule


module uart_rcv_buf_0 ( CLK, RST, LOAD_RBUF, LOAD_DATA, RCV_DATA );
  input [7:0] LOAD_DATA;
  output [7:0] RCV_DATA;
  input CLK, RST, LOAD_RBUF;
  wire   n11, n12, n13, n15, n17, n19, n21, n23, n24, n26, n34, n35, n36, n37,
         n38, n39, n40, n41;

  DFFSR \Q_int_reg[7]  ( .D(n12), .CLK(CLK), .R(n11), .S(1'b1), .Q(RCV_DATA[7]) );
  DFFSR \Q_int_reg[6]  ( .D(n13), .CLK(CLK), .R(n11), .S(1'b1), .Q(RCV_DATA[6]) );
  DFFSR \Q_int_reg[5]  ( .D(n15), .CLK(CLK), .R(n11), .S(1'b1), .Q(RCV_DATA[5]) );
  DFFSR \Q_int_reg[4]  ( .D(n17), .CLK(CLK), .R(n11), .S(1'b1), .Q(RCV_DATA[4]) );
  DFFSR \Q_int_reg[3]  ( .D(n19), .CLK(CLK), .R(n11), .S(1'b1), .Q(RCV_DATA[3]) );
  DFFSR \Q_int_reg[2]  ( .D(n21), .CLK(CLK), .R(n11), .S(1'b1), .Q(RCV_DATA[2]) );
  DFFSR \Q_int_reg[0]  ( .D(n24), .CLK(CLK), .R(n11), .S(1'b1), .Q(RCV_DATA[0]) );
  AOI22X1 U3 ( .A(LOAD_RBUF), .B(LOAD_DATA[0]), .C(RCV_DATA[0]), .D(n26), .Y(
        n41) );
  AOI22X1 U5 ( .A(LOAD_DATA[1]), .B(LOAD_RBUF), .C(RCV_DATA[1]), .D(n26), .Y(
        n40) );
  AOI22X1 U7 ( .A(LOAD_DATA[2]), .B(LOAD_RBUF), .C(RCV_DATA[2]), .D(n26), .Y(
        n39) );
  AOI22X1 U9 ( .A(LOAD_DATA[3]), .B(LOAD_RBUF), .C(RCV_DATA[3]), .D(n26), .Y(
        n38) );
  AOI22X1 U11 ( .A(LOAD_DATA[4]), .B(LOAD_RBUF), .C(RCV_DATA[4]), .D(n26), .Y(
        n37) );
  AOI22X1 U13 ( .A(LOAD_DATA[5]), .B(LOAD_RBUF), .C(RCV_DATA[5]), .D(n26), .Y(
        n36) );
  AOI22X1 U15 ( .A(LOAD_DATA[6]), .B(LOAD_RBUF), .C(RCV_DATA[6]), .D(n26), .Y(
        n35) );
  AOI22X1 U18 ( .A(LOAD_DATA[7]), .B(LOAD_RBUF), .C(RCV_DATA[7]), .D(n26), .Y(
        n34) );
  DFFSR \Q_int_reg[1]  ( .D(n23), .CLK(CLK), .R(n11), .S(1'b1), .Q(RCV_DATA[1]) );
  INVX2 U4 ( .A(RST), .Y(n11) );
  INVX2 U6 ( .A(n34), .Y(n12) );
  INVX2 U8 ( .A(n35), .Y(n13) );
  INVX2 U10 ( .A(n36), .Y(n15) );
  INVX2 U12 ( .A(n37), .Y(n17) );
  INVX2 U14 ( .A(n38), .Y(n19) );
  INVX2 U16 ( .A(n39), .Y(n21) );
  INVX2 U17 ( .A(n40), .Y(n23) );
  INVX2 U19 ( .A(n41), .Y(n24) );
  INVX2 U21 ( .A(LOAD_RBUF), .Y(n26) );
endmodule


module uart_rcv_buf_full_0 ( CLK, RST, CLR_RBUF, SET_RBUF_FULL, RBUF_FULL );
  input CLK, RST, CLR_RBUF, SET_RBUF_FULL;
  output RBUF_FULL;
  wire   n4, n6;

  DFFSR Q_int_reg ( .D(n4), .CLK(CLK), .R(n6), .S(1'b1), .Q(RBUF_FULL) );
  NOR2X1 U3 ( .A(RST), .B(CLR_RBUF), .Y(n6) );
  OR2X2 U4 ( .A(RBUF_FULL), .B(SET_RBUF_FULL), .Y(n4) );
endmodule


module uart_sb_check_0 ( RST, CLK, SBC_CLR, SBC_EN, STOP_DATA, SB_DETECT, SBE
 );
  input [1:0] STOP_DATA;
  input RST, CLK, SBC_CLR, SBC_EN;
  output SB_DETECT, SBE;
  wire   SBE_prime, sb_detect_flag, n2, n4, n5, n6, n10, n11, n12;

  DFFSR SB_DETECT_reg ( .D(sb_detect_flag), .CLK(CLK), .R(n2), .S(1'b1), .Q(
        SB_DETECT) );
  DFFSR SBE_reg ( .D(SBE_prime), .CLK(CLK), .R(n2), .S(1'b1), .Q(SBE) );
  OR2X2 U6 ( .A(SBC_CLR), .B(STOP_DATA[0]), .Y(n12) );
  NOR2X1 U10 ( .A(n12), .B(n11), .Y(sb_detect_flag) );
  NAND2X1 U11 ( .A(STOP_DATA[1]), .B(SBC_EN), .Y(n11) );
  NOR2X1 U12 ( .A(n6), .B(n10), .Y(SBE_prime) );
  OAI21X1 U13 ( .A(STOP_DATA[0]), .B(n4), .C(n5), .Y(n10) );
  INVX2 U4 ( .A(RST), .Y(n2) );
  INVX2 U7 ( .A(STOP_DATA[1]), .Y(n4) );
  INVX2 U8 ( .A(SBC_CLR), .Y(n5) );
  INVX2 U9 ( .A(SBC_EN), .Y(n6) );
endmodule


module uart_sr_10bit_0 ( CLK, RST, SHIFT_STROBE, SERIAL_IN, LOAD_DATA, 
        STOP_DATA );
  output [7:0] LOAD_DATA;
  output [1:0] STOP_DATA;
  input CLK, RST, SHIFT_STROBE, SERIAL_IN;
  wire   n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, n34, n35, n36,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48;

  DFFSR \present_val_reg[9]  ( .D(n36), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        STOP_DATA[1]) );
  OAI21X1 U2 ( .A(n35), .B(n17), .C(n48), .Y(n46) );
  NAND2X1 U3 ( .A(LOAD_DATA[0]), .B(n17), .Y(n48) );
  OAI22X1 U4 ( .A(n17), .B(n34), .C(n13), .D(n35), .Y(n45) );
  OAI22X1 U6 ( .A(n17), .B(n31), .C(n13), .D(n34), .Y(n44) );
  OAI22X1 U8 ( .A(n17), .B(n29), .C(n13), .D(n31), .Y(n43) );
  OAI22X1 U10 ( .A(n17), .B(n27), .C(n13), .D(n29), .Y(n42) );
  OAI22X1 U12 ( .A(n17), .B(n25), .C(n13), .D(n27), .Y(n41) );
  OAI22X1 U14 ( .A(n17), .B(n23), .C(n13), .D(n25), .Y(n40) );
  OAI22X1 U16 ( .A(n17), .B(n21), .C(n13), .D(n23), .Y(n39) );
  OAI22X1 U18 ( .A(n17), .B(n19), .C(n13), .D(n21), .Y(n38) );
  OAI21X1 U22 ( .A(n13), .B(n19), .C(n47), .Y(n36) );
  NAND2X1 U23 ( .A(SERIAL_IN), .B(n13), .Y(n47) );
  DFFSR \present_val_reg[8]  ( .D(n38), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        STOP_DATA[0]) );
  DFFSR \present_val_reg[7]  ( .D(n39), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[7]) );
  DFFSR \present_val_reg[6]  ( .D(n40), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[6]) );
  DFFSR \present_val_reg[5]  ( .D(n41), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[5]) );
  DFFSR \present_val_reg[4]  ( .D(n42), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[4]) );
  DFFSR \present_val_reg[3]  ( .D(n43), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[3]) );
  DFFSR \present_val_reg[2]  ( .D(n44), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[2]) );
  DFFSR \present_val_reg[1]  ( .D(n45), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[1]) );
  DFFSR \present_val_reg[0]  ( .D(n46), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[0]) );
  INVX2 U21 ( .A(RST), .Y(n15) );
  INVX2 U24 ( .A(n13), .Y(n17) );
  INVX4 U25 ( .A(n11), .Y(n13) );
  INVX2 U26 ( .A(SHIFT_STROBE), .Y(n11) );
  INVX2 U27 ( .A(STOP_DATA[1]), .Y(n19) );
  INVX2 U28 ( .A(STOP_DATA[0]), .Y(n21) );
  INVX2 U29 ( .A(LOAD_DATA[7]), .Y(n23) );
  INVX2 U30 ( .A(LOAD_DATA[6]), .Y(n25) );
  INVX2 U31 ( .A(LOAD_DATA[5]), .Y(n27) );
  INVX2 U32 ( .A(LOAD_DATA[4]), .Y(n29) );
  INVX2 U33 ( .A(LOAD_DATA[3]), .Y(n31) );
  INVX2 U35 ( .A(LOAD_DATA[2]), .Y(n34) );
  INVX2 U36 ( .A(LOAD_DATA[1]), .Y(n35) );
endmodule


module keyreg_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  AND2X2 U2 ( .A(n21), .B(n17), .Y(n1) );
  XNOR2X1 U3 ( .A(n32), .B(n33), .Y(SUM[3]) );
  XOR2X1 U4 ( .A(n27), .B(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n31), .B(n30), .Y(n2) );
  NAND2X1 U6 ( .A(n35), .B(n36), .Y(n22) );
  INVX2 U7 ( .A(n41), .Y(SUM[0]) );
  XNOR2X1 U8 ( .A(n3), .B(n4), .Y(SUM[7]) );
  XOR2X1 U9 ( .A(B[7]), .B(A[7]), .Y(n4) );
  AOI21X1 U10 ( .A(n5), .B(n6), .C(n7), .Y(n3) );
  NAND2X1 U11 ( .A(n8), .B(n9), .Y(n7) );
  NAND2X1 U12 ( .A(n10), .B(n11), .Y(n8) );
  AND2X2 U13 ( .A(n12), .B(n11), .Y(n5) );
  XNOR2X1 U14 ( .A(n13), .B(n14), .Y(SUM[6]) );
  AND2X2 U15 ( .A(n11), .B(n9), .Y(n14) );
  NAND2X1 U16 ( .A(B[6]), .B(A[6]), .Y(n9) );
  OR2X2 U17 ( .A(A[6]), .B(B[6]), .Y(n11) );
  AOI21X1 U18 ( .A(n6), .B(n12), .C(n10), .Y(n13) );
  INVX2 U19 ( .A(n15), .Y(n10) );
  XNOR2X1 U20 ( .A(n6), .B(n16), .Y(SUM[5]) );
  NAND2X1 U21 ( .A(n12), .B(n15), .Y(n16) );
  NAND2X1 U22 ( .A(B[5]), .B(A[5]), .Y(n15) );
  OR2X2 U23 ( .A(A[5]), .B(B[5]), .Y(n12) );
  NAND3X1 U24 ( .A(n17), .B(n18), .C(n19), .Y(n6) );
  NAND3X1 U25 ( .A(n20), .B(n21), .C(n22), .Y(n19) );
  INVX2 U26 ( .A(n23), .Y(n20) );
  NAND3X1 U27 ( .A(n24), .B(n21), .C(n25), .Y(n18) );
  XOR2X1 U28 ( .A(n26), .B(n1), .Y(SUM[4]) );
  NAND2X1 U29 ( .A(B[4]), .B(A[4]), .Y(n17) );
  OR2X2 U30 ( .A(A[4]), .B(B[4]), .Y(n21) );
  OAI21X1 U31 ( .A(n27), .B(n23), .C(n28), .Y(n26) );
  NAND2X1 U32 ( .A(n24), .B(n25), .Y(n28) );
  NAND2X1 U33 ( .A(n29), .B(n30), .Y(n25) );
  NAND2X1 U34 ( .A(n31), .B(n24), .Y(n23) );
  NAND2X1 U35 ( .A(n24), .B(n29), .Y(n33) );
  NAND2X1 U36 ( .A(B[3]), .B(A[3]), .Y(n29) );
  OR2X2 U37 ( .A(A[3]), .B(B[3]), .Y(n24) );
  NAND2X1 U38 ( .A(n30), .B(n34), .Y(n32) );
  NAND2X1 U39 ( .A(n22), .B(n31), .Y(n34) );
  NAND2X1 U40 ( .A(B[2]), .B(A[2]), .Y(n30) );
  OR2X2 U41 ( .A(A[2]), .B(B[2]), .Y(n31) );
  INVX2 U42 ( .A(n22), .Y(n27) );
  NAND2X1 U43 ( .A(n38), .B(n37), .Y(n35) );
  AND2X2 U44 ( .A(A[0]), .B(B[0]), .Y(n38) );
  XOR2X1 U45 ( .A(n39), .B(n40), .Y(SUM[1]) );
  NAND2X1 U46 ( .A(n37), .B(n36), .Y(n39) );
  NAND2X1 U47 ( .A(B[1]), .B(A[1]), .Y(n36) );
  OR2X2 U48 ( .A(A[1]), .B(B[1]), .Y(n37) );
  OAI21X1 U49 ( .A(A[0]), .B(B[0]), .C(n40), .Y(n41) );
  NAND2X1 U50 ( .A(B[0]), .B(A[0]), .Y(n40) );
endmodule


module keyreg_0 ( CLK, RST, SBE, OE, RBUF_FULL, RCV_DATA, PLAINKEY, KEY_ERROR, 
        PROG_ERROR, CLR_RBUFF, PARITY_ERROR );
  input [7:0] RCV_DATA;
  output [63:0] PLAINKEY;
  input CLK, RST, SBE, OE, RBUF_FULL;
  output KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR;
  wire   parityError, nextParityError, N1792, N1793, N1794, N1795, N1796,
         N1797, N1798, N1799, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n14,
         n16, n17, n19, n20, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39,
         n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63, n65, n67,
         n69, n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95,
         n97, n99, n101, n103, n105, n107, n109, n111, n113, n115, n117, n119,
         n121, n123, n125, n127, n129, n131, n133, n135, n137, n139, n141,
         n143, n145, n147, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1267, n1268, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988;
  wire   [3:0] state;
  wire   [3:0] keyCount;
  wire   [7:0] address;
  wire   [63:0] currentPlainKey;
  wire   [7:0] parityAccumulator;

  DFFPOSX1 \keyCount_reg[0]  ( .D(n1762), .CLK(CLK), .Q(keyCount[0]) );
  DFFPOSX1 \keyCount_reg[2]  ( .D(n1769), .CLK(CLK), .Q(keyCount[2]) );
  DFFPOSX1 \keyCount_reg[3]  ( .D(n1763), .CLK(CLK), .Q(keyCount[3]) );
  DFFSR \state_reg[0]  ( .D(n1765), .CLK(CLK), .R(n293), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[1]  ( .D(n1767), .CLK(CLK), .R(n290), .S(1'b1), .Q(state[1]) );
  DFFSR \state_reg[2]  ( .D(n1766), .CLK(CLK), .R(n292), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[3]  ( .D(n1764), .CLK(CLK), .R(n291), .S(1'b1), .Q(state[3]) );
  DFFPOSX1 \parityAccumulator_reg[0]  ( .D(n1770), .CLK(CLK), .Q(
        parityAccumulator[0]) );
  DFFPOSX1 \parityAccumulator_reg[1]  ( .D(n1771), .CLK(CLK), .Q(
        parityAccumulator[1]) );
  DFFPOSX1 \parityAccumulator_reg[2]  ( .D(n1772), .CLK(CLK), .Q(
        parityAccumulator[2]) );
  DFFPOSX1 \parityAccumulator_reg[3]  ( .D(n1773), .CLK(CLK), .Q(
        parityAccumulator[3]) );
  DFFPOSX1 \parityAccumulator_reg[4]  ( .D(n1774), .CLK(CLK), .Q(
        parityAccumulator[4]) );
  DFFPOSX1 \parityAccumulator_reg[5]  ( .D(n1775), .CLK(CLK), .Q(
        parityAccumulator[5]) );
  DFFPOSX1 \parityAccumulator_reg[6]  ( .D(n1776), .CLK(CLK), .Q(
        parityAccumulator[6]) );
  DFFPOSX1 \parityAccumulator_reg[7]  ( .D(n1777), .CLK(CLK), .Q(
        parityAccumulator[7]) );
  DFFPOSX1 \keyCount_reg[1]  ( .D(n1768), .CLK(CLK), .Q(keyCount[1]) );
  DFFSR PARITY_ERROR_reg ( .D(nextParityError), .CLK(CLK), .R(n292), .S(1'b1), 
        .Q(PARITY_ERROR) );
  DFFSR parityError_reg ( .D(nextParityError), .CLK(CLK), .R(n292), .S(1'b1), 
        .Q(parityError) );
  DFFPOSX1 \address_reg[7]  ( .D(n1778), .CLK(CLK), .Q(address[7]) );
  DFFPOSX1 \address_reg[6]  ( .D(n1779), .CLK(CLK), .Q(address[6]) );
  DFFPOSX1 \address_reg[5]  ( .D(n1780), .CLK(CLK), .Q(address[5]) );
  DFFPOSX1 \address_reg[4]  ( .D(n1781), .CLK(CLK), .Q(address[4]) );
  DFFPOSX1 \address_reg[3]  ( .D(n1782), .CLK(CLK), .Q(address[3]) );
  DFFPOSX1 \address_reg[2]  ( .D(n1783), .CLK(CLK), .Q(address[2]) );
  DFFPOSX1 \address_reg[1]  ( .D(n1784), .CLK(CLK), .Q(address[1]) );
  DFFPOSX1 \address_reg[0]  ( .D(n1785), .CLK(CLK), .Q(address[0]) );
  DFFPOSX1 \currentPlainKey_reg[63]  ( .D(n1849), .CLK(CLK), .Q(
        currentPlainKey[63]) );
  DFFPOSX1 \currentPlainKey_reg[62]  ( .D(n1848), .CLK(CLK), .Q(
        currentPlainKey[62]) );
  DFFPOSX1 \currentPlainKey_reg[61]  ( .D(n1847), .CLK(CLK), .Q(
        currentPlainKey[61]) );
  DFFPOSX1 \currentPlainKey_reg[60]  ( .D(n1846), .CLK(CLK), .Q(
        currentPlainKey[60]) );
  DFFPOSX1 \currentPlainKey_reg[59]  ( .D(n1845), .CLK(CLK), .Q(
        currentPlainKey[59]) );
  DFFPOSX1 \currentPlainKey_reg[58]  ( .D(n1844), .CLK(CLK), .Q(
        currentPlainKey[58]) );
  DFFPOSX1 \currentPlainKey_reg[57]  ( .D(n1843), .CLK(CLK), .Q(
        currentPlainKey[57]) );
  DFFPOSX1 \currentPlainKey_reg[56]  ( .D(n1842), .CLK(CLK), .Q(
        currentPlainKey[56]) );
  DFFPOSX1 \currentPlainKey_reg[55]  ( .D(n1841), .CLK(CLK), .Q(
        currentPlainKey[55]) );
  DFFPOSX1 \currentPlainKey_reg[54]  ( .D(n1840), .CLK(CLK), .Q(
        currentPlainKey[54]) );
  DFFPOSX1 \currentPlainKey_reg[53]  ( .D(n1839), .CLK(CLK), .Q(
        currentPlainKey[53]) );
  DFFPOSX1 \currentPlainKey_reg[52]  ( .D(n1838), .CLK(CLK), .Q(
        currentPlainKey[52]) );
  DFFPOSX1 \currentPlainKey_reg[51]  ( .D(n1837), .CLK(CLK), .Q(
        currentPlainKey[51]) );
  DFFPOSX1 \currentPlainKey_reg[50]  ( .D(n1836), .CLK(CLK), .Q(
        currentPlainKey[50]) );
  DFFPOSX1 \currentPlainKey_reg[49]  ( .D(n1835), .CLK(CLK), .Q(
        currentPlainKey[49]) );
  DFFPOSX1 \currentPlainKey_reg[48]  ( .D(n1834), .CLK(CLK), .Q(
        currentPlainKey[48]) );
  DFFPOSX1 \currentPlainKey_reg[47]  ( .D(n1833), .CLK(CLK), .Q(
        currentPlainKey[47]) );
  DFFPOSX1 \currentPlainKey_reg[46]  ( .D(n1832), .CLK(CLK), .Q(
        currentPlainKey[46]) );
  DFFPOSX1 \currentPlainKey_reg[45]  ( .D(n1831), .CLK(CLK), .Q(
        currentPlainKey[45]) );
  DFFPOSX1 \currentPlainKey_reg[44]  ( .D(n1830), .CLK(CLK), .Q(
        currentPlainKey[44]) );
  DFFPOSX1 \currentPlainKey_reg[43]  ( .D(n1829), .CLK(CLK), .Q(
        currentPlainKey[43]) );
  DFFPOSX1 \currentPlainKey_reg[42]  ( .D(n1828), .CLK(CLK), .Q(
        currentPlainKey[42]) );
  DFFPOSX1 \currentPlainKey_reg[41]  ( .D(n1827), .CLK(CLK), .Q(
        currentPlainKey[41]) );
  DFFPOSX1 \currentPlainKey_reg[40]  ( .D(n1826), .CLK(CLK), .Q(
        currentPlainKey[40]) );
  DFFPOSX1 \currentPlainKey_reg[39]  ( .D(n1825), .CLK(CLK), .Q(
        currentPlainKey[39]) );
  DFFPOSX1 \currentPlainKey_reg[38]  ( .D(n1824), .CLK(CLK), .Q(
        currentPlainKey[38]) );
  DFFPOSX1 \currentPlainKey_reg[37]  ( .D(n1823), .CLK(CLK), .Q(
        currentPlainKey[37]) );
  DFFPOSX1 \currentPlainKey_reg[36]  ( .D(n1822), .CLK(CLK), .Q(
        currentPlainKey[36]) );
  DFFPOSX1 \currentPlainKey_reg[35]  ( .D(n1821), .CLK(CLK), .Q(
        currentPlainKey[35]) );
  DFFPOSX1 \currentPlainKey_reg[34]  ( .D(n1820), .CLK(CLK), .Q(
        currentPlainKey[34]) );
  DFFPOSX1 \currentPlainKey_reg[33]  ( .D(n1819), .CLK(CLK), .Q(
        currentPlainKey[33]) );
  DFFPOSX1 \currentPlainKey_reg[32]  ( .D(n1818), .CLK(CLK), .Q(
        currentPlainKey[32]) );
  DFFPOSX1 \currentPlainKey_reg[31]  ( .D(n1817), .CLK(CLK), .Q(
        currentPlainKey[31]) );
  DFFPOSX1 \currentPlainKey_reg[30]  ( .D(n1816), .CLK(CLK), .Q(
        currentPlainKey[30]) );
  DFFPOSX1 \currentPlainKey_reg[29]  ( .D(n1815), .CLK(CLK), .Q(
        currentPlainKey[29]) );
  DFFPOSX1 \currentPlainKey_reg[28]  ( .D(n1814), .CLK(CLK), .Q(
        currentPlainKey[28]) );
  DFFPOSX1 \currentPlainKey_reg[27]  ( .D(n1813), .CLK(CLK), .Q(
        currentPlainKey[27]) );
  DFFPOSX1 \currentPlainKey_reg[26]  ( .D(n1812), .CLK(CLK), .Q(
        currentPlainKey[26]) );
  DFFPOSX1 \currentPlainKey_reg[25]  ( .D(n1811), .CLK(CLK), .Q(
        currentPlainKey[25]) );
  DFFPOSX1 \currentPlainKey_reg[24]  ( .D(n1810), .CLK(CLK), .Q(
        currentPlainKey[24]) );
  DFFPOSX1 \currentPlainKey_reg[23]  ( .D(n1809), .CLK(CLK), .Q(
        currentPlainKey[23]) );
  DFFPOSX1 \currentPlainKey_reg[22]  ( .D(n1808), .CLK(CLK), .Q(
        currentPlainKey[22]) );
  DFFPOSX1 \currentPlainKey_reg[21]  ( .D(n1807), .CLK(CLK), .Q(
        currentPlainKey[21]) );
  DFFPOSX1 \currentPlainKey_reg[20]  ( .D(n1806), .CLK(CLK), .Q(
        currentPlainKey[20]) );
  DFFPOSX1 \currentPlainKey_reg[19]  ( .D(n1805), .CLK(CLK), .Q(
        currentPlainKey[19]) );
  DFFPOSX1 \currentPlainKey_reg[18]  ( .D(n1804), .CLK(CLK), .Q(
        currentPlainKey[18]) );
  DFFPOSX1 \currentPlainKey_reg[17]  ( .D(n1803), .CLK(CLK), .Q(
        currentPlainKey[17]) );
  DFFPOSX1 \currentPlainKey_reg[16]  ( .D(n1802), .CLK(CLK), .Q(
        currentPlainKey[16]) );
  DFFPOSX1 \currentPlainKey_reg[15]  ( .D(n1801), .CLK(CLK), .Q(
        currentPlainKey[15]) );
  DFFPOSX1 \currentPlainKey_reg[14]  ( .D(n1800), .CLK(CLK), .Q(
        currentPlainKey[14]) );
  DFFPOSX1 \currentPlainKey_reg[13]  ( .D(n1799), .CLK(CLK), .Q(
        currentPlainKey[13]) );
  DFFPOSX1 \currentPlainKey_reg[12]  ( .D(n1798), .CLK(CLK), .Q(
        currentPlainKey[12]) );
  DFFPOSX1 \currentPlainKey_reg[11]  ( .D(n1797), .CLK(CLK), .Q(
        currentPlainKey[11]) );
  DFFPOSX1 \currentPlainKey_reg[10]  ( .D(n1796), .CLK(CLK), .Q(
        currentPlainKey[10]) );
  DFFPOSX1 \currentPlainKey_reg[9]  ( .D(n1795), .CLK(CLK), .Q(
        currentPlainKey[9]) );
  DFFPOSX1 \currentPlainKey_reg[8]  ( .D(n1794), .CLK(CLK), .Q(
        currentPlainKey[8]) );
  DFFPOSX1 \currentPlainKey_reg[7]  ( .D(n1793), .CLK(CLK), .Q(
        currentPlainKey[7]) );
  DFFPOSX1 \currentPlainKey_reg[6]  ( .D(n1792), .CLK(CLK), .Q(
        currentPlainKey[6]) );
  DFFPOSX1 \currentPlainKey_reg[5]  ( .D(n1791), .CLK(CLK), .Q(
        currentPlainKey[5]) );
  DFFPOSX1 \currentPlainKey_reg[4]  ( .D(n1790), .CLK(CLK), .Q(
        currentPlainKey[4]) );
  DFFPOSX1 \currentPlainKey_reg[3]  ( .D(n1789), .CLK(CLK), .Q(
        currentPlainKey[3]) );
  DFFPOSX1 \currentPlainKey_reg[2]  ( .D(n1788), .CLK(CLK), .Q(
        currentPlainKey[2]) );
  DFFPOSX1 \currentPlainKey_reg[1]  ( .D(n1787), .CLK(CLK), .Q(
        currentPlainKey[1]) );
  DFFPOSX1 \currentPlainKey_reg[0]  ( .D(n1786), .CLK(CLK), .Q(
        currentPlainKey[0]) );
  DFFPOSX1 \PLAINKEY_reg[63]  ( .D(n1856), .CLK(CLK), .Q(PLAINKEY[63]) );
  DFFPOSX1 \PLAINKEY_reg[62]  ( .D(n1857), .CLK(CLK), .Q(PLAINKEY[62]) );
  DFFPOSX1 \PLAINKEY_reg[61]  ( .D(n1858), .CLK(CLK), .Q(PLAINKEY[61]) );
  DFFPOSX1 \PLAINKEY_reg[60]  ( .D(n1859), .CLK(CLK), .Q(PLAINKEY[60]) );
  DFFPOSX1 \PLAINKEY_reg[59]  ( .D(n1860), .CLK(CLK), .Q(PLAINKEY[59]) );
  DFFPOSX1 \PLAINKEY_reg[58]  ( .D(n1861), .CLK(CLK), .Q(PLAINKEY[58]) );
  DFFPOSX1 \PLAINKEY_reg[57]  ( .D(n1862), .CLK(CLK), .Q(PLAINKEY[57]) );
  DFFPOSX1 \PLAINKEY_reg[56]  ( .D(n1863), .CLK(CLK), .Q(PLAINKEY[56]) );
  DFFPOSX1 \PLAINKEY_reg[55]  ( .D(n1864), .CLK(CLK), .Q(PLAINKEY[55]) );
  DFFPOSX1 \PLAINKEY_reg[54]  ( .D(n1865), .CLK(CLK), .Q(PLAINKEY[54]) );
  DFFPOSX1 \PLAINKEY_reg[53]  ( .D(n1866), .CLK(CLK), .Q(PLAINKEY[53]) );
  DFFPOSX1 \PLAINKEY_reg[52]  ( .D(n1867), .CLK(CLK), .Q(PLAINKEY[52]) );
  DFFPOSX1 \PLAINKEY_reg[51]  ( .D(n1868), .CLK(CLK), .Q(PLAINKEY[51]) );
  DFFPOSX1 \PLAINKEY_reg[50]  ( .D(n1869), .CLK(CLK), .Q(PLAINKEY[50]) );
  DFFPOSX1 \PLAINKEY_reg[49]  ( .D(n1870), .CLK(CLK), .Q(PLAINKEY[49]) );
  DFFPOSX1 \PLAINKEY_reg[48]  ( .D(n1871), .CLK(CLK), .Q(PLAINKEY[48]) );
  DFFPOSX1 \PLAINKEY_reg[47]  ( .D(n1872), .CLK(CLK), .Q(PLAINKEY[47]) );
  DFFPOSX1 \PLAINKEY_reg[46]  ( .D(n1873), .CLK(CLK), .Q(PLAINKEY[46]) );
  DFFPOSX1 \PLAINKEY_reg[45]  ( .D(n1874), .CLK(CLK), .Q(PLAINKEY[45]) );
  DFFPOSX1 \PLAINKEY_reg[44]  ( .D(n1875), .CLK(CLK), .Q(PLAINKEY[44]) );
  DFFPOSX1 \PLAINKEY_reg[43]  ( .D(n1876), .CLK(CLK), .Q(PLAINKEY[43]) );
  DFFPOSX1 \PLAINKEY_reg[42]  ( .D(n1877), .CLK(CLK), .Q(PLAINKEY[42]) );
  DFFPOSX1 \PLAINKEY_reg[41]  ( .D(n1878), .CLK(CLK), .Q(PLAINKEY[41]) );
  DFFPOSX1 \PLAINKEY_reg[40]  ( .D(n1879), .CLK(CLK), .Q(PLAINKEY[40]) );
  DFFPOSX1 \PLAINKEY_reg[39]  ( .D(n1880), .CLK(CLK), .Q(PLAINKEY[39]) );
  DFFPOSX1 \PLAINKEY_reg[38]  ( .D(n1881), .CLK(CLK), .Q(PLAINKEY[38]) );
  DFFPOSX1 \PLAINKEY_reg[37]  ( .D(n1882), .CLK(CLK), .Q(PLAINKEY[37]) );
  DFFPOSX1 \PLAINKEY_reg[36]  ( .D(n1883), .CLK(CLK), .Q(PLAINKEY[36]) );
  DFFPOSX1 \PLAINKEY_reg[35]  ( .D(n1884), .CLK(CLK), .Q(PLAINKEY[35]) );
  DFFPOSX1 \PLAINKEY_reg[34]  ( .D(n1885), .CLK(CLK), .Q(PLAINKEY[34]) );
  DFFPOSX1 \PLAINKEY_reg[33]  ( .D(n1886), .CLK(CLK), .Q(PLAINKEY[33]) );
  DFFPOSX1 \PLAINKEY_reg[32]  ( .D(n1887), .CLK(CLK), .Q(PLAINKEY[32]) );
  DFFPOSX1 \PLAINKEY_reg[31]  ( .D(n1888), .CLK(CLK), .Q(PLAINKEY[31]) );
  DFFPOSX1 \PLAINKEY_reg[30]  ( .D(n1889), .CLK(CLK), .Q(PLAINKEY[30]) );
  DFFPOSX1 \PLAINKEY_reg[29]  ( .D(n1890), .CLK(CLK), .Q(PLAINKEY[29]) );
  DFFPOSX1 \PLAINKEY_reg[28]  ( .D(n1891), .CLK(CLK), .Q(PLAINKEY[28]) );
  DFFPOSX1 \PLAINKEY_reg[27]  ( .D(n1892), .CLK(CLK), .Q(PLAINKEY[27]) );
  DFFPOSX1 \PLAINKEY_reg[26]  ( .D(n1893), .CLK(CLK), .Q(PLAINKEY[26]) );
  DFFPOSX1 \PLAINKEY_reg[25]  ( .D(n1894), .CLK(CLK), .Q(PLAINKEY[25]) );
  DFFPOSX1 \PLAINKEY_reg[24]  ( .D(n1895), .CLK(CLK), .Q(PLAINKEY[24]) );
  DFFPOSX1 \PLAINKEY_reg[23]  ( .D(n1896), .CLK(CLK), .Q(PLAINKEY[23]) );
  DFFPOSX1 \PLAINKEY_reg[22]  ( .D(n1897), .CLK(CLK), .Q(PLAINKEY[22]) );
  DFFPOSX1 \PLAINKEY_reg[21]  ( .D(n1898), .CLK(CLK), .Q(PLAINKEY[21]) );
  DFFPOSX1 \PLAINKEY_reg[20]  ( .D(n1899), .CLK(CLK), .Q(PLAINKEY[20]) );
  DFFPOSX1 \PLAINKEY_reg[19]  ( .D(n1900), .CLK(CLK), .Q(PLAINKEY[19]) );
  DFFPOSX1 \PLAINKEY_reg[18]  ( .D(n1901), .CLK(CLK), .Q(PLAINKEY[18]) );
  DFFPOSX1 \PLAINKEY_reg[17]  ( .D(n1902), .CLK(CLK), .Q(PLAINKEY[17]) );
  DFFPOSX1 \PLAINKEY_reg[16]  ( .D(n1903), .CLK(CLK), .Q(PLAINKEY[16]) );
  DFFPOSX1 \PLAINKEY_reg[15]  ( .D(n1904), .CLK(CLK), .Q(PLAINKEY[15]) );
  DFFPOSX1 \PLAINKEY_reg[14]  ( .D(n1905), .CLK(CLK), .Q(PLAINKEY[14]) );
  DFFPOSX1 \PLAINKEY_reg[13]  ( .D(n1906), .CLK(CLK), .Q(PLAINKEY[13]) );
  DFFPOSX1 \PLAINKEY_reg[12]  ( .D(n1907), .CLK(CLK), .Q(PLAINKEY[12]) );
  DFFPOSX1 \PLAINKEY_reg[11]  ( .D(n1908), .CLK(CLK), .Q(PLAINKEY[11]) );
  DFFPOSX1 \PLAINKEY_reg[10]  ( .D(n1909), .CLK(CLK), .Q(PLAINKEY[10]) );
  DFFPOSX1 \PLAINKEY_reg[9]  ( .D(n1910), .CLK(CLK), .Q(PLAINKEY[9]) );
  DFFPOSX1 \PLAINKEY_reg[8]  ( .D(n1911), .CLK(CLK), .Q(PLAINKEY[8]) );
  DFFPOSX1 \PLAINKEY_reg[7]  ( .D(n1912), .CLK(CLK), .Q(PLAINKEY[7]) );
  DFFPOSX1 \PLAINKEY_reg[6]  ( .D(n1913), .CLK(CLK), .Q(PLAINKEY[6]) );
  DFFPOSX1 \PLAINKEY_reg[5]  ( .D(n1914), .CLK(CLK), .Q(PLAINKEY[5]) );
  DFFPOSX1 \PLAINKEY_reg[4]  ( .D(n1915), .CLK(CLK), .Q(PLAINKEY[4]) );
  DFFPOSX1 \PLAINKEY_reg[3]  ( .D(n1916), .CLK(CLK), .Q(PLAINKEY[3]) );
  DFFPOSX1 \PLAINKEY_reg[2]  ( .D(n1917), .CLK(CLK), .Q(PLAINKEY[2]) );
  DFFPOSX1 \PLAINKEY_reg[1]  ( .D(n1918), .CLK(CLK), .Q(PLAINKEY[1]) );
  DFFPOSX1 \PLAINKEY_reg[0]  ( .D(n1919), .CLK(CLK), .Q(PLAINKEY[0]) );
  NAND3X1 U9 ( .A(parityAccumulator[7]), .B(parityAccumulator[6]), .C(n1986), 
        .Y(n1987) );
  NOR2X1 U10 ( .A(n1692), .B(n1693), .Y(n1986) );
  NAND3X1 U11 ( .A(parityAccumulator[3]), .B(parityAccumulator[2]), .C(n1985), 
        .Y(n1988) );
  NOR2X1 U12 ( .A(n1688), .B(n1689), .Y(n1985) );
  OAI21X1 U13 ( .A(RST), .B(n1759), .C(n1984), .Y(n1919) );
  NAND2X1 U14 ( .A(PLAINKEY[0]), .B(n286), .Y(n1984) );
  OAI21X1 U15 ( .A(n284), .B(n1758), .C(n1983), .Y(n1918) );
  NAND2X1 U16 ( .A(PLAINKEY[1]), .B(n288), .Y(n1983) );
  OAI21X1 U17 ( .A(n285), .B(n1757), .C(n1982), .Y(n1917) );
  NAND2X1 U18 ( .A(PLAINKEY[2]), .B(n288), .Y(n1982) );
  OAI21X1 U19 ( .A(n287), .B(n1756), .C(n1981), .Y(n1916) );
  NAND2X1 U20 ( .A(PLAINKEY[3]), .B(n288), .Y(n1981) );
  OAI21X1 U21 ( .A(RST), .B(n1755), .C(n1980), .Y(n1915) );
  NAND2X1 U22 ( .A(PLAINKEY[4]), .B(n288), .Y(n1980) );
  OAI21X1 U24 ( .A(n286), .B(n1754), .C(n1979), .Y(n1914) );
  NAND2X1 U25 ( .A(PLAINKEY[5]), .B(n288), .Y(n1979) );
  OAI21X1 U27 ( .A(n284), .B(n1753), .C(n1978), .Y(n1913) );
  NAND2X1 U28 ( .A(PLAINKEY[6]), .B(n288), .Y(n1978) );
  OAI21X1 U30 ( .A(RST), .B(n1752), .C(n1977), .Y(n1912) );
  NAND2X1 U31 ( .A(PLAINKEY[7]), .B(n288), .Y(n1977) );
  OAI21X1 U33 ( .A(n288), .B(n1751), .C(n1976), .Y(n1911) );
  NAND2X1 U34 ( .A(PLAINKEY[8]), .B(n288), .Y(n1976) );
  OAI21X1 U36 ( .A(n284), .B(n1750), .C(n1975), .Y(n1910) );
  NAND2X1 U37 ( .A(PLAINKEY[9]), .B(n288), .Y(n1975) );
  OAI21X1 U39 ( .A(n284), .B(n1749), .C(n1974), .Y(n1909) );
  NAND2X1 U40 ( .A(PLAINKEY[10]), .B(n288), .Y(n1974) );
  OAI21X1 U42 ( .A(n284), .B(n1748), .C(n1973), .Y(n1908) );
  NAND2X1 U43 ( .A(PLAINKEY[11]), .B(n288), .Y(n1973) );
  OAI21X1 U45 ( .A(n284), .B(n1747), .C(n1972), .Y(n1907) );
  NAND2X1 U46 ( .A(PLAINKEY[12]), .B(n288), .Y(n1972) );
  OAI21X1 U48 ( .A(n284), .B(n1746), .C(n1971), .Y(n1906) );
  NAND2X1 U49 ( .A(PLAINKEY[13]), .B(n288), .Y(n1971) );
  OAI21X1 U51 ( .A(n284), .B(n1745), .C(n1970), .Y(n1905) );
  NAND2X1 U52 ( .A(PLAINKEY[14]), .B(n288), .Y(n1970) );
  OAI21X1 U54 ( .A(n284), .B(n1744), .C(n1969), .Y(n1904) );
  NAND2X1 U55 ( .A(PLAINKEY[15]), .B(n288), .Y(n1969) );
  OAI21X1 U57 ( .A(n285), .B(n1743), .C(n1968), .Y(n1903) );
  NAND2X1 U58 ( .A(PLAINKEY[16]), .B(n288), .Y(n1968) );
  OAI21X1 U60 ( .A(n285), .B(n1742), .C(n1967), .Y(n1902) );
  NAND2X1 U61 ( .A(PLAINKEY[17]), .B(n288), .Y(n1967) );
  OAI21X1 U63 ( .A(n285), .B(n1741), .C(n1966), .Y(n1901) );
  NAND2X1 U64 ( .A(PLAINKEY[18]), .B(n288), .Y(n1966) );
  OAI21X1 U66 ( .A(n285), .B(n1740), .C(n1965), .Y(n1900) );
  NAND2X1 U67 ( .A(PLAINKEY[19]), .B(n288), .Y(n1965) );
  OAI21X1 U69 ( .A(n285), .B(n1739), .C(n1964), .Y(n1899) );
  NAND2X1 U70 ( .A(PLAINKEY[20]), .B(n288), .Y(n1964) );
  OAI21X1 U72 ( .A(n285), .B(n1738), .C(n1963), .Y(n1898) );
  NAND2X1 U73 ( .A(PLAINKEY[21]), .B(n288), .Y(n1963) );
  OAI21X1 U75 ( .A(n285), .B(n1737), .C(n1962), .Y(n1897) );
  NAND2X1 U76 ( .A(PLAINKEY[22]), .B(n288), .Y(n1962) );
  OAI21X1 U78 ( .A(n286), .B(n1736), .C(n1961), .Y(n1896) );
  NAND2X1 U79 ( .A(PLAINKEY[23]), .B(n287), .Y(n1961) );
  OAI21X1 U81 ( .A(n285), .B(n1735), .C(n1960), .Y(n1895) );
  NAND2X1 U82 ( .A(PLAINKEY[24]), .B(n285), .Y(n1960) );
  OAI21X1 U84 ( .A(n284), .B(n1734), .C(n1959), .Y(n1894) );
  NAND2X1 U85 ( .A(PLAINKEY[25]), .B(n287), .Y(n1959) );
  OAI21X1 U87 ( .A(n286), .B(n1733), .C(n1958), .Y(n1893) );
  NAND2X1 U88 ( .A(PLAINKEY[26]), .B(n286), .Y(n1958) );
  OAI21X1 U90 ( .A(n286), .B(n1732), .C(n1957), .Y(n1892) );
  NAND2X1 U91 ( .A(PLAINKEY[27]), .B(n285), .Y(n1957) );
  OAI21X1 U93 ( .A(n285), .B(n1731), .C(n1956), .Y(n1891) );
  NAND2X1 U94 ( .A(PLAINKEY[28]), .B(n284), .Y(n1956) );
  OAI21X1 U96 ( .A(n286), .B(n1730), .C(n1955), .Y(n1890) );
  NAND2X1 U97 ( .A(PLAINKEY[29]), .B(n284), .Y(n1955) );
  OAI21X1 U99 ( .A(n286), .B(n1729), .C(n1954), .Y(n1889) );
  NAND2X1 U100 ( .A(PLAINKEY[30]), .B(RST), .Y(n1954) );
  OAI21X1 U102 ( .A(n287), .B(n1728), .C(n1953), .Y(n1888) );
  NAND2X1 U103 ( .A(PLAINKEY[31]), .B(n288), .Y(n1953) );
  OAI21X1 U105 ( .A(n287), .B(n1727), .C(n1952), .Y(n1887) );
  NAND2X1 U106 ( .A(PLAINKEY[32]), .B(n286), .Y(n1952) );
  OAI21X1 U108 ( .A(n286), .B(n1726), .C(n1951), .Y(n1886) );
  NAND2X1 U109 ( .A(PLAINKEY[33]), .B(n287), .Y(n1951) );
  OAI21X1 U111 ( .A(n287), .B(n1725), .C(n1950), .Y(n1885) );
  NAND2X1 U112 ( .A(PLAINKEY[34]), .B(n285), .Y(n1950) );
  OAI21X1 U114 ( .A(n286), .B(n1724), .C(n1949), .Y(n1884) );
  NAND2X1 U115 ( .A(PLAINKEY[35]), .B(n284), .Y(n1949) );
  OAI21X1 U117 ( .A(n286), .B(n1723), .C(n1948), .Y(n1883) );
  NAND2X1 U118 ( .A(PLAINKEY[36]), .B(RST), .Y(n1948) );
  OAI21X1 U120 ( .A(n287), .B(n1722), .C(n1947), .Y(n1882) );
  NAND2X1 U121 ( .A(PLAINKEY[37]), .B(n286), .Y(n1947) );
  OAI21X1 U123 ( .A(n287), .B(n1721), .C(n1946), .Y(n1881) );
  NAND2X1 U124 ( .A(PLAINKEY[38]), .B(RST), .Y(n1946) );
  OAI21X1 U126 ( .A(n287), .B(n1720), .C(n1945), .Y(n1880) );
  NAND2X1 U127 ( .A(PLAINKEY[39]), .B(n288), .Y(n1945) );
  OAI21X1 U129 ( .A(n287), .B(n1719), .C(n1944), .Y(n1879) );
  NAND2X1 U130 ( .A(PLAINKEY[40]), .B(RST), .Y(n1944) );
  OAI21X1 U132 ( .A(n287), .B(n1718), .C(n1943), .Y(n1878) );
  NAND2X1 U133 ( .A(PLAINKEY[41]), .B(n287), .Y(n1943) );
  OAI21X1 U135 ( .A(n286), .B(n1717), .C(n1942), .Y(n1877) );
  NAND2X1 U136 ( .A(PLAINKEY[42]), .B(n285), .Y(n1942) );
  OAI21X1 U138 ( .A(n287), .B(n1716), .C(n1941), .Y(n1876) );
  NAND2X1 U139 ( .A(PLAINKEY[43]), .B(n286), .Y(n1941) );
  OAI21X1 U141 ( .A(n287), .B(n1715), .C(n1940), .Y(n1875) );
  NAND2X1 U142 ( .A(PLAINKEY[44]), .B(n287), .Y(n1940) );
  OAI21X1 U144 ( .A(n287), .B(n1714), .C(n1939), .Y(n1874) );
  NAND2X1 U145 ( .A(PLAINKEY[45]), .B(n284), .Y(n1939) );
  OAI21X1 U147 ( .A(n287), .B(n1713), .C(n1938), .Y(n1873) );
  NAND2X1 U148 ( .A(PLAINKEY[46]), .B(RST), .Y(n1938) );
  OAI21X1 U150 ( .A(n284), .B(n1712), .C(n1937), .Y(n1872) );
  NAND2X1 U151 ( .A(PLAINKEY[47]), .B(n287), .Y(n1937) );
  OAI21X1 U153 ( .A(n286), .B(n1711), .C(n1936), .Y(n1871) );
  NAND2X1 U154 ( .A(PLAINKEY[48]), .B(n285), .Y(n1936) );
  OAI21X1 U156 ( .A(n286), .B(n1710), .C(n1935), .Y(n1870) );
  NAND2X1 U157 ( .A(PLAINKEY[49]), .B(n287), .Y(n1935) );
  OAI21X1 U159 ( .A(n286), .B(n1709), .C(n1934), .Y(n1869) );
  NAND2X1 U160 ( .A(PLAINKEY[50]), .B(n284), .Y(n1934) );
  OAI21X1 U162 ( .A(n285), .B(n1708), .C(n1933), .Y(n1868) );
  NAND2X1 U163 ( .A(PLAINKEY[51]), .B(n286), .Y(n1933) );
  OAI21X1 U165 ( .A(n286), .B(n1707), .C(n1932), .Y(n1867) );
  NAND2X1 U166 ( .A(PLAINKEY[52]), .B(RST), .Y(n1932) );
  OAI21X1 U168 ( .A(n285), .B(n1706), .C(n1931), .Y(n1866) );
  NAND2X1 U169 ( .A(PLAINKEY[53]), .B(n285), .Y(n1931) );
  OAI21X1 U171 ( .A(n285), .B(n1705), .C(n1930), .Y(n1865) );
  NAND2X1 U172 ( .A(PLAINKEY[54]), .B(n286), .Y(n1930) );
  OAI21X1 U174 ( .A(n284), .B(n1704), .C(n1929), .Y(n1864) );
  NAND2X1 U175 ( .A(PLAINKEY[55]), .B(n287), .Y(n1929) );
  OAI21X1 U177 ( .A(n285), .B(n1703), .C(n1928), .Y(n1863) );
  NAND2X1 U178 ( .A(PLAINKEY[56]), .B(RST), .Y(n1928) );
  OAI21X1 U180 ( .A(n284), .B(n1702), .C(n1927), .Y(n1862) );
  NAND2X1 U181 ( .A(PLAINKEY[57]), .B(n288), .Y(n1927) );
  OAI21X1 U183 ( .A(n284), .B(n1701), .C(n1926), .Y(n1861) );
  NAND2X1 U184 ( .A(PLAINKEY[58]), .B(n285), .Y(n1926) );
  OAI21X1 U186 ( .A(n284), .B(n1700), .C(n1925), .Y(n1860) );
  NAND2X1 U187 ( .A(PLAINKEY[59]), .B(n287), .Y(n1925) );
  OAI21X1 U188 ( .A(RST), .B(n1699), .C(n1924), .Y(n1859) );
  NAND2X1 U189 ( .A(PLAINKEY[60]), .B(n285), .Y(n1924) );
  OAI21X1 U191 ( .A(RST), .B(n1698), .C(n1923), .Y(n1858) );
  NAND2X1 U192 ( .A(PLAINKEY[61]), .B(n288), .Y(n1923) );
  OAI21X1 U194 ( .A(n288), .B(n1685), .C(n1922), .Y(n1857) );
  NAND2X1 U195 ( .A(PLAINKEY[62]), .B(n284), .Y(n1922) );
  OAI21X1 U196 ( .A(n286), .B(n1697), .C(n1921), .Y(n1856) );
  NAND2X1 U197 ( .A(PLAINKEY[63]), .B(n284), .Y(n1921) );
  NAND2X1 U1305 ( .A(n1648), .B(n1760), .Y(n1920) );
  keyreg_0_DW01_add_1 r577 ( .A(parityAccumulator), .B({RCV_DATA[7:3], n281, 
        RCV_DATA[1], n220}), .CI(1'b0), .SUM({N1799, N1798, N1797, N1796, 
        N1795, N1794, N1793, N1792}) );
  INVX2 U3 ( .A(n747), .Y(n678) );
  INVX1 U4 ( .A(n135), .Y(n1163) );
  INVX1 U5 ( .A(n137), .Y(n849) );
  INVX2 U7 ( .A(n849), .Y(n785) );
  INVX2 U8 ( .A(n164), .Y(n303) );
  INVX4 U23 ( .A(n67), .Y(n177) );
  INVX2 U26 ( .A(n1372), .Y(n1520) );
  BUFX2 U29 ( .A(n550), .Y(n53) );
  INVX1 U32 ( .A(n691), .Y(n103) );
  INVX1 U35 ( .A(n968), .Y(n152) );
  INVX1 U38 ( .A(n1039), .Y(n107) );
  BUFX2 U41 ( .A(n190), .Y(n277) );
  INVX4 U44 ( .A(n163), .Y(n164) );
  INVX2 U47 ( .A(n1021), .Y(n1051) );
  INVX2 U50 ( .A(n1480), .Y(n1437) );
  INVX2 U53 ( .A(n744), .Y(n774) );
  INVX1 U56 ( .A(n205), .Y(n206) );
  INVX2 U59 ( .A(n1542), .Y(n205) );
  AND2X1 U62 ( .A(n188), .B(n221), .Y(n1) );
  INVX2 U65 ( .A(n847), .Y(n824) );
  AND2X2 U68 ( .A(n312), .B(n727), .Y(n2) );
  INVX2 U71 ( .A(n637), .Y(n614) );
  INVX2 U74 ( .A(n604), .Y(n585) );
  INVX2 U77 ( .A(n1481), .Y(n1444) );
  INVX2 U80 ( .A(n201), .Y(n202) );
  INVX2 U83 ( .A(n1506), .Y(n201) );
  INVX2 U86 ( .A(n1122), .Y(n1105) );
  INVX1 U89 ( .A(n283), .Y(n282) );
  INVX1 U92 ( .A(n1372), .Y(n69) );
  INVX4 U95 ( .A(n117), .Y(n275) );
  INVX2 U98 ( .A(n916), .Y(n892) );
  AND2X1 U101 ( .A(n1462), .B(n1464), .Y(n4) );
  INVX1 U104 ( .A(n1515), .Y(n5) );
  INVX1 U107 ( .A(n946), .Y(n6) );
  BUFX2 U110 ( .A(n1504), .Y(n7) );
  BUFX2 U113 ( .A(n413), .Y(n8) );
  INVX1 U116 ( .A(n1155), .Y(n9) );
  INVX2 U119 ( .A(n1121), .Y(n1155) );
  INVX1 U122 ( .A(n1190), .Y(n10) );
  INVX1 U125 ( .A(n910), .Y(n11) );
  NAND2X1 U128 ( .A(n1660), .B(n319), .Y(n14) );
  INVX4 U131 ( .A(n197), .Y(n1660) );
  BUFX4 U134 ( .A(n1482), .Y(n251) );
  BUFX4 U137 ( .A(n1466), .Y(n16) );
  OR2X2 U140 ( .A(n1529), .B(n111), .Y(n17) );
  INVX1 U143 ( .A(n17), .Y(n115) );
  INVX1 U146 ( .A(n632), .Y(n19) );
  INVX2 U149 ( .A(n1364), .Y(n20) );
  INVX1 U152 ( .A(n1460), .Y(n21) );
  INVX2 U155 ( .A(n1651), .Y(n23) );
  INVX2 U158 ( .A(n648), .Y(n25) );
  INVX2 U161 ( .A(n1444), .Y(n27) );
  INVX4 U164 ( .A(n739), .Y(n29) );
  INVX2 U167 ( .A(n708), .Y(n739) );
  INVX4 U170 ( .A(n841), .Y(n31) );
  INVX2 U173 ( .A(n814), .Y(n841) );
  INVX4 U176 ( .A(n1016), .Y(n33) );
  INVX2 U179 ( .A(n985), .Y(n1016) );
  BUFX2 U182 ( .A(n1602), .Y(n35) );
  INVX4 U185 ( .A(n809), .Y(n37) );
  INVX2 U190 ( .A(n779), .Y(n809) );
  INVX4 U193 ( .A(n1084), .Y(n39) );
  INVX2 U198 ( .A(n1056), .Y(n1084) );
  INVX1 U199 ( .A(n980), .Y(n41) );
  INVX2 U200 ( .A(n1407), .Y(n43) );
  INVX2 U201 ( .A(n926), .Y(n45) );
  INVX1 U202 ( .A(n952), .Y(n926) );
  AND2X2 U203 ( .A(n49), .B(n327), .Y(n47) );
  INVX1 U204 ( .A(n47), .Y(n1142) );
  NOR2X1 U205 ( .A(address[1]), .B(address[0]), .Y(n49) );
  INVX1 U206 ( .A(n1419), .Y(n51) );
  INVX1 U207 ( .A(n703), .Y(n55) );
  BUFX2 U208 ( .A(n567), .Y(n57) );
  INVX1 U209 ( .A(n1384), .Y(n59) );
  INVX2 U210 ( .A(n1195), .Y(n1384) );
  INVX2 U211 ( .A(n1557), .Y(n61) );
  INVX4 U212 ( .A(n1578), .Y(n1557) );
  INVX4 U213 ( .A(n1571), .Y(n63) );
  INVX4 U214 ( .A(n1503), .Y(n1571) );
  INVX2 U215 ( .A(n1437), .Y(n65) );
  INVX1 U216 ( .A(address[0]), .Y(n324) );
  OR2X2 U217 ( .A(n335), .B(n222), .Y(n67) );
  INVX2 U218 ( .A(n335), .Y(n586) );
  INVX2 U219 ( .A(n1424), .Y(n1460) );
  INVX1 U220 ( .A(n69), .Y(n71) );
  INVX2 U221 ( .A(n603), .Y(n632) );
  AND2X2 U222 ( .A(n604), .B(n603), .Y(n123) );
  INVX2 U223 ( .A(n1176), .Y(n73) );
  INVX1 U224 ( .A(n73), .Y(n75) );
  INVX2 U225 ( .A(n189), .Y(n77) );
  INVX4 U226 ( .A(n77), .Y(n79) );
  BUFX2 U227 ( .A(n131), .Y(n81) );
  INVX4 U228 ( .A(n562), .Y(n83) );
  INVX4 U229 ( .A(n545), .Y(n562) );
  MUX2X1 U230 ( .B(n271), .A(n1489), .S(n1524), .Y(n1490) );
  INVX1 U231 ( .A(n1524), .Y(n1596) );
  BUFX2 U232 ( .A(n125), .Y(n85) );
  INVX4 U233 ( .A(n497), .Y(n87) );
  INVX4 U234 ( .A(n478), .Y(n497) );
  INVX1 U235 ( .A(n1175), .Y(n89) );
  NAND2X1 U236 ( .A(n1463), .B(n4), .Y(n1842) );
  AND2X2 U237 ( .A(n916), .B(n915), .Y(n149) );
  MUX2X1 U238 ( .B(n283), .A(n1491), .S(n1529), .Y(n1492) );
  INVX1 U239 ( .A(n1529), .Y(n1598) );
  BUFX2 U240 ( .A(n174), .Y(n91) );
  INVX1 U241 ( .A(n863), .Y(n93) );
  INVX1 U242 ( .A(n125), .Y(n457) );
  INVX2 U243 ( .A(n1160), .Y(n1190) );
  AND2X2 U244 ( .A(n1090), .B(n1089), .Y(n95) );
  INVX1 U245 ( .A(n95), .Y(n1092) );
  INVX2 U246 ( .A(n1092), .Y(n1102) );
  BUFX2 U247 ( .A(n73), .Y(n159) );
  INVX2 U248 ( .A(n881), .Y(n910) );
  AND2X1 U249 ( .A(n745), .B(n744), .Y(n97) );
  INVX1 U250 ( .A(n97), .Y(n747) );
  AND2X1 U251 ( .A(n1022), .B(n1021), .Y(n99) );
  INVX1 U252 ( .A(n99), .Y(n1024) );
  INVX2 U253 ( .A(n1024), .Y(n1036) );
  INVX2 U254 ( .A(n585), .Y(n101) );
  MUX2X1 U255 ( .B(n262), .A(n665), .S(n103), .Y(n667) );
  BUFX2 U256 ( .A(address[2]), .Y(n105) );
  AND2X2 U257 ( .A(n1196), .B(n1195), .Y(n154) );
  INVX1 U258 ( .A(n37), .Y(n756) );
  MUX2X1 U259 ( .B(n261), .A(n1013), .S(n107), .Y(n1015) );
  INVX1 U260 ( .A(n29), .Y(n684) );
  NAND2X1 U261 ( .A(n299), .B(n109), .Y(n1664) );
  AND2X1 U262 ( .A(n226), .B(n164), .Y(n109) );
  OR2X2 U263 ( .A(n1529), .B(n271), .Y(n113) );
  INVX1 U264 ( .A(n168), .Y(n111) );
  AND2X2 U265 ( .A(RCV_DATA[6]), .B(n228), .Y(n117) );
  INVX2 U266 ( .A(n672), .Y(n703) );
  AND2X2 U267 ( .A(n479), .B(n478), .Y(n125) );
  INVX2 U268 ( .A(n888), .Y(n1141) );
  INVX2 U269 ( .A(n951), .Y(n980) );
  AND2X2 U270 ( .A(n1465), .B(n1453), .Y(n119) );
  INVX1 U271 ( .A(n119), .Y(n1493) );
  BUFX4 U272 ( .A(n1577), .Y(n266) );
  BUFX2 U273 ( .A(n450), .Y(n121) );
  INVX2 U274 ( .A(n1389), .Y(n1419) );
  INVX2 U275 ( .A(n782), .Y(n753) );
  INVX2 U276 ( .A(n711), .Y(n681) );
  INVX1 U277 ( .A(n123), .Y(n606) );
  AND2X2 U278 ( .A(n673), .B(n672), .Y(n141) );
  INVX2 U279 ( .A(n673), .Y(n656) );
  INVX1 U280 ( .A(n39), .Y(n1032) );
  INVX1 U281 ( .A(n1059), .Y(n993) );
  BUFX2 U282 ( .A(n14), .Y(n230) );
  INVX1 U283 ( .A(n988), .Y(n921) );
  AND2X1 U284 ( .A(n1122), .B(n1121), .Y(n127) );
  INVX2 U285 ( .A(n127), .Y(n1124) );
  INVX2 U286 ( .A(n1124), .Y(n1137) );
  BUFX4 U287 ( .A(n190), .Y(n280) );
  OR2X2 U288 ( .A(n166), .B(n1644), .Y(n1613) );
  INVX2 U289 ( .A(n166), .Y(n1609) );
  INVX2 U290 ( .A(state[0]), .Y(n163) );
  OR2X2 U291 ( .A(n230), .B(n283), .Y(n1466) );
  AND2X2 U292 ( .A(n1425), .B(n1424), .Y(n129) );
  INVX2 U293 ( .A(n129), .Y(n1427) );
  INVX2 U294 ( .A(n1427), .Y(n1441) );
  AND2X2 U295 ( .A(n546), .B(n545), .Y(n131) );
  INVX1 U296 ( .A(n131), .Y(n524) );
  INVX4 U297 ( .A(n155), .Y(n169) );
  AND2X2 U298 ( .A(n513), .B(n512), .Y(n133) );
  INVX1 U299 ( .A(n133), .Y(n491) );
  AND2X2 U300 ( .A(n1161), .B(n1160), .Y(n135) );
  AND2X1 U301 ( .A(n847), .B(n846), .Y(n137) );
  AND2X2 U302 ( .A(n882), .B(n881), .Y(n139) );
  INVX2 U303 ( .A(n139), .Y(n884) );
  INVX2 U304 ( .A(n884), .Y(n896) );
  BUFX4 U305 ( .A(n184), .Y(n242) );
  BUFX4 U306 ( .A(n1428), .Y(n231) );
  INVX2 U307 ( .A(n141), .Y(n675) );
  INVX2 U308 ( .A(n675), .Y(n688) );
  BUFX4 U309 ( .A(n184), .Y(n243) );
  INVX8 U310 ( .A(n243), .Y(n240) );
  INVX1 U311 ( .A(n1551), .Y(n143) );
  INVX2 U312 ( .A(n1519), .Y(n1551) );
  AND2X2 U313 ( .A(n1390), .B(n1389), .Y(n145) );
  INVX2 U314 ( .A(n145), .Y(n1392) );
  INVX2 U315 ( .A(n1392), .Y(n1404) );
  AND2X2 U316 ( .A(n1481), .B(n1480), .Y(n147) );
  INVX1 U317 ( .A(n147), .Y(n1454) );
  BUFX4 U318 ( .A(n1482), .Y(n249) );
  INVX4 U319 ( .A(n181), .Y(n264) );
  INVX2 U320 ( .A(n264), .Y(n263) );
  BUFX4 U321 ( .A(n184), .Y(n245) );
  INVX2 U322 ( .A(n149), .Y(n918) );
  INVX2 U323 ( .A(n918), .Y(n931) );
  AND2X1 U324 ( .A(n638), .B(n637), .Y(n150) );
  INVX1 U325 ( .A(n150), .Y(n640) );
  INVX2 U326 ( .A(n640), .Y(n653) );
  INVX4 U327 ( .A(n117), .Y(n276) );
  INVX4 U328 ( .A(n256), .Y(n253) );
  INVX1 U329 ( .A(n328), .Y(n151) );
  INVX8 U330 ( .A(n249), .Y(n248) );
  MUX2X1 U331 ( .B(n261), .A(n943), .S(n152), .Y(n945) );
  INVX1 U332 ( .A(n568), .Y(n550) );
  AND2X1 U333 ( .A(n952), .B(n951), .Y(n153) );
  INVX1 U334 ( .A(n153), .Y(n954) );
  INVX2 U335 ( .A(n954), .Y(n965) );
  INVX1 U336 ( .A(n673), .Y(n648) );
  INVX1 U337 ( .A(n154), .Y(n1268) );
  INVX2 U338 ( .A(n1268), .Y(n1368) );
  INVX4 U339 ( .A(n161), .Y(n182) );
  INVX1 U340 ( .A(n1390), .Y(n1364) );
  INVX8 U341 ( .A(n244), .Y(n239) );
  INVX8 U342 ( .A(n249), .Y(n247) );
  INVX4 U343 ( .A(n256), .Y(n254) );
  BUFX4 U344 ( .A(n1466), .Y(n238) );
  INVX1 U345 ( .A(n224), .Y(n306) );
  OR2X2 U346 ( .A(n1582), .B(n222), .Y(n155) );
  INVX2 U347 ( .A(n1582), .Y(n1561) );
  MUX2X1 U348 ( .B(n247), .A(n1052), .S(n1021), .Y(n1054) );
  NAND2X1 U349 ( .A(n1660), .B(n319), .Y(n156) );
  INVX4 U350 ( .A(n191), .Y(n204) );
  AND2X2 U351 ( .A(address[1]), .B(address[2]), .Y(n194) );
  AND2X2 U352 ( .A(n1520), .B(n223), .Y(n157) );
  BUFX2 U353 ( .A(n864), .Y(n158) );
  INVX2 U354 ( .A(n610), .Y(n864) );
  INVX1 U355 ( .A(address[6]), .Y(n1696) );
  INVX1 U356 ( .A(n1453), .Y(n1534) );
  INVX1 U357 ( .A(n782), .Y(n716) );
  INVX1 U358 ( .A(n31), .Y(n791) );
  INVX1 U359 ( .A(n817), .Y(n750) );
  INVX8 U360 ( .A(n250), .Y(n246) );
  INVX1 U361 ( .A(n711), .Y(n643) );
  INVX4 U362 ( .A(n258), .Y(n256) );
  INVX2 U363 ( .A(n256), .Y(n255) );
  INVX1 U364 ( .A(n55), .Y(n649) );
  BUFX2 U365 ( .A(address[0]), .Y(n160) );
  OR2X2 U366 ( .A(n888), .B(n222), .Y(n161) );
  BUFX2 U367 ( .A(n1520), .Y(n162) );
  INVX2 U368 ( .A(n1612), .Y(n165) );
  INVX4 U369 ( .A(n165), .Y(n166) );
  INVX4 U370 ( .A(n265), .Y(n262) );
  INVX4 U371 ( .A(n265), .Y(n261) );
  BUFX4 U372 ( .A(n1466), .Y(n237) );
  INVX1 U373 ( .A(n21), .Y(n1400) );
  INVX1 U374 ( .A(n41), .Y(n927) );
  INVX4 U375 ( .A(n264), .Y(n260) );
  INVX1 U376 ( .A(n1664), .Y(n1651) );
  INVX1 U377 ( .A(n245), .Y(n167) );
  INVX2 U378 ( .A(n264), .Y(n259) );
  INVX1 U379 ( .A(n172), .Y(n235) );
  BUFX4 U380 ( .A(n184), .Y(n244) );
  INVX4 U381 ( .A(n257), .Y(n252) );
  INVX4 U382 ( .A(n283), .Y(n281) );
  INVX2 U383 ( .A(n1505), .Y(n258) );
  INVX2 U384 ( .A(n1584), .Y(n274) );
  INVX2 U385 ( .A(address[3]), .Y(n221) );
  INVX2 U386 ( .A(n290), .Y(n286) );
  INVX2 U387 ( .A(n290), .Y(n285) );
  INVX2 U388 ( .A(n289), .Y(n284) );
  INVX2 U389 ( .A(n291), .Y(n287) );
  INVX2 U390 ( .A(n291), .Y(n288) );
  AND2X2 U391 ( .A(n1468), .B(n228), .Y(n168) );
  BUFX2 U392 ( .A(n293), .Y(n291) );
  BUFX2 U393 ( .A(n293), .Y(n290) );
  BUFX2 U394 ( .A(n293), .Y(n289) );
  BUFX2 U395 ( .A(n289), .Y(n292) );
  BUFX2 U396 ( .A(n1577), .Y(n267) );
  BUFX2 U397 ( .A(n1577), .Y(n269) );
  INVX4 U398 ( .A(n156), .Y(n229) );
  INVX4 U399 ( .A(n232), .Y(n227) );
  INVX2 U400 ( .A(n172), .Y(n233) );
  INVX2 U401 ( .A(n172), .Y(n234) );
  AND2X2 U402 ( .A(n176), .B(n1561), .Y(n170) );
  BUFX2 U403 ( .A(n1577), .Y(n270) );
  INVX2 U404 ( .A(n242), .Y(n241) );
  INVX2 U405 ( .A(RST), .Y(n293) );
  AND2X2 U406 ( .A(n325), .B(n176), .Y(n171) );
  AND2X2 U407 ( .A(n403), .B(n185), .Y(n172) );
  AND2X2 U408 ( .A(n1520), .B(n223), .Y(n173) );
  AND2X2 U409 ( .A(n73), .B(n223), .Y(n174) );
  AND2X2 U410 ( .A(n201), .B(n223), .Y(n175) );
  AND2X2 U411 ( .A(n205), .B(n223), .Y(n176) );
  INVX2 U412 ( .A(n181), .Y(n265) );
  AND2X2 U413 ( .A(n223), .B(n47), .Y(n178) );
  AND2X2 U414 ( .A(n191), .B(n223), .Y(n179) );
  INVX2 U415 ( .A(n207), .Y(n208) );
  INVX2 U416 ( .A(n207), .Y(n209) );
  AND2X2 U417 ( .A(n325), .B(n91), .Y(n180) );
  INVX2 U418 ( .A(n571), .Y(n207) );
  BUFX2 U419 ( .A(n190), .Y(n278) );
  BUFX2 U420 ( .A(n190), .Y(n279) );
  AND2X2 U421 ( .A(n343), .B(n185), .Y(n181) );
  INVX2 U422 ( .A(n274), .Y(n272) );
  INVX2 U423 ( .A(n274), .Y(n271) );
  INVX2 U424 ( .A(n1), .Y(n218) );
  AND2X2 U425 ( .A(n864), .B(n221), .Y(n183) );
  AND2X2 U426 ( .A(n339), .B(n185), .Y(n184) );
  AND2X2 U427 ( .A(n319), .B(n309), .Y(n185) );
  INVX2 U428 ( .A(n258), .Y(n257) );
  AND2X2 U429 ( .A(n194), .B(n324), .Y(n186) );
  AND2X2 U430 ( .A(n226), .B(n225), .Y(n187) );
  INVX2 U431 ( .A(n221), .Y(n223) );
  INVX2 U432 ( .A(n274), .Y(n273) );
  INVX2 U433 ( .A(n221), .Y(n222) );
  INVX2 U434 ( .A(RCV_DATA[2]), .Y(n283) );
  BUFX4 U435 ( .A(state[2]), .Y(n225) );
  BUFX4 U436 ( .A(state[1]), .Y(n226) );
  INVX2 U437 ( .A(n210), .Y(n211) );
  INVX2 U438 ( .A(n712), .Y(n210) );
  INVX2 U439 ( .A(n214), .Y(n215) );
  INVX2 U440 ( .A(n989), .Y(n214) );
  INVX4 U441 ( .A(n212), .Y(n213) );
  INVX2 U442 ( .A(n850), .Y(n212) );
  INVX4 U443 ( .A(n216), .Y(n217) );
  INVX2 U444 ( .A(n1125), .Y(n216) );
  INVX4 U445 ( .A(n219), .Y(n220) );
  INVX2 U446 ( .A(RCV_DATA[0]), .Y(n219) );
  AND2X2 U447 ( .A(address[4]), .B(address[5]), .Y(n188) );
  NOR2X1 U448 ( .A(address[6]), .B(address[7]), .Y(n189) );
  AND2X2 U449 ( .A(RCV_DATA[6]), .B(n228), .Y(n190) );
  AND2X2 U450 ( .A(n194), .B(n160), .Y(n191) );
  INVX4 U451 ( .A(n2), .Y(n203) );
  NOR2X1 U452 ( .A(n224), .B(n164), .Y(n192) );
  NOR2X1 U453 ( .A(n226), .B(n164), .Y(n193) );
  INVX2 U454 ( .A(n1469), .Y(n195) );
  INVX1 U455 ( .A(n195), .Y(n196) );
  BUFX4 U456 ( .A(n1672), .Y(n197) );
  BUFX2 U457 ( .A(n1672), .Y(n198) );
  INVX1 U458 ( .A(n186), .Y(n199) );
  INVX1 U459 ( .A(n186), .Y(n200) );
  BUFX4 U460 ( .A(state[3]), .Y(n224) );
  INVX1 U461 ( .A(n166), .Y(n1611) );
  BUFX2 U462 ( .A(n14), .Y(n232) );
  INVX8 U463 ( .A(n231), .Y(n228) );
  BUFX4 U464 ( .A(n1466), .Y(n236) );
  BUFX4 U465 ( .A(n1482), .Y(n250) );
  BUFX4 U466 ( .A(n1577), .Y(n268) );
  NOR2X1 U467 ( .A(n224), .B(n225), .Y(n294) );
  NAND3X1 U468 ( .A(n226), .B(n303), .C(n294), .Y(n1672) );
  INVX2 U469 ( .A(n226), .Y(n297) );
  NOR2X1 U470 ( .A(n224), .B(n297), .Y(n295) );
  NAND3X1 U471 ( .A(n225), .B(n164), .C(n295), .Y(n1642) );
  NAND2X1 U472 ( .A(n197), .B(n1642), .Y(CLR_RBUFF) );
  NOR2X1 U473 ( .A(n224), .B(n164), .Y(n296) );
  NAND3X1 U474 ( .A(n225), .B(n297), .C(n296), .Y(n1620) );
  INVX2 U475 ( .A(n1620), .Y(PROG_ERROR) );
  NOR2X1 U476 ( .A(n226), .B(n225), .Y(n298) );
  NAND2X1 U477 ( .A(n298), .B(n303), .Y(n1662) );
  NOR2X1 U478 ( .A(n224), .B(n225), .Y(n299) );
  OAI21X1 U479 ( .A(n224), .B(n1662), .C(n1664), .Y(n301) );
  NAND2X1 U480 ( .A(n187), .B(n192), .Y(n1661) );
  NAND2X1 U481 ( .A(n1661), .B(n1620), .Y(n300) );
  NOR3X1 U482 ( .A(CLR_RBUFF), .B(n301), .C(n300), .Y(n1602) );
  NOR2X1 U483 ( .A(n225), .B(n306), .Y(n302) );
  NAND2X1 U484 ( .A(n302), .B(n193), .Y(n1663) );
  NOR2X1 U485 ( .A(n224), .B(n303), .Y(n304) );
  NAND3X1 U486 ( .A(n225), .B(n297), .C(n304), .Y(n1669) );
  INVX2 U487 ( .A(n1669), .Y(n1647) );
  NOR2X1 U488 ( .A(n226), .B(n225), .Y(n305) );
  NAND3X1 U489 ( .A(n164), .B(n306), .C(n305), .Y(n1657) );
  INVX2 U490 ( .A(n1657), .Y(n1615) );
  AOI21X1 U491 ( .A(n1647), .B(parityError), .C(n1615), .Y(n307) );
  NAND3X1 U492 ( .A(n35), .B(n1663), .C(n307), .Y(KEY_ERROR) );
  INVX2 U493 ( .A(currentPlainKey[63]), .Y(n1697) );
  INVX2 U494 ( .A(currentPlainKey[62]), .Y(n1685) );
  INVX2 U495 ( .A(currentPlainKey[3]), .Y(n1756) );
  INVX2 U496 ( .A(currentPlainKey[2]), .Y(n1757) );
  INVX2 U497 ( .A(currentPlainKey[1]), .Y(n1758) );
  INVX2 U498 ( .A(currentPlainKey[0]), .Y(n1759) );
  INVX2 U499 ( .A(parityAccumulator[4]), .Y(n1692) );
  INVX2 U500 ( .A(parityAccumulator[5]), .Y(n1693) );
  AOI21X1 U501 ( .A(n187), .B(n192), .C(n287), .Y(n308) );
  AND2X2 U502 ( .A(n308), .B(n1664), .Y(n319) );
  AND2X2 U503 ( .A(n1657), .B(n1620), .Y(n309) );
  NAND3X1 U504 ( .A(n1663), .B(n1642), .C(n185), .Y(n310) );
  INVX2 U505 ( .A(n310), .Y(n1683) );
  NAND2X1 U506 ( .A(n1683), .B(n1669), .Y(n1577) );
  NAND2X1 U507 ( .A(n270), .B(currentPlainKey[0]), .Y(n333) );
  NAND3X1 U508 ( .A(address[6]), .B(address[7]), .C(n188), .Y(n329) );
  INVX2 U509 ( .A(n329), .Y(n325) );
  INVX2 U510 ( .A(address[1]), .Y(n328) );
  NAND3X1 U511 ( .A(address[2]), .B(n324), .C(n328), .Y(n1372) );
  NAND2X1 U512 ( .A(n325), .B(n173), .Y(n311) );
  INVX2 U513 ( .A(n311), .Y(n380) );
  INVX2 U514 ( .A(RCV_DATA[4]), .Y(n342) );
  NAND2X1 U515 ( .A(n380), .B(n342), .Y(n323) );
  NAND2X1 U516 ( .A(n186), .B(n223), .Y(n1581) );
  INVX2 U517 ( .A(n1581), .Y(n1130) );
  NAND2X1 U518 ( .A(n325), .B(n1130), .Y(n412) );
  INVX2 U519 ( .A(n412), .Y(n384) );
  INVX2 U520 ( .A(address[2]), .Y(n327) );
  NAND3X1 U521 ( .A(address[1]), .B(address[0]), .C(n327), .Y(n1506) );
  NAND2X1 U522 ( .A(n325), .B(n175), .Y(n345) );
  NAND2X1 U523 ( .A(n345), .B(n311), .Y(n361) );
  AOI21X1 U524 ( .A(n384), .B(n281), .C(n361), .Y(n318) );
  NOR2X1 U525 ( .A(address[4]), .B(n222), .Y(n312) );
  INVX2 U526 ( .A(address[5]), .Y(n727) );
  INVX2 U527 ( .A(n203), .Y(n368) );
  NAND2X1 U528 ( .A(n368), .B(n47), .Y(n313) );
  NAND2X1 U529 ( .A(n220), .B(n47), .Y(n1144) );
  INVX2 U530 ( .A(n1144), .Y(n1445) );
  AOI22X1 U531 ( .A(n313), .B(currentPlainKey[0]), .C(n368), .D(n1445), .Y(
        n315) );
  NAND2X1 U532 ( .A(n325), .B(n179), .Y(n413) );
  NAND2X1 U533 ( .A(n412), .B(n413), .Y(n391) );
  INVX2 U534 ( .A(n413), .Y(n430) );
  NAND2X1 U535 ( .A(n430), .B(RCV_DATA[1]), .Y(n314) );
  OAI21X1 U536 ( .A(n315), .B(n391), .C(n314), .Y(n316) );
  NAND3X1 U537 ( .A(address[2]), .B(address[0]), .C(n328), .Y(n1542) );
  MUX2X1 U538 ( .B(n316), .A(RCV_DATA[3]), .S(n171), .Y(n317) );
  NAND2X1 U539 ( .A(n318), .B(n317), .Y(n322) );
  NAND2X1 U540 ( .A(n1660), .B(n319), .Y(n1428) );
  NAND2X1 U541 ( .A(n229), .B(n345), .Y(n320) );
  NAND3X1 U542 ( .A(n185), .B(RCV_DATA[5]), .C(n1660), .Y(n1505) );
  NAND2X1 U543 ( .A(n320), .B(n257), .Y(n321) );
  NAND3X1 U544 ( .A(n323), .B(n322), .C(n321), .Y(n326) );
  NAND3X1 U545 ( .A(address[1]), .B(n324), .C(n327), .Y(n1176) );
  MUX2X1 U546 ( .B(n326), .A(n276), .S(n180), .Y(n331) );
  NAND2X1 U547 ( .A(RCV_DATA[7]), .B(n228), .Y(n1482) );
  NAND3X1 U548 ( .A(n328), .B(address[0]), .C(n327), .Y(n1469) );
  NAND2X1 U549 ( .A(n195), .B(n223), .Y(n484) );
  NOR2X1 U550 ( .A(n484), .B(n329), .Y(n330) );
  MUX2X1 U551 ( .B(n331), .A(n248), .S(n330), .Y(n332) );
  NAND2X1 U552 ( .A(n333), .B(n332), .Y(n1786) );
  NAND2X1 U553 ( .A(n270), .B(currentPlainKey[1]), .Y(n350) );
  INVX2 U554 ( .A(n391), .Y(n411) );
  NAND2X1 U555 ( .A(n368), .B(n195), .Y(n334) );
  NAND2X1 U556 ( .A(n220), .B(n195), .Y(n469) );
  INVX2 U557 ( .A(n469), .Y(n1470) );
  AOI22X1 U558 ( .A(n334), .B(currentPlainKey[1]), .C(n368), .D(n1470), .Y(
        n336) );
  INVX2 U559 ( .A(RCV_DATA[1]), .Y(n1584) );
  INVX2 U560 ( .A(address[4]), .Y(n1004) );
  NAND3X1 U561 ( .A(n79), .B(n1004), .C(n727), .Y(n335) );
  NAND2X1 U562 ( .A(n177), .B(n47), .Y(n446) );
  INVX2 U563 ( .A(n446), .Y(n417) );
  MUX2X1 U564 ( .B(n336), .A(n271), .S(n417), .Y(n338) );
  NOR2X1 U565 ( .A(n283), .B(n413), .Y(n337) );
  AOI21X1 U566 ( .A(n411), .B(n338), .C(n337), .Y(n341) );
  INVX2 U567 ( .A(RCV_DATA[3]), .Y(n1589) );
  NOR2X1 U568 ( .A(n1589), .B(n198), .Y(n339) );
  NAND2X1 U569 ( .A(n384), .B(n245), .Y(n340) );
  OAI21X1 U570 ( .A(n341), .B(n230), .C(n340), .Y(n344) );
  NOR2X1 U571 ( .A(n342), .B(n198), .Y(n343) );
  MUX2X1 U572 ( .B(n344), .A(n261), .S(n171), .Y(n347) );
  INVX2 U573 ( .A(n345), .Y(n351) );
  AOI22X1 U574 ( .A(n380), .B(n253), .C(n351), .D(n280), .Y(n346) );
  OAI21X1 U575 ( .A(n347), .B(n361), .C(n346), .Y(n348) );
  MUX2X1 U576 ( .B(n348), .A(n247), .S(n180), .Y(n349) );
  NAND2X1 U577 ( .A(n350), .B(n349), .Y(n1787) );
  AOI22X1 U578 ( .A(n267), .B(currentPlainKey[2]), .C(n351), .D(n246), .Y(n367) );
  NOR2X1 U579 ( .A(n265), .B(n412), .Y(n364) );
  NOR2X1 U580 ( .A(n241), .B(n8), .Y(n359) );
  NAND2X1 U581 ( .A(n417), .B(n281), .Y(n357) );
  OAI21X1 U582 ( .A(n75), .B(n203), .C(currentPlainKey[2]), .Y(n353) );
  NAND2X1 U583 ( .A(n73), .B(n220), .Y(n1179) );
  INVX2 U584 ( .A(n1179), .Y(n1486) );
  NAND2X1 U585 ( .A(n368), .B(n1486), .Y(n352) );
  NAND2X1 U586 ( .A(n177), .B(n195), .Y(n445) );
  NAND2X1 U587 ( .A(n446), .B(n445), .Y(n424) );
  AOI21X1 U588 ( .A(n353), .B(n352), .C(n424), .Y(n355) );
  INVX2 U589 ( .A(n445), .Y(n463) );
  AND2X2 U590 ( .A(n463), .B(RCV_DATA[1]), .Y(n354) );
  OAI21X1 U591 ( .A(n355), .B(n354), .C(n8), .Y(n356) );
  AOI21X1 U592 ( .A(n357), .B(n356), .C(n230), .Y(n358) );
  OAI21X1 U593 ( .A(n359), .B(n358), .C(n412), .Y(n360) );
  MUX2X1 U594 ( .B(n360), .A(n257), .S(n171), .Y(n363) );
  INVX2 U595 ( .A(n361), .Y(n362) );
  OAI21X1 U596 ( .A(n364), .B(n363), .C(n362), .Y(n366) );
  NAND2X1 U597 ( .A(n380), .B(n278), .Y(n365) );
  NAND3X1 U598 ( .A(n367), .B(n366), .C(n365), .Y(n1788) );
  NAND2X1 U599 ( .A(n269), .B(currentPlainKey[3]), .Y(n383) );
  NOR2X1 U600 ( .A(n257), .B(n412), .Y(n378) );
  OAI21X1 U601 ( .A(n202), .B(n203), .C(currentPlainKey[3]), .Y(n370) );
  NAND2X1 U602 ( .A(n220), .B(n201), .Y(n503) );
  INVX2 U603 ( .A(n503), .Y(n1357) );
  NAND2X1 U604 ( .A(n368), .B(n1357), .Y(n369) );
  NAND2X1 U605 ( .A(n370), .B(n369), .Y(n371) );
  NAND2X1 U606 ( .A(n177), .B(n159), .Y(n479) );
  INVX2 U607 ( .A(n479), .Y(n450) );
  MUX2X1 U608 ( .B(n371), .A(RCV_DATA[1]), .S(n450), .Y(n373) );
  NAND2X1 U609 ( .A(n463), .B(n282), .Y(n372) );
  OAI21X1 U610 ( .A(n373), .B(n424), .C(n372), .Y(n374) );
  AOI22X1 U611 ( .A(n417), .B(n242), .C(n374), .D(n227), .Y(n376) );
  NAND2X1 U612 ( .A(n430), .B(n263), .Y(n375) );
  OAI21X1 U613 ( .A(n376), .B(n391), .C(n375), .Y(n377) );
  NOR2X1 U614 ( .A(n378), .B(n377), .Y(n379) );
  MUX2X1 U615 ( .B(n379), .A(n276), .S(n171), .Y(n381) );
  MUX2X1 U616 ( .B(n381), .A(n247), .S(n380), .Y(n382) );
  NAND2X1 U617 ( .A(n383), .B(n382), .Y(n1789) );
  NAND2X1 U618 ( .A(n384), .B(n278), .Y(n400) );
  NAND2X1 U619 ( .A(n177), .B(n201), .Y(n478) );
  NAND2X1 U620 ( .A(n220), .B(n1520), .Y(n1521) );
  OAI21X1 U621 ( .A(n71), .B(n203), .C(currentPlainKey[4]), .Y(n385) );
  OAI21X1 U622 ( .A(n1521), .B(n203), .C(n385), .Y(n387) );
  NOR2X1 U623 ( .A(n271), .B(n87), .Y(n386) );
  AOI21X1 U624 ( .A(n125), .B(n387), .C(n386), .Y(n389) );
  NAND2X1 U625 ( .A(n450), .B(n282), .Y(n388) );
  OAI21X1 U626 ( .A(n463), .B(n389), .C(n388), .Y(n390) );
  NAND2X1 U627 ( .A(n229), .B(n390), .Y(n393) );
  NAND2X1 U628 ( .A(n463), .B(n245), .Y(n392) );
  AOI21X1 U629 ( .A(n393), .B(n392), .C(n391), .Y(n394) );
  MUX2X1 U630 ( .B(n394), .A(n262), .S(n417), .Y(n396) );
  NAND2X1 U631 ( .A(n430), .B(n254), .Y(n395) );
  NAND2X1 U632 ( .A(n396), .B(n395), .Y(n397) );
  MUX2X1 U633 ( .B(n397), .A(n247), .S(n171), .Y(n399) );
  NAND2X1 U634 ( .A(currentPlainKey[4]), .B(n266), .Y(n398) );
  NAND3X1 U635 ( .A(n400), .B(n399), .C(n398), .Y(n1790) );
  NAND2X1 U636 ( .A(n463), .B(n263), .Y(n409) );
  NAND2X1 U637 ( .A(n220), .B(n205), .Y(n1544) );
  OAI21X1 U638 ( .A(n206), .B(n203), .C(currentPlainKey[5]), .Y(n401) );
  OAI21X1 U639 ( .A(n1544), .B(n203), .C(n401), .Y(n402) );
  NAND3X1 U640 ( .A(n125), .B(n228), .C(n402), .Y(n404) );
  NOR2X1 U641 ( .A(n273), .B(n198), .Y(n403) );
  NAND2X1 U642 ( .A(n177), .B(n162), .Y(n513) );
  INVX2 U643 ( .A(n513), .Y(n483) );
  MUX2X1 U644 ( .B(n404), .A(n233), .S(n483), .Y(n406) );
  OAI22X1 U645 ( .A(n241), .B(n479), .C(n236), .D(n87), .Y(n405) );
  INVX2 U646 ( .A(n424), .Y(n444) );
  OAI21X1 U647 ( .A(n406), .B(n405), .C(n444), .Y(n408) );
  NAND2X1 U648 ( .A(n417), .B(n254), .Y(n407) );
  NAND3X1 U649 ( .A(n409), .B(n408), .C(n407), .Y(n410) );
  NAND2X1 U650 ( .A(n411), .B(n410), .Y(n416) );
  OAI22X1 U651 ( .A(n276), .B(n8), .C(n251), .D(n412), .Y(n414) );
  AOI21X1 U652 ( .A(currentPlainKey[5]), .B(n269), .C(n414), .Y(n415) );
  NAND2X1 U653 ( .A(n416), .B(n415), .Y(n1791) );
  NAND2X1 U654 ( .A(n417), .B(n280), .Y(n434) );
  NAND2X1 U655 ( .A(n177), .B(n205), .Y(n512) );
  NAND2X1 U656 ( .A(n220), .B(n186), .Y(n1556) );
  OAI21X1 U657 ( .A(n200), .B(n203), .C(currentPlainKey[6]), .Y(n418) );
  OAI21X1 U658 ( .A(n1556), .B(n203), .C(n418), .Y(n420) );
  NOR2X1 U659 ( .A(n273), .B(n512), .Y(n419) );
  AOI21X1 U660 ( .A(n133), .B(n420), .C(n419), .Y(n422) );
  NAND2X1 U661 ( .A(n483), .B(n282), .Y(n421) );
  OAI21X1 U662 ( .A(n497), .B(n422), .C(n421), .Y(n423) );
  NAND2X1 U663 ( .A(n229), .B(n423), .Y(n426) );
  NAND2X1 U664 ( .A(n497), .B(n245), .Y(n425) );
  AOI21X1 U665 ( .A(n426), .B(n425), .C(n424), .Y(n427) );
  MUX2X1 U666 ( .B(n427), .A(n262), .S(n121), .Y(n429) );
  NAND2X1 U667 ( .A(n463), .B(n254), .Y(n428) );
  NAND2X1 U668 ( .A(n429), .B(n428), .Y(n431) );
  MUX2X1 U669 ( .B(n431), .A(n246), .S(n430), .Y(n433) );
  NAND2X1 U670 ( .A(currentPlainKey[6]), .B(n268), .Y(n432) );
  NAND3X1 U671 ( .A(n434), .B(n433), .C(n432), .Y(n1792) );
  NAND2X1 U672 ( .A(n497), .B(n263), .Y(n442) );
  NAND2X1 U673 ( .A(n220), .B(n191), .Y(n572) );
  OAI21X1 U674 ( .A(n204), .B(n203), .C(currentPlainKey[7]), .Y(n435) );
  OAI21X1 U675 ( .A(n572), .B(n203), .C(n435), .Y(n436) );
  NAND3X1 U676 ( .A(n133), .B(n228), .C(n436), .Y(n437) );
  NAND2X1 U677 ( .A(n177), .B(n186), .Y(n546) );
  INVX2 U678 ( .A(n546), .Y(n517) );
  MUX2X1 U679 ( .B(n437), .A(n233), .S(n517), .Y(n439) );
  OAI22X1 U680 ( .A(n240), .B(n513), .C(n236), .D(n512), .Y(n438) );
  OAI21X1 U681 ( .A(n439), .B(n438), .C(n85), .Y(n441) );
  NAND2X1 U682 ( .A(n121), .B(n254), .Y(n440) );
  NAND3X1 U683 ( .A(n442), .B(n441), .C(n440), .Y(n443) );
  NAND2X1 U684 ( .A(n444), .B(n443), .Y(n449) );
  OAI22X1 U685 ( .A(n250), .B(n446), .C(n276), .D(n445), .Y(n447) );
  AOI21X1 U686 ( .A(currentPlainKey[7]), .B(n269), .C(n447), .Y(n448) );
  NAND2X1 U687 ( .A(n449), .B(n448), .Y(n1793) );
  NAND2X1 U688 ( .A(n121), .B(n279), .Y(n467) );
  INVX2 U689 ( .A(n512), .Y(n530) );
  NAND2X1 U690 ( .A(n177), .B(n191), .Y(n545) );
  NAND3X1 U691 ( .A(n222), .B(n1004), .C(n727), .Y(n571) );
  OAI21X1 U692 ( .A(n1142), .B(n209), .C(currentPlainKey[8]), .Y(n451) );
  OAI21X1 U693 ( .A(n1144), .B(n208), .C(n451), .Y(n453) );
  NOR2X1 U694 ( .A(n273), .B(n83), .Y(n452) );
  AOI21X1 U695 ( .A(n131), .B(n453), .C(n452), .Y(n455) );
  NAND2X1 U696 ( .A(n517), .B(n282), .Y(n454) );
  OAI21X1 U697 ( .A(n530), .B(n455), .C(n454), .Y(n456) );
  NAND2X1 U698 ( .A(n229), .B(n456), .Y(n459) );
  NAND2X1 U699 ( .A(n530), .B(n245), .Y(n458) );
  AOI21X1 U700 ( .A(n459), .B(n458), .C(n457), .Y(n460) );
  MUX2X1 U701 ( .B(n460), .A(n262), .S(n483), .Y(n462) );
  NAND2X1 U702 ( .A(n497), .B(n255), .Y(n461) );
  NAND2X1 U703 ( .A(n462), .B(n461), .Y(n464) );
  MUX2X1 U704 ( .B(n464), .A(n246), .S(n463), .Y(n466) );
  NAND2X1 U705 ( .A(currentPlainKey[8]), .B(n266), .Y(n465) );
  NAND3X1 U706 ( .A(n467), .B(n466), .C(n465), .Y(n1794) );
  NAND2X1 U707 ( .A(n530), .B(n263), .Y(n476) );
  OAI21X1 U708 ( .A(n196), .B(n209), .C(currentPlainKey[9]), .Y(n468) );
  OAI21X1 U709 ( .A(n469), .B(n208), .C(n468), .Y(n470) );
  NAND3X1 U710 ( .A(n131), .B(n228), .C(n470), .Y(n471) );
  NAND2X1 U711 ( .A(n586), .B(n178), .Y(n568) );
  MUX2X1 U712 ( .B(n471), .A(n233), .S(n53), .Y(n473) );
  OAI22X1 U713 ( .A(n240), .B(n546), .C(n238), .D(n83), .Y(n472) );
  OAI21X1 U714 ( .A(n473), .B(n472), .C(n133), .Y(n475) );
  NAND2X1 U715 ( .A(n483), .B(n255), .Y(n474) );
  NAND3X1 U716 ( .A(n476), .B(n475), .C(n474), .Y(n477) );
  NAND2X1 U717 ( .A(n85), .B(n477), .Y(n482) );
  OAI22X1 U718 ( .A(n251), .B(n479), .C(n275), .D(n87), .Y(n480) );
  AOI21X1 U719 ( .A(currentPlainKey[9]), .B(n266), .C(n480), .Y(n481) );
  NAND2X1 U720 ( .A(n481), .B(n482), .Y(n1795) );
  NAND2X1 U721 ( .A(n483), .B(n277), .Y(n501) );
  INVX2 U722 ( .A(n484), .Y(n1488) );
  NAND2X1 U723 ( .A(n586), .B(n1488), .Y(n567) );
  NAND2X1 U724 ( .A(n568), .B(n567), .Y(n570) );
  INVX2 U725 ( .A(n570), .Y(n538) );
  OAI21X1 U726 ( .A(n75), .B(n209), .C(currentPlainKey[10]), .Y(n485) );
  OAI21X1 U727 ( .A(n1179), .B(n208), .C(n485), .Y(n487) );
  NOR2X1 U728 ( .A(n273), .B(n567), .Y(n486) );
  AOI21X1 U729 ( .A(n538), .B(n487), .C(n486), .Y(n489) );
  NAND2X1 U730 ( .A(n550), .B(n282), .Y(n488) );
  OAI21X1 U731 ( .A(n562), .B(n489), .C(n488), .Y(n490) );
  NAND2X1 U732 ( .A(n229), .B(n490), .Y(n493) );
  NAND2X1 U733 ( .A(n562), .B(n245), .Y(n492) );
  AOI21X1 U734 ( .A(n493), .B(n492), .C(n491), .Y(n494) );
  MUX2X1 U735 ( .B(n494), .A(n262), .S(n517), .Y(n496) );
  NAND2X1 U736 ( .A(n530), .B(n255), .Y(n495) );
  NAND2X1 U737 ( .A(n496), .B(n495), .Y(n498) );
  MUX2X1 U738 ( .B(n498), .A(n246), .S(n497), .Y(n500) );
  NAND2X1 U739 ( .A(currentPlainKey[10]), .B(n266), .Y(n499) );
  NAND3X1 U740 ( .A(n501), .B(n500), .C(n499), .Y(n1796) );
  NAND2X1 U741 ( .A(n562), .B(n262), .Y(n510) );
  OAI21X1 U742 ( .A(n202), .B(n209), .C(currentPlainKey[11]), .Y(n502) );
  OAI21X1 U743 ( .A(n503), .B(n208), .C(n502), .Y(n504) );
  NAND3X1 U744 ( .A(n538), .B(n228), .C(n504), .Y(n505) );
  NAND2X1 U745 ( .A(n586), .B(n174), .Y(n604) );
  MUX2X1 U746 ( .B(n505), .A(n233), .S(n585), .Y(n507) );
  OAI22X1 U747 ( .A(n240), .B(n568), .C(n236), .D(n57), .Y(n506) );
  OAI21X1 U748 ( .A(n507), .B(n506), .C(n81), .Y(n509) );
  NAND2X1 U749 ( .A(n517), .B(n253), .Y(n508) );
  NAND3X1 U750 ( .A(n510), .B(n509), .C(n508), .Y(n511) );
  NAND2X1 U751 ( .A(n133), .B(n511), .Y(n516) );
  OAI22X1 U752 ( .A(n249), .B(n513), .C(n276), .D(n512), .Y(n514) );
  AOI21X1 U753 ( .A(currentPlainKey[11]), .B(n268), .C(n514), .Y(n515) );
  NAND2X1 U754 ( .A(n516), .B(n515), .Y(n1797) );
  NAND2X1 U755 ( .A(n517), .B(n278), .Y(n534) );
  INVX2 U756 ( .A(n567), .Y(n598) );
  NAND2X1 U757 ( .A(n586), .B(n175), .Y(n603) );
  OAI21X1 U758 ( .A(n71), .B(n209), .C(currentPlainKey[12]), .Y(n518) );
  OAI21X1 U759 ( .A(n1521), .B(n208), .C(n518), .Y(n520) );
  NOR2X1 U760 ( .A(n273), .B(n603), .Y(n519) );
  AOI21X1 U761 ( .A(n123), .B(n520), .C(n519), .Y(n522) );
  NAND2X1 U762 ( .A(n585), .B(n282), .Y(n521) );
  OAI21X1 U763 ( .A(n522), .B(n598), .C(n521), .Y(n523) );
  NAND2X1 U764 ( .A(n229), .B(n523), .Y(n526) );
  NAND2X1 U765 ( .A(n598), .B(n245), .Y(n525) );
  AOI21X1 U766 ( .A(n526), .B(n525), .C(n524), .Y(n527) );
  MUX2X1 U767 ( .B(n527), .A(n262), .S(n53), .Y(n529) );
  NAND2X1 U768 ( .A(n562), .B(n255), .Y(n528) );
  NAND2X1 U769 ( .A(n529), .B(n528), .Y(n531) );
  MUX2X1 U770 ( .B(n531), .A(n246), .S(n530), .Y(n533) );
  NAND2X1 U771 ( .A(currentPlainKey[12]), .B(n270), .Y(n532) );
  NAND3X1 U772 ( .A(n534), .B(n533), .C(n532), .Y(n1798) );
  NAND2X1 U773 ( .A(n598), .B(n263), .Y(n543) );
  OAI21X1 U774 ( .A(n206), .B(n209), .C(currentPlainKey[13]), .Y(n535) );
  OAI21X1 U775 ( .A(n1544), .B(n208), .C(n535), .Y(n536) );
  NAND3X1 U776 ( .A(n123), .B(n228), .C(n536), .Y(n537) );
  NAND2X1 U777 ( .A(n586), .B(n157), .Y(n638) );
  INVX2 U778 ( .A(n638), .Y(n620) );
  MUX2X1 U779 ( .B(n537), .A(n233), .S(n620), .Y(n540) );
  OAI22X1 U780 ( .A(n240), .B(n101), .C(n16), .D(n19), .Y(n539) );
  OAI21X1 U781 ( .A(n540), .B(n539), .C(n538), .Y(n542) );
  NAND2X1 U782 ( .A(n53), .B(n255), .Y(n541) );
  NAND3X1 U783 ( .A(n543), .B(n542), .C(n541), .Y(n544) );
  NAND2X1 U784 ( .A(n81), .B(n544), .Y(n549) );
  OAI22X1 U785 ( .A(n249), .B(n546), .C(n276), .D(n83), .Y(n547) );
  AOI21X1 U786 ( .A(currentPlainKey[13]), .B(n268), .C(n547), .Y(n548) );
  NAND2X1 U787 ( .A(n548), .B(n549), .Y(n1799) );
  NAND2X1 U788 ( .A(n53), .B(n279), .Y(n566) );
  NAND2X1 U789 ( .A(n586), .B(n176), .Y(n637) );
  OAI21X1 U790 ( .A(n199), .B(n209), .C(currentPlainKey[14]), .Y(n551) );
  OAI21X1 U791 ( .A(n1556), .B(n208), .C(n551), .Y(n553) );
  NOR2X1 U792 ( .A(n272), .B(n637), .Y(n552) );
  AOI21X1 U793 ( .A(n150), .B(n553), .C(n552), .Y(n555) );
  NAND2X1 U794 ( .A(n620), .B(n282), .Y(n554) );
  OAI21X1 U795 ( .A(n632), .B(n555), .C(n554), .Y(n556) );
  NAND2X1 U796 ( .A(n229), .B(n556), .Y(n558) );
  NAND2X1 U797 ( .A(n632), .B(n245), .Y(n557) );
  AOI21X1 U798 ( .A(n558), .B(n557), .C(n570), .Y(n559) );
  MUX2X1 U799 ( .B(n559), .A(n262), .S(n585), .Y(n561) );
  NAND2X1 U800 ( .A(n598), .B(n255), .Y(n560) );
  NAND2X1 U801 ( .A(n561), .B(n560), .Y(n563) );
  MUX2X1 U802 ( .B(n563), .A(n246), .S(n562), .Y(n565) );
  NAND2X1 U803 ( .A(currentPlainKey[14]), .B(n266), .Y(n564) );
  NAND3X1 U804 ( .A(n566), .B(n565), .C(n564), .Y(n1800) );
  OAI22X1 U805 ( .A(n249), .B(n568), .C(n276), .D(n57), .Y(n569) );
  AOI21X1 U806 ( .A(currentPlainKey[15]), .B(n266), .C(n569), .Y(n584) );
  OAI21X1 U807 ( .A(n204), .B(n209), .C(currentPlainKey[15]), .Y(n575) );
  INVX2 U808 ( .A(n208), .Y(n573) );
  INVX2 U809 ( .A(n572), .Y(n1430) );
  NAND2X1 U810 ( .A(n573), .B(n1430), .Y(n574) );
  NAND2X1 U811 ( .A(n575), .B(n574), .Y(n576) );
  NAND3X1 U812 ( .A(n228), .B(n576), .C(n653), .Y(n577) );
  NAND2X1 U813 ( .A(n586), .B(n1130), .Y(n673) );
  MUX2X1 U814 ( .B(n577), .A(n233), .S(n656), .Y(n579) );
  OAI22X1 U815 ( .A(n240), .B(n638), .C(n16), .D(n637), .Y(n578) );
  OAI21X1 U816 ( .A(n579), .B(n578), .C(n123), .Y(n581) );
  AOI22X1 U817 ( .A(n632), .B(n260), .C(n585), .D(n253), .Y(n580) );
  NAND2X1 U818 ( .A(n581), .B(n580), .Y(n582) );
  NAND2X1 U819 ( .A(n538), .B(n582), .Y(n583) );
  NAND2X1 U820 ( .A(n584), .B(n583), .Y(n1801) );
  NAND2X1 U821 ( .A(n585), .B(n277), .Y(n602) );
  NAND2X1 U822 ( .A(n586), .B(n179), .Y(n672) );
  NAND3X1 U823 ( .A(address[4]), .B(n221), .C(n727), .Y(n712) );
  OAI21X1 U824 ( .A(n1142), .B(n211), .C(currentPlainKey[16]), .Y(n587) );
  OAI21X1 U825 ( .A(n1144), .B(n211), .C(n587), .Y(n589) );
  NOR2X1 U826 ( .A(n272), .B(n672), .Y(n588) );
  AOI21X1 U827 ( .A(n141), .B(n589), .C(n588), .Y(n591) );
  NAND2X1 U828 ( .A(n656), .B(n282), .Y(n590) );
  OAI21X1 U829 ( .A(n614), .B(n591), .C(n590), .Y(n592) );
  NAND2X1 U830 ( .A(n229), .B(n592), .Y(n594) );
  NAND2X1 U831 ( .A(n614), .B(n245), .Y(n593) );
  AOI21X1 U832 ( .A(n594), .B(n593), .C(n606), .Y(n595) );
  MUX2X1 U833 ( .B(n595), .A(n262), .S(n620), .Y(n597) );
  NAND2X1 U834 ( .A(n632), .B(n255), .Y(n596) );
  NAND2X1 U835 ( .A(n597), .B(n596), .Y(n599) );
  MUX2X1 U836 ( .B(n599), .A(n246), .S(n598), .Y(n601) );
  NAND2X1 U837 ( .A(currentPlainKey[16]), .B(n268), .Y(n600) );
  NAND3X1 U838 ( .A(n602), .B(n601), .C(n600), .Y(n1802) );
  OAI22X1 U839 ( .A(n250), .B(n101), .C(n276), .D(n19), .Y(n605) );
  AOI21X1 U840 ( .A(currentPlainKey[17]), .B(n266), .C(n605), .Y(n619) );
  OAI21X1 U841 ( .A(n196), .B(n211), .C(currentPlainKey[17]), .Y(n608) );
  INVX2 U842 ( .A(n211), .Y(n713) );
  NAND2X1 U843 ( .A(n713), .B(n1470), .Y(n607) );
  NAND2X1 U844 ( .A(n608), .B(n607), .Y(n609) );
  NAND3X1 U845 ( .A(n227), .B(n609), .C(n688), .Y(n611) );
  NAND3X1 U846 ( .A(n79), .B(address[4]), .C(n727), .Y(n610) );
  NAND2X1 U847 ( .A(n183), .B(n47), .Y(n709) );
  INVX2 U848 ( .A(n709), .Y(n691) );
  MUX2X1 U849 ( .B(n611), .A(n233), .S(n691), .Y(n613) );
  OAI22X1 U850 ( .A(n240), .B(n25), .C(n238), .D(n55), .Y(n612) );
  OAI21X1 U851 ( .A(n613), .B(n612), .C(n653), .Y(n616) );
  AOI22X1 U852 ( .A(n614), .B(n260), .C(n620), .D(n253), .Y(n615) );
  NAND2X1 U853 ( .A(n616), .B(n615), .Y(n617) );
  NAND2X1 U854 ( .A(n123), .B(n617), .Y(n618) );
  NAND2X1 U855 ( .A(n619), .B(n618), .Y(n1803) );
  NAND2X1 U856 ( .A(n620), .B(n279), .Y(n636) );
  NAND2X1 U857 ( .A(n183), .B(n195), .Y(n708) );
  NAND2X1 U858 ( .A(n709), .B(n708), .Y(n711) );
  OAI21X1 U859 ( .A(n75), .B(n211), .C(currentPlainKey[18]), .Y(n621) );
  OAI21X1 U860 ( .A(n1179), .B(n211), .C(n621), .Y(n623) );
  NOR2X1 U861 ( .A(n272), .B(n29), .Y(n622) );
  AOI21X1 U862 ( .A(n681), .B(n623), .C(n622), .Y(n625) );
  NAND2X1 U863 ( .A(n691), .B(n282), .Y(n624) );
  OAI21X1 U864 ( .A(n703), .B(n625), .C(n624), .Y(n626) );
  NAND2X1 U865 ( .A(n229), .B(n626), .Y(n628) );
  NAND2X1 U866 ( .A(n703), .B(n245), .Y(n627) );
  AOI21X1 U867 ( .A(n628), .B(n627), .C(n640), .Y(n629) );
  MUX2X1 U868 ( .B(n629), .A(n262), .S(n656), .Y(n631) );
  NAND2X1 U869 ( .A(n614), .B(n255), .Y(n630) );
  NAND2X1 U870 ( .A(n631), .B(n630), .Y(n633) );
  MUX2X1 U871 ( .B(n633), .A(n246), .S(n632), .Y(n635) );
  NAND2X1 U872 ( .A(currentPlainKey[18]), .B(n268), .Y(n634) );
  NAND3X1 U873 ( .A(n636), .B(n635), .C(n634), .Y(n1804) );
  OAI22X1 U874 ( .A(n250), .B(n638), .C(n276), .D(n637), .Y(n639) );
  AOI21X1 U875 ( .A(currentPlainKey[19]), .B(n266), .C(n639), .Y(n655) );
  OAI21X1 U876 ( .A(n202), .B(n211), .C(currentPlainKey[19]), .Y(n642) );
  NAND2X1 U877 ( .A(n713), .B(n1357), .Y(n641) );
  NAND2X1 U878 ( .A(n642), .B(n641), .Y(n644) );
  NAND3X1 U879 ( .A(n228), .B(n644), .C(n643), .Y(n645) );
  NAND2X1 U880 ( .A(n183), .B(n159), .Y(n745) );
  INVX2 U881 ( .A(n745), .Y(n726) );
  MUX2X1 U882 ( .B(n645), .A(n233), .S(n726), .Y(n647) );
  OAI22X1 U883 ( .A(n240), .B(n709), .C(n238), .D(n29), .Y(n646) );
  OAI21X1 U884 ( .A(n647), .B(n646), .C(n688), .Y(n651) );
  AOI22X1 U885 ( .A(n649), .B(n260), .C(n648), .D(n253), .Y(n650) );
  NAND2X1 U886 ( .A(n651), .B(n650), .Y(n652) );
  NAND2X1 U887 ( .A(n653), .B(n652), .Y(n654) );
  NAND2X1 U888 ( .A(n655), .B(n654), .Y(n1805) );
  NAND2X1 U889 ( .A(n656), .B(n277), .Y(n671) );
  NAND2X1 U890 ( .A(n183), .B(n201), .Y(n744) );
  OAI21X1 U891 ( .A(n71), .B(n211), .C(currentPlainKey[20]), .Y(n657) );
  OAI21X1 U892 ( .A(n1521), .B(n211), .C(n657), .Y(n659) );
  NOR2X1 U893 ( .A(n272), .B(n744), .Y(n658) );
  AOI21X1 U894 ( .A(n97), .B(n659), .C(n658), .Y(n661) );
  NAND2X1 U895 ( .A(n726), .B(n281), .Y(n660) );
  OAI21X1 U896 ( .A(n661), .B(n739), .C(n660), .Y(n662) );
  NAND2X1 U897 ( .A(n229), .B(n662), .Y(n664) );
  NAND2X1 U898 ( .A(n739), .B(n245), .Y(n663) );
  AOI21X1 U899 ( .A(n664), .B(n663), .C(n675), .Y(n665) );
  NAND2X1 U900 ( .A(n703), .B(n255), .Y(n666) );
  NAND2X1 U901 ( .A(n667), .B(n666), .Y(n668) );
  MUX2X1 U902 ( .B(n668), .A(n246), .S(n614), .Y(n670) );
  NAND2X1 U903 ( .A(currentPlainKey[20]), .B(n269), .Y(n669) );
  NAND3X1 U904 ( .A(n671), .B(n670), .C(n669), .Y(n1806) );
  OAI22X1 U905 ( .A(n250), .B(n25), .C(n275), .D(n55), .Y(n674) );
  AOI21X1 U906 ( .A(currentPlainKey[21]), .B(n268), .C(n674), .Y(n690) );
  OAI21X1 U907 ( .A(n206), .B(n211), .C(currentPlainKey[21]), .Y(n677) );
  INVX2 U908 ( .A(n1544), .Y(n1393) );
  NAND2X1 U909 ( .A(n713), .B(n1393), .Y(n676) );
  NAND2X1 U910 ( .A(n677), .B(n676), .Y(n679) );
  NAND3X1 U911 ( .A(n228), .B(n679), .C(n678), .Y(n680) );
  NAND2X1 U912 ( .A(n183), .B(n1520), .Y(n780) );
  INVX2 U913 ( .A(n780), .Y(n762) );
  MUX2X1 U914 ( .B(n680), .A(n233), .S(n762), .Y(n683) );
  OAI22X1 U915 ( .A(n240), .B(n745), .C(n16), .D(n744), .Y(n682) );
  OAI21X1 U916 ( .A(n683), .B(n682), .C(n681), .Y(n686) );
  AOI22X1 U917 ( .A(n684), .B(n260), .C(n691), .D(n253), .Y(n685) );
  NAND2X1 U918 ( .A(n686), .B(n685), .Y(n687) );
  NAND2X1 U919 ( .A(n688), .B(n687), .Y(n689) );
  NAND2X1 U920 ( .A(n690), .B(n689), .Y(n1807) );
  NAND2X1 U921 ( .A(n691), .B(n280), .Y(n707) );
  NAND2X1 U922 ( .A(n183), .B(n205), .Y(n779) );
  NAND2X1 U923 ( .A(n780), .B(n779), .Y(n782) );
  OAI21X1 U924 ( .A(n200), .B(n211), .C(currentPlainKey[22]), .Y(n692) );
  OAI21X1 U925 ( .A(n1556), .B(n211), .C(n692), .Y(n694) );
  NOR2X1 U926 ( .A(n272), .B(n37), .Y(n693) );
  AOI21X1 U927 ( .A(n753), .B(n694), .C(n693), .Y(n696) );
  NAND2X1 U928 ( .A(n762), .B(n281), .Y(n695) );
  OAI21X1 U929 ( .A(n774), .B(n696), .C(n695), .Y(n697) );
  NAND2X1 U930 ( .A(n229), .B(n697), .Y(n699) );
  NAND2X1 U931 ( .A(n774), .B(n243), .Y(n698) );
  AOI21X1 U932 ( .A(n699), .B(n698), .C(n711), .Y(n700) );
  MUX2X1 U933 ( .B(n700), .A(n262), .S(n726), .Y(n702) );
  NAND2X1 U934 ( .A(n739), .B(n255), .Y(n701) );
  NAND2X1 U935 ( .A(n702), .B(n701), .Y(n704) );
  MUX2X1 U936 ( .B(n704), .A(n248), .S(n703), .Y(n706) );
  NAND2X1 U937 ( .A(currentPlainKey[22]), .B(n266), .Y(n705) );
  NAND3X1 U938 ( .A(n707), .B(n706), .C(n705), .Y(n1808) );
  OAI22X1 U939 ( .A(n251), .B(n709), .C(n276), .D(n29), .Y(n710) );
  AOI21X1 U940 ( .A(currentPlainKey[23]), .B(n270), .C(n710), .Y(n725) );
  OAI21X1 U941 ( .A(n204), .B(n211), .C(currentPlainKey[23]), .Y(n715) );
  NAND2X1 U942 ( .A(n713), .B(n1430), .Y(n714) );
  NAND2X1 U943 ( .A(n715), .B(n714), .Y(n717) );
  NAND3X1 U944 ( .A(n228), .B(n717), .C(n716), .Y(n718) );
  NAND2X1 U945 ( .A(n183), .B(n186), .Y(n815) );
  INVX2 U946 ( .A(n815), .Y(n797) );
  MUX2X1 U947 ( .B(n718), .A(n233), .S(n797), .Y(n720) );
  OAI22X1 U948 ( .A(n240), .B(n780), .C(n238), .D(n37), .Y(n719) );
  OAI21X1 U949 ( .A(n720), .B(n719), .C(n678), .Y(n722) );
  AOI22X1 U950 ( .A(n774), .B(n260), .C(n726), .D(n253), .Y(n721) );
  NAND2X1 U951 ( .A(n722), .B(n721), .Y(n723) );
  NAND2X1 U952 ( .A(n643), .B(n723), .Y(n724) );
  NAND2X1 U953 ( .A(n725), .B(n724), .Y(n1809) );
  NAND2X1 U954 ( .A(n726), .B(n278), .Y(n743) );
  NAND2X1 U955 ( .A(n183), .B(n191), .Y(n814) );
  NAND2X1 U956 ( .A(n815), .B(n814), .Y(n817) );
  INVX2 U957 ( .A(n817), .Y(n788) );
  NAND3X1 U958 ( .A(n222), .B(address[4]), .C(n727), .Y(n850) );
  OAI21X1 U959 ( .A(n1142), .B(n213), .C(currentPlainKey[24]), .Y(n728) );
  OAI21X1 U960 ( .A(n1144), .B(n213), .C(n728), .Y(n730) );
  NOR2X1 U961 ( .A(n272), .B(n31), .Y(n729) );
  AOI21X1 U962 ( .A(n788), .B(n730), .C(n729), .Y(n732) );
  NAND2X1 U963 ( .A(n797), .B(n281), .Y(n731) );
  OAI21X1 U964 ( .A(n809), .B(n732), .C(n731), .Y(n733) );
  NAND2X1 U965 ( .A(n229), .B(n733), .Y(n735) );
  NAND2X1 U966 ( .A(n809), .B(n242), .Y(n734) );
  AOI21X1 U967 ( .A(n735), .B(n734), .C(n747), .Y(n736) );
  MUX2X1 U968 ( .B(n736), .A(n261), .S(n762), .Y(n738) );
  NAND2X1 U969 ( .A(n774), .B(n253), .Y(n737) );
  NAND2X1 U970 ( .A(n738), .B(n737), .Y(n740) );
  MUX2X1 U971 ( .B(n740), .A(n248), .S(n739), .Y(n742) );
  NAND2X1 U972 ( .A(currentPlainKey[24]), .B(n266), .Y(n741) );
  NAND3X1 U973 ( .A(n743), .B(n742), .C(n741), .Y(n1810) );
  OAI22X1 U974 ( .A(n251), .B(n745), .C(n276), .D(n744), .Y(n746) );
  AOI21X1 U975 ( .A(currentPlainKey[25]), .B(n266), .C(n746), .Y(n761) );
  OAI21X1 U976 ( .A(n196), .B(n213), .C(currentPlainKey[25]), .Y(n749) );
  INVX2 U977 ( .A(n213), .Y(n851) );
  NAND2X1 U978 ( .A(n851), .B(n1470), .Y(n748) );
  NAND2X1 U979 ( .A(n749), .B(n748), .Y(n751) );
  NAND3X1 U980 ( .A(n228), .B(n751), .C(n750), .Y(n752) );
  NAND2X1 U981 ( .A(n158), .B(n178), .Y(n847) );
  MUX2X1 U982 ( .B(n752), .A(n233), .S(n824), .Y(n755) );
  OAI22X1 U983 ( .A(n240), .B(n815), .C(n237), .D(n31), .Y(n754) );
  OAI21X1 U984 ( .A(n755), .B(n754), .C(n753), .Y(n758) );
  AOI22X1 U985 ( .A(n756), .B(n260), .C(n762), .D(n253), .Y(n757) );
  NAND2X1 U986 ( .A(n758), .B(n757), .Y(n759) );
  NAND2X1 U987 ( .A(n678), .B(n759), .Y(n760) );
  NAND2X1 U988 ( .A(n761), .B(n760), .Y(n1811) );
  NAND2X1 U989 ( .A(n762), .B(n279), .Y(n778) );
  NAND2X1 U990 ( .A(n158), .B(n1488), .Y(n846) );
  OAI21X1 U991 ( .A(n75), .B(n213), .C(currentPlainKey[26]), .Y(n763) );
  OAI21X1 U992 ( .A(n1179), .B(n213), .C(n763), .Y(n765) );
  NOR2X1 U993 ( .A(n272), .B(n846), .Y(n764) );
  AOI21X1 U994 ( .A(n137), .B(n765), .C(n764), .Y(n767) );
  NAND2X1 U995 ( .A(n824), .B(n281), .Y(n766) );
  OAI21X1 U996 ( .A(n841), .B(n767), .C(n766), .Y(n768) );
  NAND2X1 U997 ( .A(n229), .B(n768), .Y(n770) );
  NAND2X1 U998 ( .A(n841), .B(n243), .Y(n769) );
  AOI21X1 U999 ( .A(n770), .B(n769), .C(n782), .Y(n771) );
  MUX2X1 U1000 ( .B(n771), .A(n262), .S(n797), .Y(n773) );
  NAND2X1 U1001 ( .A(n809), .B(n254), .Y(n772) );
  NAND2X1 U1002 ( .A(n773), .B(n772), .Y(n775) );
  MUX2X1 U1003 ( .B(n775), .A(n248), .S(n774), .Y(n777) );
  NAND2X1 U1004 ( .A(currentPlainKey[26]), .B(n268), .Y(n776) );
  NAND3X1 U1005 ( .A(n778), .B(n777), .C(n776), .Y(n1812) );
  OAI22X1 U1006 ( .A(n251), .B(n780), .C(n276), .D(n37), .Y(n781) );
  AOI21X1 U1007 ( .A(currentPlainKey[27]), .B(n268), .C(n781), .Y(n796) );
  OAI21X1 U1008 ( .A(n202), .B(n213), .C(currentPlainKey[27]), .Y(n784) );
  NAND2X1 U1009 ( .A(n851), .B(n1357), .Y(n783) );
  NAND2X1 U1010 ( .A(n784), .B(n783), .Y(n786) );
  NAND3X1 U1011 ( .A(n228), .B(n786), .C(n785), .Y(n787) );
  NAND2X1 U1012 ( .A(n158), .B(n174), .Y(n882) );
  INVX2 U1013 ( .A(n882), .Y(n863) );
  MUX2X1 U1014 ( .B(n787), .A(n233), .S(n863), .Y(n790) );
  OAI22X1 U1015 ( .A(n240), .B(n847), .C(n238), .D(n846), .Y(n789) );
  OAI21X1 U1016 ( .A(n790), .B(n789), .C(n788), .Y(n793) );
  AOI22X1 U1017 ( .A(n791), .B(n260), .C(n797), .D(n253), .Y(n792) );
  NAND2X1 U1018 ( .A(n793), .B(n792), .Y(n794) );
  NAND2X1 U1019 ( .A(n716), .B(n794), .Y(n795) );
  NAND2X1 U1020 ( .A(n796), .B(n795), .Y(n1813) );
  NAND2X1 U1021 ( .A(n797), .B(n277), .Y(n813) );
  INVX2 U1022 ( .A(n846), .Y(n876) );
  NAND2X1 U1023 ( .A(n158), .B(n175), .Y(n881) );
  OAI21X1 U1024 ( .A(n71), .B(n213), .C(currentPlainKey[28]), .Y(n798) );
  OAI21X1 U1025 ( .A(n1521), .B(n213), .C(n798), .Y(n800) );
  NOR2X1 U1026 ( .A(n272), .B(n881), .Y(n799) );
  AOI21X1 U1027 ( .A(n139), .B(n800), .C(n799), .Y(n802) );
  NAND2X1 U1028 ( .A(n863), .B(n281), .Y(n801) );
  OAI21X1 U1029 ( .A(n802), .B(n876), .C(n801), .Y(n803) );
  NAND2X1 U1030 ( .A(n229), .B(n803), .Y(n805) );
  NAND2X1 U1031 ( .A(n876), .B(n243), .Y(n804) );
  AOI21X1 U1032 ( .A(n805), .B(n804), .C(n817), .Y(n806) );
  MUX2X1 U1033 ( .B(n806), .A(n261), .S(n824), .Y(n808) );
  NAND2X1 U1034 ( .A(n841), .B(n253), .Y(n807) );
  NAND2X1 U1035 ( .A(n808), .B(n807), .Y(n810) );
  MUX2X1 U1036 ( .B(n810), .A(n247), .S(n809), .Y(n812) );
  NAND2X1 U1037 ( .A(currentPlainKey[28]), .B(n266), .Y(n811) );
  NAND3X1 U1038 ( .A(n813), .B(n812), .C(n811), .Y(n1814) );
  OAI22X1 U1039 ( .A(n251), .B(n815), .C(n276), .D(n31), .Y(n816) );
  AOI21X1 U1040 ( .A(currentPlainKey[29]), .B(n268), .C(n816), .Y(n829) );
  OAI21X1 U1041 ( .A(n206), .B(n213), .C(currentPlainKey[29]), .Y(n819) );
  NAND2X1 U1042 ( .A(n851), .B(n1393), .Y(n818) );
  NAND2X1 U1043 ( .A(n819), .B(n818), .Y(n820) );
  NAND3X1 U1044 ( .A(n227), .B(n820), .C(n896), .Y(n821) );
  NAND2X1 U1045 ( .A(n158), .B(n173), .Y(n916) );
  MUX2X1 U1046 ( .B(n821), .A(n234), .S(n892), .Y(n823) );
  OAI22X1 U1047 ( .A(n240), .B(n882), .C(n238), .D(n11), .Y(n822) );
  OAI21X1 U1048 ( .A(n823), .B(n822), .C(n785), .Y(n826) );
  AOI22X1 U1049 ( .A(n876), .B(n260), .C(n824), .D(n253), .Y(n825) );
  NAND2X1 U1050 ( .A(n826), .B(n825), .Y(n827) );
  NAND2X1 U1051 ( .A(n750), .B(n827), .Y(n828) );
  NAND2X1 U1052 ( .A(n829), .B(n828), .Y(n1815) );
  NAND2X1 U1053 ( .A(n824), .B(n279), .Y(n845) );
  NAND2X1 U1054 ( .A(n158), .B(n176), .Y(n915) );
  OAI21X1 U1055 ( .A(n200), .B(n213), .C(currentPlainKey[30]), .Y(n830) );
  OAI21X1 U1056 ( .A(n1556), .B(n213), .C(n830), .Y(n832) );
  NOR2X1 U1057 ( .A(n272), .B(n915), .Y(n831) );
  AOI21X1 U1058 ( .A(n149), .B(n832), .C(n831), .Y(n834) );
  NAND2X1 U1059 ( .A(n892), .B(n281), .Y(n833) );
  OAI21X1 U1060 ( .A(n834), .B(n910), .C(n833), .Y(n835) );
  NAND2X1 U1061 ( .A(n229), .B(n835), .Y(n837) );
  NAND2X1 U1062 ( .A(n910), .B(n244), .Y(n836) );
  AOI21X1 U1063 ( .A(n837), .B(n836), .C(n849), .Y(n838) );
  MUX2X1 U1064 ( .B(n838), .A(n261), .S(n863), .Y(n840) );
  NAND2X1 U1065 ( .A(n876), .B(n253), .Y(n839) );
  NAND2X1 U1066 ( .A(n840), .B(n839), .Y(n842) );
  MUX2X1 U1067 ( .B(n842), .A(n247), .S(n841), .Y(n844) );
  NAND2X1 U1068 ( .A(currentPlainKey[30]), .B(n268), .Y(n843) );
  NAND3X1 U1069 ( .A(n845), .B(n844), .C(n843), .Y(n1816) );
  OAI22X1 U1070 ( .A(n251), .B(n847), .C(n275), .D(n846), .Y(n848) );
  AOI21X1 U1071 ( .A(currentPlainKey[31]), .B(n267), .C(n848), .Y(n862) );
  OAI21X1 U1072 ( .A(n204), .B(n213), .C(currentPlainKey[31]), .Y(n853) );
  NAND2X1 U1073 ( .A(n851), .B(n1430), .Y(n852) );
  NAND2X1 U1074 ( .A(n853), .B(n852), .Y(n854) );
  NAND3X1 U1075 ( .A(n228), .B(n854), .C(n931), .Y(n855) );
  NAND2X1 U1076 ( .A(n158), .B(n1130), .Y(n952) );
  INVX2 U1077 ( .A(n952), .Y(n934) );
  MUX2X1 U1078 ( .B(n855), .A(n234), .S(n934), .Y(n857) );
  OAI22X1 U1079 ( .A(n240), .B(n916), .C(n237), .D(n6), .Y(n856) );
  OAI21X1 U1080 ( .A(n857), .B(n856), .C(n896), .Y(n859) );
  AOI22X1 U1081 ( .A(n910), .B(n259), .C(n863), .D(n252), .Y(n858) );
  NAND2X1 U1082 ( .A(n859), .B(n858), .Y(n860) );
  NAND2X1 U1083 ( .A(n785), .B(n860), .Y(n861) );
  NAND2X1 U1084 ( .A(n862), .B(n861), .Y(n1817) );
  NAND2X1 U1085 ( .A(n863), .B(n280), .Y(n880) );
  INVX2 U1086 ( .A(n915), .Y(n946) );
  NAND2X1 U1087 ( .A(n158), .B(n179), .Y(n951) );
  NAND3X1 U1088 ( .A(address[5]), .B(n221), .C(n1004), .Y(n989) );
  OAI21X1 U1089 ( .A(n1142), .B(n215), .C(currentPlainKey[32]), .Y(n865) );
  OAI21X1 U1090 ( .A(n1144), .B(n215), .C(n865), .Y(n867) );
  NOR2X1 U1091 ( .A(n272), .B(n951), .Y(n866) );
  AOI21X1 U1092 ( .A(n153), .B(n867), .C(n866), .Y(n869) );
  NAND2X1 U1093 ( .A(n934), .B(n281), .Y(n868) );
  OAI21X1 U1094 ( .A(n946), .B(n869), .C(n868), .Y(n870) );
  NAND2X1 U1095 ( .A(n229), .B(n870), .Y(n872) );
  NAND2X1 U1096 ( .A(n946), .B(n243), .Y(n871) );
  AOI21X1 U1097 ( .A(n872), .B(n871), .C(n884), .Y(n873) );
  MUX2X1 U1098 ( .B(n873), .A(n261), .S(n892), .Y(n875) );
  NAND2X1 U1099 ( .A(n910), .B(n253), .Y(n874) );
  NAND2X1 U1100 ( .A(n875), .B(n874), .Y(n877) );
  MUX2X1 U1101 ( .B(n877), .A(n247), .S(n876), .Y(n879) );
  NAND2X1 U1102 ( .A(currentPlainKey[32]), .B(n266), .Y(n878) );
  NAND3X1 U1103 ( .A(n880), .B(n879), .C(n878), .Y(n1818) );
  OAI22X1 U1104 ( .A(n251), .B(n93), .C(n275), .D(n11), .Y(n883) );
  AOI21X1 U1105 ( .A(currentPlainKey[33]), .B(n267), .C(n883), .Y(n898) );
  OAI21X1 U1106 ( .A(n196), .B(n215), .C(currentPlainKey[33]), .Y(n886) );
  INVX2 U1107 ( .A(n215), .Y(n990) );
  NAND2X1 U1108 ( .A(n990), .B(n1470), .Y(n885) );
  NAND2X1 U1109 ( .A(n886), .B(n885), .Y(n887) );
  NAND3X1 U1110 ( .A(n227), .B(n887), .C(n965), .Y(n889) );
  NAND3X1 U1111 ( .A(n79), .B(address[5]), .C(n1004), .Y(n888) );
  NAND2X1 U1112 ( .A(n182), .B(n47), .Y(n986) );
  INVX2 U1113 ( .A(n986), .Y(n968) );
  MUX2X1 U1114 ( .B(n889), .A(n234), .S(n968), .Y(n891) );
  OAI22X1 U1115 ( .A(n239), .B(n45), .C(n16), .D(n41), .Y(n890) );
  OAI21X1 U1116 ( .A(n891), .B(n890), .C(n931), .Y(n894) );
  AOI22X1 U1117 ( .A(n946), .B(n259), .C(n892), .D(n252), .Y(n893) );
  NAND2X1 U1118 ( .A(n894), .B(n893), .Y(n895) );
  NAND2X1 U1119 ( .A(n896), .B(n895), .Y(n897) );
  NAND2X1 U1120 ( .A(n898), .B(n897), .Y(n1819) );
  NAND2X1 U1121 ( .A(n892), .B(n279), .Y(n914) );
  NAND2X1 U1122 ( .A(n182), .B(n195), .Y(n985) );
  NAND2X1 U1123 ( .A(n986), .B(n985), .Y(n988) );
  INVX2 U1124 ( .A(n988), .Y(n959) );
  OAI21X1 U1125 ( .A(n75), .B(n215), .C(currentPlainKey[34]), .Y(n899) );
  OAI21X1 U1126 ( .A(n1179), .B(n215), .C(n899), .Y(n901) );
  NOR2X1 U1127 ( .A(n272), .B(n33), .Y(n900) );
  AOI21X1 U1128 ( .A(n959), .B(n901), .C(n900), .Y(n903) );
  NAND2X1 U1129 ( .A(n968), .B(n281), .Y(n902) );
  OAI21X1 U1130 ( .A(n980), .B(n903), .C(n902), .Y(n904) );
  NAND2X1 U1131 ( .A(n229), .B(n904), .Y(n906) );
  NAND2X1 U1132 ( .A(n980), .B(n243), .Y(n905) );
  AOI21X1 U1133 ( .A(n906), .B(n905), .C(n918), .Y(n907) );
  MUX2X1 U1134 ( .B(n907), .A(n261), .S(n934), .Y(n909) );
  NAND2X1 U1135 ( .A(n946), .B(n254), .Y(n908) );
  NAND2X1 U1136 ( .A(n909), .B(n908), .Y(n911) );
  MUX2X1 U1137 ( .B(n911), .A(n247), .S(n910), .Y(n913) );
  NAND2X1 U1138 ( .A(currentPlainKey[34]), .B(n268), .Y(n912) );
  NAND3X1 U1139 ( .A(n914), .B(n913), .C(n912), .Y(n1820) );
  OAI22X1 U1140 ( .A(n251), .B(n916), .C(n275), .D(n6), .Y(n917) );
  AOI21X1 U1141 ( .A(currentPlainKey[35]), .B(n269), .C(n917), .Y(n933) );
  OAI21X1 U1142 ( .A(n202), .B(n215), .C(currentPlainKey[35]), .Y(n920) );
  NAND2X1 U1143 ( .A(n990), .B(n1357), .Y(n919) );
  NAND2X1 U1144 ( .A(n920), .B(n919), .Y(n922) );
  NAND3X1 U1145 ( .A(n228), .B(n922), .C(n921), .Y(n923) );
  NAND2X1 U1146 ( .A(n182), .B(n159), .Y(n1022) );
  INVX2 U1147 ( .A(n1022), .Y(n1003) );
  MUX2X1 U1148 ( .B(n923), .A(n234), .S(n1003), .Y(n925) );
  OAI22X1 U1149 ( .A(n239), .B(n986), .C(n237), .D(n33), .Y(n924) );
  OAI21X1 U1150 ( .A(n925), .B(n924), .C(n965), .Y(n929) );
  AOI22X1 U1151 ( .A(n927), .B(n259), .C(n926), .D(n252), .Y(n928) );
  NAND2X1 U1152 ( .A(n929), .B(n928), .Y(n930) );
  NAND2X1 U1153 ( .A(n931), .B(n930), .Y(n932) );
  NAND2X1 U1154 ( .A(n933), .B(n932), .Y(n1821) );
  NAND2X1 U1155 ( .A(n934), .B(n277), .Y(n950) );
  NAND2X1 U1156 ( .A(n182), .B(n201), .Y(n1021) );
  OAI21X1 U1157 ( .A(n71), .B(n215), .C(currentPlainKey[36]), .Y(n935) );
  OAI21X1 U1158 ( .A(n1521), .B(n215), .C(n935), .Y(n937) );
  NOR2X1 U1159 ( .A(n272), .B(n1021), .Y(n936) );
  AOI21X1 U1160 ( .A(n99), .B(n937), .C(n936), .Y(n939) );
  NAND2X1 U1161 ( .A(n1003), .B(n281), .Y(n938) );
  OAI21X1 U1162 ( .A(n1016), .B(n939), .C(n938), .Y(n940) );
  NAND2X1 U1163 ( .A(n229), .B(n940), .Y(n942) );
  NAND2X1 U1164 ( .A(n1016), .B(n243), .Y(n941) );
  AOI21X1 U1165 ( .A(n942), .B(n941), .C(n954), .Y(n943) );
  NAND2X1 U1166 ( .A(n980), .B(n254), .Y(n944) );
  NAND2X1 U1167 ( .A(n944), .B(n945), .Y(n947) );
  MUX2X1 U1168 ( .B(n947), .A(n247), .S(n946), .Y(n949) );
  NAND2X1 U1169 ( .A(currentPlainKey[36]), .B(n270), .Y(n948) );
  NAND3X1 U1170 ( .A(n950), .B(n949), .C(n948), .Y(n1822) );
  OAI22X1 U1171 ( .A(n251), .B(n45), .C(n275), .D(n41), .Y(n953) );
  AOI21X1 U1172 ( .A(currentPlainKey[37]), .B(n270), .C(n953), .Y(n967) );
  OAI21X1 U1173 ( .A(n206), .B(n215), .C(currentPlainKey[37]), .Y(n956) );
  NAND2X1 U1174 ( .A(n990), .B(n1393), .Y(n955) );
  NAND2X1 U1175 ( .A(n956), .B(n955), .Y(n957) );
  NAND3X1 U1176 ( .A(n227), .B(n957), .C(n1036), .Y(n958) );
  NAND2X1 U1177 ( .A(n182), .B(n1520), .Y(n1057) );
  INVX2 U1178 ( .A(n1057), .Y(n1039) );
  MUX2X1 U1179 ( .B(n958), .A(n234), .S(n1039), .Y(n961) );
  OAI22X1 U1180 ( .A(n239), .B(n1022), .C(n237), .D(n1021), .Y(n960) );
  OAI21X1 U1181 ( .A(n961), .B(n960), .C(n959), .Y(n963) );
  AOI22X1 U1182 ( .A(n1016), .B(n259), .C(n968), .D(n252), .Y(n962) );
  NAND2X1 U1183 ( .A(n963), .B(n962), .Y(n964) );
  NAND2X1 U1184 ( .A(n965), .B(n964), .Y(n966) );
  NAND2X1 U1185 ( .A(n967), .B(n966), .Y(n1823) );
  NAND2X1 U1186 ( .A(n968), .B(n280), .Y(n984) );
  NAND2X1 U1187 ( .A(n182), .B(n205), .Y(n1056) );
  NAND2X1 U1188 ( .A(n1057), .B(n1056), .Y(n1059) );
  INVX2 U1189 ( .A(n1059), .Y(n1029) );
  OAI21X1 U1190 ( .A(n199), .B(n215), .C(currentPlainKey[38]), .Y(n969) );
  OAI21X1 U1191 ( .A(n1556), .B(n215), .C(n969), .Y(n971) );
  NOR2X1 U1192 ( .A(n272), .B(n39), .Y(n970) );
  AOI21X1 U1193 ( .A(n1029), .B(n971), .C(n970), .Y(n973) );
  NAND2X1 U1194 ( .A(n1039), .B(n281), .Y(n972) );
  OAI21X1 U1195 ( .A(n1051), .B(n973), .C(n972), .Y(n974) );
  NAND2X1 U1196 ( .A(n229), .B(n974), .Y(n976) );
  NAND2X1 U1197 ( .A(n1051), .B(n244), .Y(n975) );
  AOI21X1 U1198 ( .A(n976), .B(n975), .C(n988), .Y(n977) );
  MUX2X1 U1199 ( .B(n977), .A(n261), .S(n1003), .Y(n979) );
  NAND2X1 U1200 ( .A(n1016), .B(n254), .Y(n978) );
  NAND2X1 U1201 ( .A(n979), .B(n978), .Y(n981) );
  MUX2X1 U1202 ( .B(n981), .A(n247), .S(n980), .Y(n983) );
  NAND2X1 U1203 ( .A(currentPlainKey[38]), .B(n268), .Y(n982) );
  NAND3X1 U1204 ( .A(n984), .B(n983), .C(n982), .Y(n1824) );
  OAI22X1 U1205 ( .A(n250), .B(n986), .C(n275), .D(n33), .Y(n987) );
  AOI21X1 U1206 ( .A(currentPlainKey[39]), .B(n269), .C(n987), .Y(n1002) );
  OAI21X1 U1207 ( .A(n204), .B(n215), .C(currentPlainKey[39]), .Y(n992) );
  NAND2X1 U1208 ( .A(n990), .B(n1430), .Y(n991) );
  NAND2X1 U1209 ( .A(n992), .B(n991), .Y(n994) );
  NAND3X1 U1210 ( .A(n227), .B(n994), .C(n993), .Y(n995) );
  NAND2X1 U1211 ( .A(n182), .B(n186), .Y(n1090) );
  INVX2 U1212 ( .A(n1090), .Y(n1072) );
  MUX2X1 U1213 ( .B(n995), .A(n234), .S(n1072), .Y(n997) );
  OAI22X1 U1214 ( .A(n239), .B(n1057), .C(n238), .D(n39), .Y(n996) );
  OAI21X1 U1215 ( .A(n997), .B(n996), .C(n1036), .Y(n999) );
  AOI22X1 U1216 ( .A(n1051), .B(n259), .C(n1003), .D(n252), .Y(n998) );
  NAND2X1 U1217 ( .A(n999), .B(n998), .Y(n1000) );
  NAND2X1 U1218 ( .A(n921), .B(n1000), .Y(n1001) );
  NAND2X1 U1219 ( .A(n1002), .B(n1001), .Y(n1825) );
  NAND2X1 U1220 ( .A(n1003), .B(n277), .Y(n1020) );
  NAND2X1 U1221 ( .A(n182), .B(n191), .Y(n1089) );
  NAND3X1 U1222 ( .A(n222), .B(address[5]), .C(n1004), .Y(n1125) );
  OAI21X1 U1223 ( .A(n1142), .B(n217), .C(currentPlainKey[40]), .Y(n1005) );
  OAI21X1 U1224 ( .A(n1144), .B(n217), .C(n1005), .Y(n1007) );
  NOR2X1 U1225 ( .A(n272), .B(n1089), .Y(n1006) );
  AOI21X1 U1226 ( .A(n95), .B(n1007), .C(n1006), .Y(n1009) );
  NAND2X1 U1227 ( .A(n1072), .B(n281), .Y(n1008) );
  OAI21X1 U1228 ( .A(n1084), .B(n1009), .C(n1008), .Y(n1010) );
  NAND2X1 U1229 ( .A(n229), .B(n1010), .Y(n1012) );
  NAND2X1 U1230 ( .A(n1084), .B(n244), .Y(n1011) );
  AOI21X1 U1231 ( .A(n1012), .B(n1011), .C(n1024), .Y(n1013) );
  NAND2X1 U1232 ( .A(n1051), .B(n254), .Y(n1014) );
  NAND2X1 U1233 ( .A(n1014), .B(n1015), .Y(n1017) );
  MUX2X1 U1234 ( .B(n1017), .A(n247), .S(n1016), .Y(n1019) );
  NAND2X1 U1235 ( .A(currentPlainKey[40]), .B(n266), .Y(n1018) );
  NAND3X1 U1236 ( .A(n1020), .B(n1019), .C(n1018), .Y(n1826) );
  OAI22X1 U1237 ( .A(n250), .B(n1022), .C(n275), .D(n1021), .Y(n1023) );
  AOI21X1 U1238 ( .A(currentPlainKey[41]), .B(n266), .C(n1023), .Y(n1038) );
  OAI21X1 U1239 ( .A(n196), .B(n217), .C(currentPlainKey[41]), .Y(n1026) );
  INVX2 U1240 ( .A(n217), .Y(n1126) );
  NAND2X1 U1241 ( .A(n1126), .B(n1470), .Y(n1025) );
  NAND2X1 U1242 ( .A(n1026), .B(n1025), .Y(n1027) );
  NAND3X1 U1243 ( .A(n227), .B(n1027), .C(n1102), .Y(n1028) );
  NAND2X1 U1244 ( .A(n1141), .B(n178), .Y(n1122) );
  MUX2X1 U1245 ( .B(n1028), .A(n234), .S(n1105), .Y(n1031) );
  OAI22X1 U1246 ( .A(n239), .B(n1090), .C(n16), .D(n1089), .Y(n1030) );
  OAI21X1 U1247 ( .A(n1031), .B(n1030), .C(n1029), .Y(n1034) );
  AOI22X1 U1248 ( .A(n1032), .B(n259), .C(n1039), .D(n252), .Y(n1033) );
  NAND2X1 U1249 ( .A(n1034), .B(n1033), .Y(n1035) );
  NAND2X1 U1250 ( .A(n1036), .B(n1035), .Y(n1037) );
  NAND2X1 U1251 ( .A(n1038), .B(n1037), .Y(n1827) );
  NAND2X1 U1252 ( .A(n1039), .B(n278), .Y(n1055) );
  NAND2X1 U1253 ( .A(n1141), .B(n1488), .Y(n1121) );
  OAI21X1 U1254 ( .A(n75), .B(n217), .C(currentPlainKey[42]), .Y(n1040) );
  OAI21X1 U1255 ( .A(n1179), .B(n217), .C(n1040), .Y(n1042) );
  NOR2X1 U1256 ( .A(n272), .B(n1121), .Y(n1041) );
  AOI21X1 U1257 ( .A(n127), .B(n1042), .C(n1041), .Y(n1044) );
  NAND2X1 U1258 ( .A(n1105), .B(n281), .Y(n1043) );
  OAI21X1 U1259 ( .A(n1066), .B(n1044), .C(n1043), .Y(n1045) );
  NAND2X1 U1260 ( .A(n229), .B(n1045), .Y(n1047) );
  NAND2X1 U1261 ( .A(n1066), .B(n244), .Y(n1046) );
  AOI21X1 U1262 ( .A(n1047), .B(n1046), .C(n1059), .Y(n1048) );
  MUX2X1 U1263 ( .B(n1048), .A(n261), .S(n1072), .Y(n1050) );
  NAND2X1 U1264 ( .A(n1084), .B(n254), .Y(n1049) );
  NAND2X1 U1265 ( .A(n1050), .B(n1049), .Y(n1052) );
  NAND2X1 U1266 ( .A(currentPlainKey[42]), .B(n268), .Y(n1053) );
  NAND3X1 U1267 ( .A(n1055), .B(n1053), .C(n1054), .Y(n1828) );
  OAI22X1 U1268 ( .A(n250), .B(n1057), .C(n275), .D(n39), .Y(n1058) );
  AOI21X1 U1269 ( .A(currentPlainKey[43]), .B(n268), .C(n1058), .Y(n1071) );
  OAI21X1 U1270 ( .A(n202), .B(n217), .C(currentPlainKey[43]), .Y(n1061) );
  NAND2X1 U1271 ( .A(n1126), .B(n1357), .Y(n1060) );
  NAND2X1 U1272 ( .A(n1061), .B(n1060), .Y(n1062) );
  NAND3X1 U1273 ( .A(n227), .B(n1062), .C(n1137), .Y(n1063) );
  NAND2X1 U1274 ( .A(n1141), .B(n174), .Y(n1161) );
  INVX2 U1275 ( .A(n1161), .Y(n1140) );
  MUX2X1 U1276 ( .B(n1063), .A(n234), .S(n1140), .Y(n1065) );
  OAI22X1 U1277 ( .A(n239), .B(n1122), .C(n16), .D(n9), .Y(n1064) );
  OAI21X1 U1278 ( .A(n1065), .B(n1064), .C(n1102), .Y(n1068) );
  INVX2 U1279 ( .A(n1089), .Y(n1066) );
  AOI22X1 U1280 ( .A(n1066), .B(n259), .C(n1072), .D(n252), .Y(n1067) );
  NAND2X1 U1281 ( .A(n1068), .B(n1067), .Y(n1069) );
  NAND2X1 U1282 ( .A(n993), .B(n1069), .Y(n1070) );
  NAND2X1 U1283 ( .A(n1071), .B(n1070), .Y(n1829) );
  NAND2X1 U1284 ( .A(n1072), .B(n280), .Y(n1088) );
  NAND2X1 U1285 ( .A(n1141), .B(n175), .Y(n1160) );
  OAI21X1 U1286 ( .A(n71), .B(n217), .C(currentPlainKey[44]), .Y(n1073) );
  OAI21X1 U1287 ( .A(n1521), .B(n217), .C(n1073), .Y(n1075) );
  NOR2X1 U1288 ( .A(n271), .B(n1160), .Y(n1074) );
  AOI21X1 U1289 ( .A(n135), .B(n1075), .C(n1074), .Y(n1077) );
  NAND2X1 U1290 ( .A(n1140), .B(n281), .Y(n1076) );
  OAI21X1 U1291 ( .A(n1077), .B(n1155), .C(n1076), .Y(n1078) );
  NAND2X1 U1292 ( .A(n229), .B(n1078), .Y(n1080) );
  NAND2X1 U1293 ( .A(n1155), .B(n244), .Y(n1079) );
  AOI21X1 U1294 ( .A(n1080), .B(n1079), .C(n1092), .Y(n1081) );
  MUX2X1 U1295 ( .B(n1081), .A(n261), .S(n1105), .Y(n1083) );
  NAND2X1 U1296 ( .A(n1066), .B(n254), .Y(n1082) );
  NAND2X1 U1297 ( .A(n1083), .B(n1082), .Y(n1085) );
  MUX2X1 U1298 ( .B(n1085), .A(n247), .S(n1084), .Y(n1087) );
  NAND2X1 U1299 ( .A(currentPlainKey[44]), .B(n266), .Y(n1086) );
  NAND3X1 U1300 ( .A(n1088), .B(n1087), .C(n1086), .Y(n1830) );
  OAI22X1 U1301 ( .A(n251), .B(n1090), .C(n275), .D(n1089), .Y(n1091) );
  AOI21X1 U1302 ( .A(currentPlainKey[45]), .B(n266), .C(n1091), .Y(n1104) );
  OAI21X1 U1303 ( .A(n206), .B(n217), .C(currentPlainKey[45]), .Y(n1094) );
  NAND2X1 U1304 ( .A(n1126), .B(n1393), .Y(n1093) );
  NAND2X1 U1306 ( .A(n1094), .B(n1093), .Y(n1095) );
  NAND3X1 U1307 ( .A(n227), .B(n1095), .C(n135), .Y(n1096) );
  NAND2X1 U1308 ( .A(n1141), .B(n173), .Y(n1196) );
  INVX2 U1309 ( .A(n1196), .Y(n1175) );
  MUX2X1 U1310 ( .B(n1096), .A(n234), .S(n1175), .Y(n1098) );
  OAI22X1 U1311 ( .A(n239), .B(n1161), .C(n16), .D(n10), .Y(n1097) );
  OAI21X1 U1312 ( .A(n1098), .B(n1097), .C(n1137), .Y(n1100) );
  AOI22X1 U1313 ( .A(n1155), .B(n259), .C(n1105), .D(n252), .Y(n1099) );
  NAND2X1 U1314 ( .A(n1100), .B(n1099), .Y(n1101) );
  NAND2X1 U1315 ( .A(n1102), .B(n1101), .Y(n1103) );
  NAND2X1 U1316 ( .A(n1104), .B(n1103), .Y(n1831) );
  NAND2X1 U1317 ( .A(n1105), .B(n280), .Y(n1120) );
  NAND2X1 U1318 ( .A(n1141), .B(n176), .Y(n1195) );
  OAI21X1 U1319 ( .A(n199), .B(n217), .C(currentPlainKey[46]), .Y(n1106) );
  OAI21X1 U1320 ( .A(n1556), .B(n217), .C(n1106), .Y(n1108) );
  NOR2X1 U1321 ( .A(n271), .B(n1195), .Y(n1107) );
  AOI21X1 U1322 ( .A(n154), .B(n1108), .C(n1107), .Y(n1110) );
  NAND2X1 U1323 ( .A(n1175), .B(n281), .Y(n1109) );
  OAI21X1 U1324 ( .A(n1110), .B(n1190), .C(n1109), .Y(n1111) );
  NAND2X1 U1325 ( .A(n229), .B(n1111), .Y(n1113) );
  NAND2X1 U1326 ( .A(n1190), .B(n245), .Y(n1112) );
  AOI21X1 U1327 ( .A(n1113), .B(n1112), .C(n1124), .Y(n1114) );
  MUX2X1 U1328 ( .B(n1114), .A(n261), .S(n1140), .Y(n1116) );
  NAND2X1 U1329 ( .A(n1155), .B(n254), .Y(n1115) );
  NAND2X1 U1330 ( .A(n1116), .B(n1115), .Y(n1117) );
  MUX2X1 U1331 ( .B(n1117), .A(n246), .S(n1066), .Y(n1119) );
  NAND2X1 U1332 ( .A(currentPlainKey[46]), .B(n268), .Y(n1118) );
  NAND3X1 U1333 ( .A(n1120), .B(n1119), .C(n1118), .Y(n1832) );
  OAI22X1 U1334 ( .A(n249), .B(n1122), .C(n276), .D(n9), .Y(n1123) );
  AOI21X1 U1335 ( .A(currentPlainKey[47]), .B(n268), .C(n1123), .Y(n1139) );
  OAI21X1 U1336 ( .A(n204), .B(n217), .C(currentPlainKey[47]), .Y(n1128) );
  NAND2X1 U1337 ( .A(n1126), .B(n1430), .Y(n1127) );
  NAND2X1 U1338 ( .A(n1128), .B(n1127), .Y(n1129) );
  NAND3X1 U1339 ( .A(n227), .B(n1129), .C(n1368), .Y(n1131) );
  NAND2X1 U1340 ( .A(n1141), .B(n1130), .Y(n1390) );
  INVX2 U1341 ( .A(n1390), .Y(n1371) );
  MUX2X1 U1342 ( .B(n1131), .A(n234), .S(n1371), .Y(n1133) );
  OAI22X1 U1343 ( .A(n239), .B(n89), .C(n237), .D(n59), .Y(n1132) );
  OAI21X1 U1344 ( .A(n1133), .B(n1132), .C(n135), .Y(n1135) );
  AOI22X1 U1345 ( .A(n1190), .B(n259), .C(n1140), .D(n252), .Y(n1134) );
  NAND2X1 U1346 ( .A(n1135), .B(n1134), .Y(n1136) );
  NAND2X1 U1347 ( .A(n1137), .B(n1136), .Y(n1138) );
  NAND2X1 U1348 ( .A(n1139), .B(n1138), .Y(n1833) );
  NAND2X1 U1349 ( .A(n1140), .B(n279), .Y(n1159) );
  NAND2X1 U1350 ( .A(n1141), .B(n179), .Y(n1389) );
  OAI21X1 U1351 ( .A(n1142), .B(n218), .C(currentPlainKey[48]), .Y(n1143) );
  OAI21X1 U1358 ( .A(n1144), .B(n218), .C(n1143), .Y(n1146) );
  NOR2X1 U1359 ( .A(n271), .B(n1389), .Y(n1145) );
  AOI21X1 U1360 ( .A(n145), .B(n1146), .C(n1145), .Y(n1148) );
  NAND2X1 U1361 ( .A(n1371), .B(n281), .Y(n1147) );
  OAI21X1 U1362 ( .A(n1384), .B(n1148), .C(n1147), .Y(n1149) );
  NAND2X1 U1363 ( .A(n229), .B(n1149), .Y(n1151) );
  NAND2X1 U1364 ( .A(n1384), .B(n245), .Y(n1150) );
  AOI21X1 U1365 ( .A(n1151), .B(n1150), .C(n1163), .Y(n1152) );
  MUX2X1 U1366 ( .B(n1152), .A(n261), .S(n1175), .Y(n1154) );
  NAND2X1 U1367 ( .A(n1190), .B(n254), .Y(n1153) );
  NAND2X1 U1368 ( .A(n1154), .B(n1153), .Y(n1156) );
  MUX2X1 U1369 ( .B(n1156), .A(n248), .S(n1155), .Y(n1158) );
  NAND2X1 U1370 ( .A(currentPlainKey[48]), .B(n268), .Y(n1157) );
  NAND3X1 U1371 ( .A(n1159), .B(n1158), .C(n1157), .Y(n1834) );
  OAI22X1 U1372 ( .A(n251), .B(n1161), .C(n275), .D(n10), .Y(n1162) );
  AOI21X1 U1373 ( .A(currentPlainKey[49]), .B(n270), .C(n1162), .Y(n1174) );
  OAI21X1 U1374 ( .A(n196), .B(n218), .C(currentPlainKey[49]), .Y(n1165) );
  INVX2 U1375 ( .A(n218), .Y(n1429) );
  NAND2X1 U1376 ( .A(n1429), .B(n1470), .Y(n1164) );
  NAND2X1 U1377 ( .A(n1165), .B(n1164), .Y(n1166) );
  NAND3X1 U1378 ( .A(n227), .B(n1166), .C(n1404), .Y(n1167) );
  NAND2X1 U1379 ( .A(n79), .B(n188), .Y(n1582) );
  NAND2X1 U1380 ( .A(n169), .B(n47), .Y(n1425) );
  INVX2 U1381 ( .A(n1425), .Y(n1407) );
  MUX2X1 U1382 ( .B(n1167), .A(n234), .S(n1407), .Y(n1169) );
  OAI22X1 U1383 ( .A(n239), .B(n20), .C(n16), .D(n51), .Y(n1168) );
  OAI21X1 U1384 ( .A(n1169), .B(n1168), .C(n1368), .Y(n1171) );
  AOI22X1 U1385 ( .A(n1384), .B(n259), .C(n1175), .D(n252), .Y(n1170) );
  NAND2X1 U1386 ( .A(n1171), .B(n1170), .Y(n1172) );
  NAND2X1 U1387 ( .A(n135), .B(n1172), .Y(n1173) );
  NAND2X1 U1388 ( .A(n1174), .B(n1173), .Y(n1835) );
  NAND2X1 U1389 ( .A(n1175), .B(n278), .Y(n1194) );
  NAND2X1 U1390 ( .A(n169), .B(n195), .Y(n1424) );
  OAI21X1 U1391 ( .A(n75), .B(n218), .C(currentPlainKey[50]), .Y(n1177) );
  OAI21X1 U1392 ( .A(n1179), .B(n218), .C(n1177), .Y(n1181) );
  NOR2X1 U1393 ( .A(n271), .B(n1424), .Y(n1180) );
  AOI21X1 U1394 ( .A(n129), .B(n1181), .C(n1180), .Y(n1183) );
  NAND2X1 U1395 ( .A(n1407), .B(n281), .Y(n1182) );
  OAI21X1 U1396 ( .A(n1419), .B(n1183), .C(n1182), .Y(n1184) );
  NAND2X1 U1397 ( .A(n229), .B(n1184), .Y(n1186) );
  NAND2X1 U1398 ( .A(n1419), .B(n242), .Y(n1185) );
  AOI21X1 U1399 ( .A(n1186), .B(n1185), .C(n1268), .Y(n1187) );
  MUX2X1 U1400 ( .B(n1187), .A(n260), .S(n1371), .Y(n1189) );
  NAND2X1 U1401 ( .A(n1384), .B(n254), .Y(n1188) );
  NAND2X1 U1402 ( .A(n1189), .B(n1188), .Y(n1191) );
  MUX2X1 U1403 ( .B(n1191), .A(n248), .S(n1190), .Y(n1193) );
  NAND2X1 U1404 ( .A(currentPlainKey[50]), .B(n270), .Y(n1192) );
  NAND3X1 U1405 ( .A(n1194), .B(n1193), .C(n1192), .Y(n1836) );
  OAI22X1 U1406 ( .A(n251), .B(n89), .C(n275), .D(n59), .Y(n1267) );
  AOI21X1 U1407 ( .A(currentPlainKey[51]), .B(n269), .C(n1267), .Y(n1370) );
  OAI21X1 U1408 ( .A(n202), .B(n218), .C(currentPlainKey[51]), .Y(n1359) );
  NAND2X1 U1409 ( .A(n1357), .B(n1429), .Y(n1358) );
  NAND2X1 U1410 ( .A(n1359), .B(n1358), .Y(n1360) );
  NAND3X1 U1411 ( .A(n227), .B(n1360), .C(n1441), .Y(n1361) );
  NAND2X1 U1412 ( .A(n169), .B(n159), .Y(n1481) );
  MUX2X1 U1413 ( .B(n1361), .A(n234), .S(n1444), .Y(n1363) );
  OAI22X1 U1414 ( .A(n239), .B(n43), .C(n237), .D(n21), .Y(n1362) );
  OAI21X1 U1415 ( .A(n1363), .B(n1362), .C(n1404), .Y(n1366) );
  AOI22X1 U1416 ( .A(n1419), .B(n259), .C(n1364), .D(n252), .Y(n1365) );
  NAND2X1 U1417 ( .A(n1366), .B(n1365), .Y(n1367) );
  NAND2X1 U1418 ( .A(n1368), .B(n1367), .Y(n1369) );
  NAND2X1 U1419 ( .A(n1370), .B(n1369), .Y(n1837) );
  NAND2X1 U1420 ( .A(n1371), .B(n278), .Y(n1388) );
  NAND2X1 U1421 ( .A(n169), .B(n201), .Y(n1480) );
  OAI21X1 U1422 ( .A(n71), .B(n218), .C(currentPlainKey[52]), .Y(n1373) );
  OAI21X1 U1423 ( .A(n1521), .B(n218), .C(n1373), .Y(n1375) );
  NOR2X1 U1424 ( .A(n271), .B(n1480), .Y(n1374) );
  AOI21X1 U1425 ( .A(n147), .B(n1375), .C(n1374), .Y(n1377) );
  NAND2X1 U1426 ( .A(n1444), .B(n281), .Y(n1376) );
  OAI21X1 U1427 ( .A(n1460), .B(n1377), .C(n1376), .Y(n1378) );
  NAND2X1 U1428 ( .A(n229), .B(n1378), .Y(n1380) );
  NAND2X1 U1429 ( .A(n1460), .B(n242), .Y(n1379) );
  AOI21X1 U1430 ( .A(n1380), .B(n1379), .C(n1392), .Y(n1381) );
  MUX2X1 U1431 ( .B(n1381), .A(n260), .S(n1407), .Y(n1383) );
  NAND2X1 U1432 ( .A(n1419), .B(n254), .Y(n1382) );
  NAND2X1 U1433 ( .A(n1383), .B(n1382), .Y(n1385) );
  MUX2X1 U1434 ( .B(n1385), .A(n248), .S(n1384), .Y(n1387) );
  NAND2X1 U1435 ( .A(currentPlainKey[52]), .B(n269), .Y(n1386) );
  NAND3X1 U1436 ( .A(n1388), .B(n1387), .C(n1386), .Y(n1838) );
  OAI22X1 U1437 ( .A(n251), .B(n20), .C(n275), .D(n51), .Y(n1391) );
  AOI21X1 U1438 ( .A(currentPlainKey[53]), .B(n267), .C(n1391), .Y(n1406) );
  OAI21X1 U1439 ( .A(n206), .B(n218), .C(currentPlainKey[53]), .Y(n1395) );
  NAND2X1 U1440 ( .A(n1429), .B(n1393), .Y(n1394) );
  NAND2X1 U1441 ( .A(n1395), .B(n1394), .Y(n1396) );
  NAND3X1 U1442 ( .A(n227), .B(n1396), .C(n147), .Y(n1397) );
  NAND2X1 U1443 ( .A(n169), .B(n1520), .Y(n1465) );
  INVX2 U1444 ( .A(n1465), .Y(n1515) );
  MUX2X1 U1445 ( .B(n1397), .A(n235), .S(n1515), .Y(n1399) );
  OAI22X1 U1446 ( .A(n239), .B(n27), .C(n238), .D(n65), .Y(n1398) );
  OAI21X1 U1447 ( .A(n1399), .B(n1398), .C(n1441), .Y(n1402) );
  AOI22X1 U1448 ( .A(n1400), .B(n259), .C(n1407), .D(n252), .Y(n1401) );
  NAND2X1 U1449 ( .A(n1402), .B(n1401), .Y(n1403) );
  NAND2X1 U1450 ( .A(n1404), .B(n1403), .Y(n1405) );
  NAND2X1 U1451 ( .A(n1406), .B(n1405), .Y(n1839) );
  NAND2X1 U1452 ( .A(n1407), .B(n278), .Y(n1423) );
  NAND2X1 U1453 ( .A(n169), .B(n205), .Y(n1453) );
  OAI21X1 U1454 ( .A(n199), .B(n218), .C(currentPlainKey[54]), .Y(n1408) );
  OAI21X1 U1455 ( .A(n218), .B(n1556), .C(n1408), .Y(n1410) );
  NOR2X1 U1456 ( .A(n271), .B(n1453), .Y(n1409) );
  AOI21X1 U1457 ( .A(n119), .B(n1410), .C(n1409), .Y(n1412) );
  NAND2X1 U1458 ( .A(n1515), .B(n281), .Y(n1411) );
  OAI21X1 U1459 ( .A(n1437), .B(n1412), .C(n1411), .Y(n1413) );
  NAND2X1 U1460 ( .A(n229), .B(n1413), .Y(n1415) );
  NAND2X1 U1461 ( .A(n1437), .B(n242), .Y(n1414) );
  AOI21X1 U1462 ( .A(n1415), .B(n1414), .C(n1427), .Y(n1416) );
  MUX2X1 U1463 ( .B(n1416), .A(n260), .S(n1444), .Y(n1418) );
  NAND2X1 U1464 ( .A(n1460), .B(n254), .Y(n1417) );
  NAND2X1 U1465 ( .A(n1418), .B(n1417), .Y(n1420) );
  MUX2X1 U1466 ( .B(n1420), .A(n248), .S(n1419), .Y(n1422) );
  NAND2X1 U1467 ( .A(currentPlainKey[54]), .B(n268), .Y(n1421) );
  NAND3X1 U1468 ( .A(n1423), .B(n1422), .C(n1421), .Y(n1840) );
  OAI22X1 U1469 ( .A(n251), .B(n43), .C(n275), .D(n21), .Y(n1426) );
  AOI21X1 U1470 ( .A(currentPlainKey[55]), .B(n268), .C(n1426), .Y(n1443) );
  OAI21X1 U1471 ( .A(n204), .B(n218), .C(currentPlainKey[55]), .Y(n1432) );
  NAND2X1 U1472 ( .A(n1430), .B(n1429), .Y(n1431) );
  NAND2X1 U1473 ( .A(n1432), .B(n1431), .Y(n1433) );
  NAND3X1 U1474 ( .A(n227), .B(n1433), .C(n119), .Y(n1434) );
  NAND2X1 U1475 ( .A(n169), .B(n186), .Y(n1504) );
  INVX2 U1476 ( .A(n1504), .Y(n1552) );
  MUX2X1 U1477 ( .B(n1434), .A(n235), .S(n1552), .Y(n1436) );
  OAI22X1 U1478 ( .A(n5), .B(n239), .C(n1453), .D(n237), .Y(n1435) );
  OAI21X1 U1479 ( .A(n1436), .B(n1435), .C(n147), .Y(n1439) );
  AOI22X1 U1480 ( .A(n1437), .B(n259), .C(n1444), .D(n252), .Y(n1438) );
  NAND2X1 U1481 ( .A(n1439), .B(n1438), .Y(n1440) );
  NAND2X1 U1482 ( .A(n1441), .B(n1440), .Y(n1442) );
  NAND2X1 U1483 ( .A(n1443), .B(n1442), .Y(n1841) );
  NAND2X1 U1484 ( .A(n1444), .B(n280), .Y(n1464) );
  NAND2X1 U1485 ( .A(n1552), .B(n281), .Y(n1451) );
  NAND2X1 U1486 ( .A(n223), .B(n188), .Y(n1578) );
  NAND2X1 U1487 ( .A(n1557), .B(n47), .Y(n1446) );
  AOI22X1 U1488 ( .A(currentPlainKey[56]), .B(n1446), .C(n1445), .D(n1557), 
        .Y(n1448) );
  NAND2X1 U1489 ( .A(n169), .B(n191), .Y(n1503) );
  NAND2X1 U1490 ( .A(n1504), .B(n1503), .Y(n1467) );
  NAND2X1 U1491 ( .A(n1571), .B(RCV_DATA[1]), .Y(n1447) );
  OAI21X1 U1492 ( .A(n1448), .B(n1467), .C(n1447), .Y(n1449) );
  NAND2X1 U1493 ( .A(n1449), .B(n1453), .Y(n1450) );
  NAND2X1 U1494 ( .A(n1451), .B(n1450), .Y(n1452) );
  NAND2X1 U1495 ( .A(n229), .B(n1452), .Y(n1456) );
  NAND2X1 U1496 ( .A(n244), .B(n1534), .Y(n1455) );
  AOI21X1 U1497 ( .A(n1456), .B(n1455), .C(n1454), .Y(n1457) );
  MUX2X1 U1498 ( .B(n1457), .A(n260), .S(n1515), .Y(n1459) );
  NAND2X1 U1499 ( .A(n1437), .B(n254), .Y(n1458) );
  NAND2X1 U1500 ( .A(n1459), .B(n1458), .Y(n1461) );
  MUX2X1 U1501 ( .B(n1461), .A(n248), .S(n1460), .Y(n1463) );
  NAND2X1 U1502 ( .A(currentPlainKey[56]), .B(n267), .Y(n1462) );
  NOR2X1 U1503 ( .A(n257), .B(n5), .Y(n1479) );
  OAI22X1 U1504 ( .A(n7), .B(n167), .C(n63), .D(n236), .Y(n1475) );
  NAND2X1 U1505 ( .A(n1561), .B(n178), .Y(n1529) );
  INVX2 U1506 ( .A(n1467), .Y(n1468) );
  NOR2X1 U1507 ( .A(n111), .B(n113), .Y(n1474) );
  OAI21X1 U1508 ( .A(n196), .B(n61), .C(currentPlainKey[57]), .Y(n1472) );
  NAND2X1 U1509 ( .A(n1470), .B(n1557), .Y(n1471) );
  NAND2X1 U1510 ( .A(n168), .B(n1529), .Y(n1519) );
  AOI21X1 U1511 ( .A(n1472), .B(n1471), .C(n1519), .Y(n1473) );
  NOR3X1 U1512 ( .A(n1473), .B(n1474), .C(n1475), .Y(n1477) );
  NAND2X1 U1513 ( .A(n1534), .B(n262), .Y(n1476) );
  OAI21X1 U1514 ( .A(n1493), .B(n1477), .C(n1476), .Y(n1478) );
  OAI21X1 U1515 ( .A(n1479), .B(n1478), .C(n147), .Y(n1485) );
  OAI22X1 U1516 ( .A(n251), .B(n27), .C(n275), .D(n65), .Y(n1483) );
  AOI21X1 U1517 ( .A(currentPlainKey[57]), .B(n266), .C(n1483), .Y(n1484) );
  NAND2X1 U1518 ( .A(n1485), .B(n1484), .Y(n1843) );
  NAND2X1 U1519 ( .A(n1515), .B(n279), .Y(n1502) );
  NAND2X1 U1520 ( .A(n244), .B(n1571), .Y(n1495) );
  NAND2X1 U1521 ( .A(n159), .B(n1557), .Y(n1487) );
  AOI22X1 U1522 ( .A(currentPlainKey[58]), .B(n1487), .C(n1557), .D(n1486), 
        .Y(n1489) );
  NAND2X1 U1523 ( .A(n1488), .B(n1561), .Y(n1524) );
  NAND2X1 U1524 ( .A(n1490), .B(n63), .Y(n1491) );
  NAND2X1 U1525 ( .A(n229), .B(n1492), .Y(n1494) );
  AOI21X1 U1526 ( .A(n1495), .B(n1494), .C(n1493), .Y(n1496) );
  MUX2X1 U1527 ( .B(n1496), .A(n260), .S(n1552), .Y(n1498) );
  NAND2X1 U1528 ( .A(n1534), .B(n254), .Y(n1497) );
  NAND2X1 U1529 ( .A(n1498), .B(n1497), .Y(n1499) );
  MUX2X1 U1530 ( .B(n1499), .A(n248), .S(n1437), .Y(n1501) );
  NAND2X1 U1531 ( .A(currentPlainKey[58]), .B(n270), .Y(n1500) );
  NAND3X1 U1532 ( .A(n1502), .B(n1501), .C(n1500), .Y(n1844) );
  NAND2X1 U1533 ( .A(n1534), .B(n278), .Y(n1518) );
  OAI22X1 U1534 ( .A(n256), .B(n7), .C(n264), .D(n63), .Y(n1514) );
  NOR2X1 U1535 ( .A(n283), .B(n1524), .Y(n1511) );
  NOR2X1 U1536 ( .A(n61), .B(n202), .Y(n1507) );
  MUX2X1 U1537 ( .B(n1700), .A(n1761), .S(n1507), .Y(n1508) );
  NAND2X1 U1538 ( .A(n1508), .B(n1524), .Y(n1509) );
  NAND2X1 U1539 ( .A(n174), .B(n1561), .Y(n1568) );
  INVX2 U1540 ( .A(n1568), .Y(n1592) );
  MUX2X1 U1541 ( .B(n1509), .A(n271), .S(n1592), .Y(n1510) );
  NOR2X1 U1542 ( .A(n1511), .B(n1510), .Y(n1512) );
  OAI22X1 U1543 ( .A(n1512), .B(n143), .C(n1589), .D(n17), .Y(n1513) );
  OAI21X1 U1544 ( .A(n1514), .B(n1513), .C(n119), .Y(n1517) );
  AOI22X1 U1545 ( .A(n1515), .B(n246), .C(currentPlainKey[59]), .D(n267), .Y(
        n1516) );
  NAND3X1 U1546 ( .A(n1518), .B(n1517), .C(n1516), .Y(n1845) );
  AOI22X1 U1547 ( .A(n1552), .B(n279), .C(currentPlainKey[60]), .D(n270), .Y(
        n1537) );
  AOI22X1 U1548 ( .A(n1592), .B(n281), .C(n1596), .D(RCV_DATA[3]), .Y(n1528)
         );
  NAND2X1 U1549 ( .A(n162), .B(n1557), .Y(n1523) );
  INVX2 U1550 ( .A(n1521), .Y(n1522) );
  AOI22X1 U1551 ( .A(currentPlainKey[60]), .B(n1523), .C(n1522), .D(n1557), 
        .Y(n1525) );
  NAND2X1 U1552 ( .A(n1568), .B(n1524), .Y(n1538) );
  NOR2X1 U1553 ( .A(n1525), .B(n1538), .Y(n1526) );
  NAND2X1 U1554 ( .A(n175), .B(n1561), .Y(n1540) );
  INVX2 U1555 ( .A(n1540), .Y(n1590) );
  MUX2X1 U1556 ( .B(n1526), .A(RCV_DATA[1]), .S(n1590), .Y(n1527) );
  NAND2X1 U1557 ( .A(n1528), .B(n1527), .Y(n1531) );
  NOR2X1 U1558 ( .A(n265), .B(n1529), .Y(n1530) );
  AOI21X1 U1559 ( .A(n1551), .B(n1531), .C(n1530), .Y(n1533) );
  NAND2X1 U1560 ( .A(n255), .B(n1571), .Y(n1532) );
  NAND2X1 U1561 ( .A(n1533), .B(n1532), .Y(n1535) );
  MUX2X1 U1562 ( .B(n1535), .A(n248), .S(n1534), .Y(n1536) );
  NAND2X1 U1563 ( .A(n1537), .B(n1536), .Y(n1846) );
  NAND2X1 U1564 ( .A(n157), .B(n1561), .Y(n1587) );
  INVX2 U1565 ( .A(n1538), .Y(n1539) );
  NAND3X1 U1566 ( .A(n1587), .B(n1540), .C(n1539), .Y(n1541) );
  INVX2 U1567 ( .A(n1541), .Y(n1565) );
  OAI21X1 U1568 ( .A(n61), .B(n206), .C(currentPlainKey[61]), .Y(n1543) );
  OAI21X1 U1569 ( .A(n61), .B(n1544), .C(n1543), .Y(n1546) );
  NOR2X1 U1570 ( .A(n271), .B(n1587), .Y(n1545) );
  AOI21X1 U1571 ( .A(n1565), .B(n1546), .C(n1545), .Y(n1549) );
  NAND2X1 U1572 ( .A(n1590), .B(n281), .Y(n1548) );
  AOI22X1 U1573 ( .A(n1592), .B(RCV_DATA[3]), .C(n1596), .D(RCV_DATA[4]), .Y(
        n1547) );
  NAND3X1 U1574 ( .A(n1549), .B(n1548), .C(n1547), .Y(n1550) );
  AOI22X1 U1575 ( .A(n115), .B(RCV_DATA[5]), .C(n1551), .D(n1550), .Y(n1555)
         );
  NAND2X1 U1576 ( .A(n280), .B(n1571), .Y(n1554) );
  AOI22X1 U1577 ( .A(n1552), .B(n246), .C(currentPlainKey[61]), .D(n267), .Y(
        n1553) );
  NAND3X1 U1578 ( .A(n1555), .B(n1554), .C(n1553), .Y(n1847) );
  AOI22X1 U1579 ( .A(n246), .B(n1571), .C(n269), .D(currentPlainKey[62]), .Y(
        n1576) );
  INVX2 U1580 ( .A(n1556), .Y(n1560) );
  AOI21X1 U1581 ( .A(n186), .B(n1557), .C(n1685), .Y(n1559) );
  NAND2X1 U1582 ( .A(n61), .B(n1685), .Y(n1558) );
  OAI21X1 U1583 ( .A(n1560), .B(n1559), .C(n1558), .Y(n1562) );
  MUX2X1 U1584 ( .B(n1562), .A(n271), .S(n170), .Y(n1564) );
  NOR2X1 U1585 ( .A(n283), .B(n1587), .Y(n1563) );
  AOI21X1 U1586 ( .A(n1565), .B(n1564), .C(n1563), .Y(n1567) );
  NAND2X1 U1587 ( .A(n1590), .B(RCV_DATA[3]), .Y(n1566) );
  NAND2X1 U1588 ( .A(n1567), .B(n1566), .Y(n1570) );
  NOR2X1 U1589 ( .A(n265), .B(n1568), .Y(n1569) );
  AOI21X1 U1590 ( .A(n227), .B(n1570), .C(n1569), .Y(n1573) );
  NAND2X1 U1591 ( .A(n1596), .B(n254), .Y(n1572) );
  AOI21X1 U1592 ( .A(n1573), .B(n1572), .C(n1571), .Y(n1574) );
  MUX2X1 U1593 ( .B(n1574), .A(n278), .S(n1598), .Y(n1575) );
  NAND2X1 U1594 ( .A(n1576), .B(n1575), .Y(n1848) );
  NAND2X1 U1595 ( .A(n266), .B(currentPlainKey[63]), .Y(n1601) );
  INVX2 U1596 ( .A(n1761), .Y(n1580) );
  NOR2X1 U1597 ( .A(n1578), .B(n204), .Y(n1579) );
  MUX2X1 U1598 ( .B(currentPlainKey[63]), .A(n1580), .S(n1579), .Y(n1585) );
  NOR2X1 U1599 ( .A(n1582), .B(n1581), .Y(n1583) );
  MUX2X1 U1600 ( .B(n1585), .A(n271), .S(n1583), .Y(n1586) );
  MUX2X1 U1601 ( .B(n1586), .A(n281), .S(n170), .Y(n1588) );
  MUX2X1 U1602 ( .B(n1589), .A(n1588), .S(n1587), .Y(n1591) );
  MUX2X1 U1603 ( .B(n1591), .A(RCV_DATA[4]), .S(n1590), .Y(n1594) );
  INVX2 U1604 ( .A(RCV_DATA[5]), .Y(n1593) );
  MUX2X1 U1605 ( .B(n1594), .A(n1593), .S(n1592), .Y(n1595) );
  NAND2X1 U1606 ( .A(n229), .B(n1595), .Y(n1597) );
  MUX2X1 U1607 ( .B(n1597), .A(n276), .S(n1596), .Y(n1599) );
  MUX2X1 U1608 ( .B(n1599), .A(n247), .S(n1598), .Y(n1600) );
  NAND2X1 U1609 ( .A(n1601), .B(n1600), .Y(n1849) );
  NAND2X1 U1610 ( .A(n1669), .B(n1602), .Y(n1614) );
  INVX2 U1611 ( .A(n1614), .Y(n1603) );
  NAND3X1 U1612 ( .A(n1603), .B(n292), .C(n1663), .Y(n1612) );
  NAND2X1 U1613 ( .A(n160), .B(n166), .Y(n1604) );
  NAND2X1 U1614 ( .A(n1613), .B(n1604), .Y(n1785) );
  NAND2X1 U1615 ( .A(n151), .B(n166), .Y(n1605) );
  NAND2X1 U1616 ( .A(n1613), .B(n1605), .Y(n1784) );
  NAND2X1 U1617 ( .A(n105), .B(n166), .Y(n1606) );
  NAND2X1 U1618 ( .A(n1613), .B(n1606), .Y(n1783) );
  MUX2X1 U1619 ( .B(n222), .A(keyCount[0]), .S(n1609), .Y(n1607) );
  NAND2X1 U1620 ( .A(n1613), .B(n1607), .Y(n1782) );
  MUX2X1 U1621 ( .B(address[4]), .A(keyCount[1]), .S(n1609), .Y(n1608) );
  NAND2X1 U1622 ( .A(n1613), .B(n1608), .Y(n1781) );
  MUX2X1 U1623 ( .B(address[5]), .A(keyCount[2]), .S(n1609), .Y(n1610) );
  NAND2X1 U1624 ( .A(n1613), .B(n1610), .Y(n1780) );
  OAI21X1 U1625 ( .A(n1696), .B(n1611), .C(n1613), .Y(n1779) );
  OAI21X1 U1626 ( .A(n1695), .B(n1611), .C(n1613), .Y(n1778) );
  OAI21X1 U1627 ( .A(n1615), .B(n1614), .C(parityError), .Y(n1618) );
  INVX2 U1628 ( .A(n1663), .Y(n1616) );
  OAI21X1 U1629 ( .A(n1988), .B(n1987), .C(n1616), .Y(n1617) );
  NAND2X1 U1630 ( .A(n1618), .B(n1617), .Y(nextParityError) );
  OAI21X1 U1631 ( .A(keyCount[0]), .B(n198), .C(n1683), .Y(n1619) );
  INVX2 U1632 ( .A(n1619), .Y(n1671) );
  NAND2X1 U1633 ( .A(n1660), .B(n1683), .Y(n1684) );
  INVX2 U1634 ( .A(n1684), .Y(n1674) );
  NAND2X1 U1635 ( .A(keyCount[0]), .B(n1674), .Y(n1679) );
  MUX2X1 U1636 ( .B(n1671), .A(n1679), .S(n1694), .Y(n1768) );
  NAND3X1 U1637 ( .A(n1661), .B(n23), .C(n1663), .Y(n1622) );
  NAND3X1 U1638 ( .A(n1620), .B(n292), .C(n1657), .Y(n1621) );
  OR2X2 U1639 ( .A(n1622), .B(n1621), .Y(n1635) );
  NAND2X1 U1640 ( .A(n1638), .B(CLR_RBUFF), .Y(n1637) );
  INVX2 U1641 ( .A(n1637), .Y(n1633) );
  NAND2X1 U1642 ( .A(N1799), .B(n1633), .Y(n1624) );
  NAND2X1 U1643 ( .A(parityAccumulator[7]), .B(n1635), .Y(n1623) );
  NAND2X1 U1644 ( .A(n1624), .B(n1623), .Y(n1777) );
  NAND2X1 U1645 ( .A(N1798), .B(n1633), .Y(n1626) );
  NAND2X1 U1646 ( .A(parityAccumulator[6]), .B(n1635), .Y(n1625) );
  NAND2X1 U1647 ( .A(n1626), .B(n1625), .Y(n1776) );
  NAND2X1 U1648 ( .A(N1797), .B(n1633), .Y(n1628) );
  NAND2X1 U1649 ( .A(n1635), .B(parityAccumulator[5]), .Y(n1627) );
  NAND2X1 U1650 ( .A(n1628), .B(n1627), .Y(n1775) );
  NAND2X1 U1651 ( .A(N1796), .B(n1633), .Y(n1630) );
  NAND2X1 U1652 ( .A(n1635), .B(parityAccumulator[4]), .Y(n1629) );
  NAND2X1 U1653 ( .A(n1630), .B(n1629), .Y(n1774) );
  NAND2X1 U1654 ( .A(N1795), .B(n1633), .Y(n1631) );
  OAI21X1 U1655 ( .A(n1691), .B(n1638), .C(n1631), .Y(n1773) );
  NAND2X1 U1656 ( .A(N1794), .B(n1633), .Y(n1632) );
  OAI21X1 U1657 ( .A(n1690), .B(n1638), .C(n1632), .Y(n1772) );
  NAND2X1 U1658 ( .A(N1793), .B(n1633), .Y(n1634) );
  OAI21X1 U1659 ( .A(n1689), .B(n1638), .C(n1634), .Y(n1771) );
  INVX2 U1660 ( .A(n1635), .Y(n1638) );
  INVX2 U1661 ( .A(N1792), .Y(n1636) );
  OAI22X1 U1662 ( .A(n1688), .B(n1638), .C(n1637), .D(n1636), .Y(n1770) );
  AOI21X1 U1663 ( .A(n1644), .B(RBUF_FULL), .C(n1920), .Y(n1639) );
  NAND2X1 U1664 ( .A(n1639), .B(n1651), .Y(n1640) );
  OAI21X1 U1665 ( .A(n224), .B(n193), .C(n1662), .Y(n1645) );
  NAND2X1 U1666 ( .A(n1640), .B(n1645), .Y(n1655) );
  NAND2X1 U1667 ( .A(n224), .B(n1655), .Y(n1641) );
  NAND2X1 U1668 ( .A(n1642), .B(n1641), .Y(n1764) );
  INVX2 U1669 ( .A(keyCount[3]), .Y(n1644) );
  AND2X2 U1670 ( .A(keyCount[2]), .B(keyCount[0]), .Y(n1643) );
  NAND3X1 U1671 ( .A(keyCount[1]), .B(n1644), .C(n1643), .Y(n1659) );
  INVX2 U1672 ( .A(n1659), .Y(n1675) );
  INVX2 U1673 ( .A(n1645), .Y(n1658) );
  AOI22X1 U1674 ( .A(n1675), .B(n1660), .C(n1658), .D(n225), .Y(n1654) );
  INVX2 U1675 ( .A(RBUF_FULL), .Y(n1646) );
  NAND2X1 U1676 ( .A(n1647), .B(n1646), .Y(n1653) );
  INVX2 U1677 ( .A(OE), .Y(n1648) );
  NAND2X1 U1678 ( .A(n1760), .B(n1648), .Y(n1650) );
  NAND2X1 U1679 ( .A(n1661), .B(n1663), .Y(n1649) );
  AOI21X1 U1680 ( .A(n1651), .B(n1650), .C(n1649), .Y(n1652) );
  NAND3X1 U1681 ( .A(n1654), .B(n1653), .C(n1652), .Y(n1766) );
  AOI21X1 U1682 ( .A(n226), .B(n1655), .C(n1660), .Y(n1656) );
  NAND3X1 U1683 ( .A(n1661), .B(n1657), .C(n1656), .Y(n1767) );
  AOI22X1 U1684 ( .A(n1660), .B(n1659), .C(n1658), .D(n164), .Y(n1670) );
  NAND2X1 U1685 ( .A(n1662), .B(n1661), .Y(n1667) );
  NAND2X1 U1686 ( .A(n1760), .B(n1648), .Y(n1665) );
  OAI21X1 U1687 ( .A(n1665), .B(n23), .C(n1663), .Y(n1666) );
  AOI21X1 U1688 ( .A(RBUF_FULL), .B(n1667), .C(n1666), .Y(n1668) );
  NAND3X1 U1689 ( .A(n1670), .B(n1669), .C(n1668), .Y(n1765) );
  NOR2X1 U1690 ( .A(keyCount[2]), .B(n198), .Y(n1673) );
  OAI21X1 U1691 ( .A(keyCount[1]), .B(n198), .C(n1671), .Y(n1678) );
  OAI21X1 U1692 ( .A(n1673), .B(n1678), .C(keyCount[3]), .Y(n1677) );
  NAND2X1 U1693 ( .A(n1675), .B(n1674), .Y(n1676) );
  NAND2X1 U1694 ( .A(n1677), .B(n1676), .Y(n1763) );
  INVX2 U1695 ( .A(n1678), .Y(n1682) );
  INVX2 U1696 ( .A(n1679), .Y(n1680) );
  NAND2X1 U1697 ( .A(n1680), .B(keyCount[1]), .Y(n1681) );
  MUX2X1 U1698 ( .B(n1682), .A(n1681), .S(n1686), .Y(n1769) );
  MUX2X1 U1699 ( .B(n1684), .A(n1683), .S(keyCount[0]), .Y(n1762) );
  INVX2 U1700 ( .A(keyCount[2]), .Y(n1686) );
  INVX2 U1701 ( .A(parityAccumulator[0]), .Y(n1688) );
  INVX2 U1702 ( .A(parityAccumulator[1]), .Y(n1689) );
  INVX2 U1703 ( .A(parityAccumulator[2]), .Y(n1690) );
  INVX2 U1704 ( .A(parityAccumulator[3]), .Y(n1691) );
  INVX2 U1705 ( .A(keyCount[1]), .Y(n1694) );
  INVX2 U1706 ( .A(address[7]), .Y(n1695) );
  INVX2 U1707 ( .A(currentPlainKey[61]), .Y(n1698) );
  INVX2 U1708 ( .A(currentPlainKey[60]), .Y(n1699) );
  INVX2 U1709 ( .A(currentPlainKey[59]), .Y(n1700) );
  INVX2 U1710 ( .A(currentPlainKey[58]), .Y(n1701) );
  INVX2 U1711 ( .A(currentPlainKey[57]), .Y(n1702) );
  INVX2 U1712 ( .A(currentPlainKey[56]), .Y(n1703) );
  INVX2 U1713 ( .A(currentPlainKey[55]), .Y(n1704) );
  INVX2 U1714 ( .A(currentPlainKey[54]), .Y(n1705) );
  INVX2 U1715 ( .A(currentPlainKey[53]), .Y(n1706) );
  INVX2 U1716 ( .A(currentPlainKey[52]), .Y(n1707) );
  INVX2 U1717 ( .A(currentPlainKey[51]), .Y(n1708) );
  INVX2 U1718 ( .A(currentPlainKey[50]), .Y(n1709) );
  INVX2 U1719 ( .A(currentPlainKey[49]), .Y(n1710) );
  INVX2 U1720 ( .A(currentPlainKey[48]), .Y(n1711) );
  INVX2 U1721 ( .A(currentPlainKey[47]), .Y(n1712) );
  INVX2 U1722 ( .A(currentPlainKey[46]), .Y(n1713) );
  INVX2 U1723 ( .A(currentPlainKey[45]), .Y(n1714) );
  INVX2 U1724 ( .A(currentPlainKey[44]), .Y(n1715) );
  INVX2 U1725 ( .A(currentPlainKey[43]), .Y(n1716) );
  INVX2 U1726 ( .A(currentPlainKey[42]), .Y(n1717) );
  INVX2 U1727 ( .A(currentPlainKey[41]), .Y(n1718) );
  INVX2 U1728 ( .A(currentPlainKey[40]), .Y(n1719) );
  INVX2 U1729 ( .A(currentPlainKey[39]), .Y(n1720) );
  INVX2 U1730 ( .A(currentPlainKey[38]), .Y(n1721) );
  INVX2 U1731 ( .A(currentPlainKey[37]), .Y(n1722) );
  INVX2 U1732 ( .A(currentPlainKey[36]), .Y(n1723) );
  INVX2 U1733 ( .A(currentPlainKey[35]), .Y(n1724) );
  INVX2 U1734 ( .A(currentPlainKey[34]), .Y(n1725) );
  INVX2 U1735 ( .A(currentPlainKey[33]), .Y(n1726) );
  INVX2 U1736 ( .A(currentPlainKey[32]), .Y(n1727) );
  INVX2 U1737 ( .A(currentPlainKey[31]), .Y(n1728) );
  INVX2 U1738 ( .A(currentPlainKey[30]), .Y(n1729) );
  INVX2 U1739 ( .A(currentPlainKey[29]), .Y(n1730) );
  INVX2 U1740 ( .A(currentPlainKey[28]), .Y(n1731) );
  INVX2 U1741 ( .A(currentPlainKey[27]), .Y(n1732) );
  INVX2 U1742 ( .A(currentPlainKey[26]), .Y(n1733) );
  INVX2 U1743 ( .A(currentPlainKey[25]), .Y(n1734) );
  INVX2 U1744 ( .A(currentPlainKey[24]), .Y(n1735) );
  INVX2 U1745 ( .A(currentPlainKey[23]), .Y(n1736) );
  INVX2 U1746 ( .A(currentPlainKey[22]), .Y(n1737) );
  INVX2 U1747 ( .A(currentPlainKey[21]), .Y(n1738) );
  INVX2 U1748 ( .A(currentPlainKey[20]), .Y(n1739) );
  INVX2 U1749 ( .A(currentPlainKey[19]), .Y(n1740) );
  INVX2 U1750 ( .A(currentPlainKey[18]), .Y(n1741) );
  INVX2 U1751 ( .A(currentPlainKey[17]), .Y(n1742) );
  INVX2 U1752 ( .A(currentPlainKey[16]), .Y(n1743) );
  INVX2 U1753 ( .A(currentPlainKey[15]), .Y(n1744) );
  INVX2 U1754 ( .A(currentPlainKey[14]), .Y(n1745) );
  INVX2 U1755 ( .A(currentPlainKey[13]), .Y(n1746) );
  INVX2 U1756 ( .A(currentPlainKey[12]), .Y(n1747) );
  INVX2 U1757 ( .A(currentPlainKey[11]), .Y(n1748) );
  INVX2 U1758 ( .A(currentPlainKey[10]), .Y(n1749) );
  INVX2 U1759 ( .A(currentPlainKey[9]), .Y(n1750) );
  INVX2 U1760 ( .A(currentPlainKey[8]), .Y(n1751) );
  INVX2 U1761 ( .A(currentPlainKey[7]), .Y(n1752) );
  INVX2 U1762 ( .A(currentPlainKey[6]), .Y(n1753) );
  INVX2 U1763 ( .A(currentPlainKey[5]), .Y(n1754) );
  INVX2 U1764 ( .A(currentPlainKey[4]), .Y(n1755) );
  INVX2 U1765 ( .A(SBE), .Y(n1760) );
  INVX2 U1766 ( .A(n220), .Y(n1761) );
endmodule


module uart_timer_0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module uart_timer_0 ( CLK, RST, TIMER_TRIG, STOP_RCVING, SHIFT_STROBE );
  input CLK, RST, TIMER_TRIG;
  output STOP_RCVING, SHIFT_STROBE;
  wire   N26, N27, N28, N29, N30, N31, N32, N33, N60, n17, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110;
  wire   [7:0] state;
  wire   [7:0] nextState;
  assign SHIFT_STROBE = N60;

  DFFSR \nextState_reg[0]  ( .D(n74), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[0]) );
  DFFSR \nextState_reg[1]  ( .D(n75), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[1]) );
  DFFSR \nextState_reg[2]  ( .D(n76), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[2]) );
  DFFSR \nextState_reg[3]  ( .D(n77), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[3]) );
  DFFSR \nextState_reg[4]  ( .D(n78), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[4]) );
  DFFSR \nextState_reg[5]  ( .D(n79), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[5]) );
  DFFSR \nextState_reg[6]  ( .D(n80), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[6]) );
  DFFSR STOP_RCVING_reg ( .D(n73), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        STOP_RCVING) );
  DFFSR \state_reg[7]  ( .D(nextState[7]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[7]) );
  DFFSR \state_reg[6]  ( .D(nextState[6]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[6]) );
  DFFSR \state_reg[5]  ( .D(nextState[5]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[5]) );
  DFFSR \state_reg[4]  ( .D(nextState[4]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[3]  ( .D(nextState[3]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        state[0]) );
  OR2X2 U21 ( .A(state[7]), .B(n95), .Y(n96) );
  OAI21X1 U38 ( .A(n20), .B(n27), .C(n110), .Y(n81) );
  NAND2X1 U39 ( .A(N33), .B(n109), .Y(n110) );
  OAI21X1 U40 ( .A(n26), .B(n20), .C(n108), .Y(n80) );
  NAND2X1 U41 ( .A(N32), .B(n109), .Y(n108) );
  OAI21X1 U42 ( .A(n25), .B(n20), .C(n107), .Y(n79) );
  NAND2X1 U43 ( .A(N31), .B(n109), .Y(n107) );
  OAI21X1 U44 ( .A(n20), .B(n24), .C(n106), .Y(n78) );
  NAND2X1 U45 ( .A(N30), .B(n109), .Y(n106) );
  OAI21X1 U46 ( .A(n23), .B(n20), .C(n105), .Y(n77) );
  NAND2X1 U47 ( .A(N29), .B(n109), .Y(n105) );
  OAI21X1 U48 ( .A(n22), .B(n20), .C(n104), .Y(n76) );
  NAND2X1 U49 ( .A(N28), .B(n109), .Y(n104) );
  OAI21X1 U50 ( .A(n20), .B(n21), .C(n103), .Y(n75) );
  NAND2X1 U51 ( .A(N27), .B(n109), .Y(n103) );
  OAI21X1 U52 ( .A(n19), .B(n20), .C(n102), .Y(n74) );
  NAND2X1 U53 ( .A(N26), .B(n109), .Y(n102) );
  NOR2X1 U54 ( .A(n101), .B(n73), .Y(n109) );
  NOR2X1 U55 ( .A(n73), .B(TIMER_TRIG), .Y(n101) );
  NOR2X1 U56 ( .A(n100), .B(n99), .Y(n73) );
  NAND3X1 U57 ( .A(nextState[6]), .B(nextState[5]), .C(n98), .Y(n99) );
  NOR2X1 U58 ( .A(n22), .B(n23), .Y(n98) );
  NAND3X1 U59 ( .A(nextState[0]), .B(n21), .C(n97), .Y(n100) );
  NOR2X1 U60 ( .A(nextState[7]), .B(nextState[4]), .Y(n97) );
  NOR2X1 U61 ( .A(state[0]), .B(n96), .Y(N60) );
  AOI21X1 U62 ( .A(n94), .B(n32), .C(n93), .Y(n95) );
  OAI21X1 U63 ( .A(n33), .B(n92), .C(n91), .Y(n93) );
  NAND3X1 U64 ( .A(state[6]), .B(state[1]), .C(n90), .Y(n91) );
  AOI21X1 U65 ( .A(n89), .B(n88), .C(state[3]), .Y(n90) );
  NAND3X1 U66 ( .A(n33), .B(n31), .C(state[4]), .Y(n88) );
  NAND3X1 U67 ( .A(state[2]), .B(n32), .C(state[5]), .Y(n89) );
  NAND2X1 U68 ( .A(state[4]), .B(n87), .Y(n92) );
  OAI21X1 U69 ( .A(state[2]), .B(n28), .C(n86), .Y(n94) );
  NAND3X1 U70 ( .A(state[2]), .B(n29), .C(n30), .Y(n86) );
  OAI22X1 U71 ( .A(state[6]), .B(n84), .C(n29), .D(n85), .Y(n87) );
  NAND3X1 U72 ( .A(n34), .B(n31), .C(state[3]), .Y(n85) );
  AOI22X1 U73 ( .A(n83), .B(state[1]), .C(n82), .D(state[5]), .Y(n84) );
  XOR2X1 U74 ( .A(n34), .B(state[3]), .Y(n82) );
  NOR2X1 U75 ( .A(state[5]), .B(state[3]), .Y(n83) );
  uart_timer_0_DW01_inc_0 add_39 ( .A(nextState), .SUM({N33, N32, N31, N30, 
        N29, N28, N27, N26}) );
  DFFSR \nextState_reg[7]  ( .D(n81), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        nextState[7]) );
  INVX2 U19 ( .A(RST), .Y(n17) );
  INVX2 U22 ( .A(nextState[0]), .Y(n19) );
  INVX2 U23 ( .A(n101), .Y(n20) );
  INVX2 U24 ( .A(nextState[1]), .Y(n21) );
  INVX2 U25 ( .A(nextState[2]), .Y(n22) );
  INVX2 U26 ( .A(nextState[3]), .Y(n23) );
  INVX2 U27 ( .A(nextState[4]), .Y(n24) );
  INVX2 U28 ( .A(nextState[5]), .Y(n25) );
  INVX2 U29 ( .A(nextState[6]), .Y(n26) );
  INVX2 U30 ( .A(nextState[7]), .Y(n27) );
  INVX2 U31 ( .A(n87), .Y(n28) );
  INVX2 U32 ( .A(state[6]), .Y(n29) );
  INVX2 U33 ( .A(n85), .Y(n30) );
  INVX2 U34 ( .A(state[5]), .Y(n31) );
  INVX2 U35 ( .A(state[4]), .Y(n32) );
  INVX2 U36 ( .A(state[2]), .Y(n33) );
  INVX2 U37 ( .A(state[1]), .Y(n34) );
endmodule


module uart_rcv_block_0 ( CLK, RST, SERIAL_IN, KEY_ERROR, PROG_ERROR, PLAINKEY, 
        RBUF_FULL, PARITY_ERROR );
  output [63:0] PLAINKEY;
  input CLK, RST, SERIAL_IN;
  output KEY_ERROR, PROG_ERROR, RBUF_FULL, PARITY_ERROR;
  wire   START_BIT, CHK_ERROR, OE, SB_DETECT, STOP_RCVING, RBUF_LOAD, SBC_CLR,
         SBC_EN, SET_RBUF_FULL, TIMER_TRIG, CLR_RBUF, SBE, SHIFT_STROBE, n1,
         n2;
  wire   [7:0] LOAD_DATA;
  wire   [7:0] RCV_DATA;
  wire   [1:0] STOP_DATA;

  uart_edge_detector_0 U_0 ( .CLK(CLK), .RST(n1), .SERIAL_IN(SERIAL_IN), 
        .START_BIT(START_BIT) );
  uart_error_0 U_1 ( .RST(n1), .CLK(CLK), .RBUF_FULL(RBUF_FULL), .CHK_ERROR(
        CHK_ERROR), .OE(OE) );
  uart_rcu_0 U_2 ( .CLK(CLK), .RST(n1), .START_BIT(START_BIT), .STOP_RCVING(
        STOP_RCVING), .SB_DETECT(SB_DETECT), .RBUF_LOAD(RBUF_LOAD), 
        .TIMER_TRIG(TIMER_TRIG), .CHK_ERROR(CHK_ERROR), .SET_RBUF_FULL(
        SET_RBUF_FULL), .SBC_EN(SBC_EN), .SBC_CLR(SBC_CLR) );
  uart_rcv_buf_0 U_3 ( .CLK(CLK), .RST(n1), .LOAD_RBUF(RBUF_LOAD), .LOAD_DATA(
        LOAD_DATA), .RCV_DATA(RCV_DATA) );
  uart_rcv_buf_full_0 U_4 ( .CLK(CLK), .RST(n1), .CLR_RBUF(CLR_RBUF), 
        .SET_RBUF_FULL(SET_RBUF_FULL), .RBUF_FULL(RBUF_FULL) );
  uart_sb_check_0 U_5 ( .RST(n1), .CLK(CLK), .SBC_CLR(SBC_CLR), .SBC_EN(SBC_EN), .STOP_DATA(STOP_DATA), .SB_DETECT(SB_DETECT), .SBE(SBE) );
  uart_sr_10bit_0 U_6 ( .CLK(CLK), .RST(n1), .SHIFT_STROBE(SHIFT_STROBE), 
        .SERIAL_IN(SERIAL_IN), .LOAD_DATA(LOAD_DATA), .STOP_DATA(STOP_DATA) );
  keyreg_0 U_8 ( .CLK(CLK), .RST(n1), .SBE(SBE), .OE(OE), .RBUF_FULL(RBUF_FULL), .RCV_DATA(RCV_DATA), .PLAINKEY(PLAINKEY), .KEY_ERROR(KEY_ERROR), 
        .PROG_ERROR(PROG_ERROR), .CLR_RBUFF(CLR_RBUF), .PARITY_ERROR(
        PARITY_ERROR) );
  uart_timer_0 U_7 ( .CLK(CLK), .RST(n1), .TIMER_TRIG(TIMER_TRIG), 
        .STOP_RCVING(STOP_RCVING), .SHIFT_STROBE(SHIFT_STROBE) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module EDBlock_0 ( BYTE, BYTE_READY, CLK, OPCODE, RST, SERIAL_IN, DATA_IN, 
        KEY_ERROR, PARITY_ERROR, PDATA_READY, PROCESSED_DATA, PROG_ERROR, 
        RBUF_FULL, W_ENABLE, R_ENABLE, DATA, ADDR );
  input [7:0] BYTE;
  input [1:0] OPCODE;
  input [7:0] DATA_IN;
  output [7:0] PROCESSED_DATA;
  output [7:0] DATA;
  output [7:0] ADDR;
  input BYTE_READY, CLK, RST, SERIAL_IN;
  output KEY_ERROR, PARITY_ERROR, PDATA_READY, PROG_ERROR, RBUF_FULL, W_ENABLE,
         R_ENABLE;

  wire   [63:0] PLAINKEY;

  KSA_0 U_0 ( .KEY(PLAINKEY), .CLK(CLK), .RST(RST), .KEY_ERROR(KEY_ERROR), 
        .BYTE_READY(BYTE_READY), .BYTE(BYTE), .OPCODE(OPCODE), .DATA_IN(
        DATA_IN), .PROCESSED_DATA(PROCESSED_DATA), .PDATA_READY(PDATA_READY), 
        .W_ENABLE(W_ENABLE), .R_ENABLE(R_ENABLE), .ADDR(ADDR), .DATA(DATA) );
  uart_rcv_block_0 U_1 ( .CLK(CLK), .RST(RST), .SERIAL_IN(SERIAL_IN), 
        .KEY_ERROR(KEY_ERROR), .PROG_ERROR(PROG_ERROR), .PLAINKEY(PLAINKEY), 
        .RBUF_FULL(RBUF_FULL), .PARITY_ERROR(PARITY_ERROR) );
endmodule


module RBUFFER_0 ( CLK, RST, NEXT_BYTE, DATA, OPCODE, BYTE_COUNT, EOP, B_READY, 
        R_ENABLE, PRGA_IN, PRGA_OPCODE );
  input [7:0] DATA;
  input [1:0] OPCODE;
  input [4:0] BYTE_COUNT;
  output [7:0] PRGA_IN;
  output [1:0] PRGA_OPCODE;
  input CLK, RST, NEXT_BYTE, EOP;
  output B_READY, R_ENABLE;
  wire   N39, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n86, n88, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103;
  wire   [2:0] state;
  wire   [2:0] nextState;
  wire   [7:0] tempData;
  wire   [1:0] tempOpcode;
  assign N39 = BYTE_COUNT[4];

  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n1), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n1), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n1), .S(1'b1), .Q(
        state[1]) );
  DFFPOSX1 B_READY_reg ( .D(n92), .CLK(CLK), .Q(B_READY) );
  DFFPOSX1 \tempData_reg[7]  ( .D(n68), .CLK(CLK), .Q(tempData[7]) );
  DFFPOSX1 \tempData_reg[6]  ( .D(n69), .CLK(CLK), .Q(tempData[6]) );
  DFFPOSX1 \tempData_reg[5]  ( .D(n70), .CLK(CLK), .Q(tempData[5]) );
  DFFPOSX1 \tempData_reg[4]  ( .D(n71), .CLK(CLK), .Q(tempData[4]) );
  DFFPOSX1 \tempData_reg[3]  ( .D(n72), .CLK(CLK), .Q(tempData[3]) );
  DFFPOSX1 \tempData_reg[2]  ( .D(n73), .CLK(CLK), .Q(tempData[2]) );
  DFFPOSX1 \tempData_reg[1]  ( .D(n74), .CLK(CLK), .Q(tempData[1]) );
  DFFPOSX1 \tempData_reg[0]  ( .D(n75), .CLK(CLK), .Q(tempData[0]) );
  DFFPOSX1 \tempOpcode_reg[1]  ( .D(n86), .CLK(CLK), .Q(tempOpcode[1]) );
  DFFPOSX1 \PRGA_OPCODE_reg[1]  ( .D(n93), .CLK(CLK), .Q(PRGA_OPCODE[1]) );
  DFFPOSX1 \tempOpcode_reg[0]  ( .D(n88), .CLK(CLK), .Q(tempOpcode[0]) );
  DFFPOSX1 \PRGA_OPCODE_reg[0]  ( .D(n94), .CLK(CLK), .Q(PRGA_OPCODE[0]) );
  DFFPOSX1 R_ENABLE_reg ( .D(n95), .CLK(CLK), .Q(R_ENABLE) );
  DFFPOSX1 \PRGA_IN_reg[7]  ( .D(n96), .CLK(CLK), .Q(PRGA_IN[7]) );
  DFFPOSX1 \PRGA_IN_reg[6]  ( .D(n97), .CLK(CLK), .Q(PRGA_IN[6]) );
  DFFPOSX1 \PRGA_IN_reg[5]  ( .D(n98), .CLK(CLK), .Q(PRGA_IN[5]) );
  DFFPOSX1 \PRGA_IN_reg[4]  ( .D(n99), .CLK(CLK), .Q(PRGA_IN[4]) );
  DFFPOSX1 \PRGA_IN_reg[3]  ( .D(n100), .CLK(CLK), .Q(PRGA_IN[3]) );
  DFFPOSX1 \PRGA_IN_reg[2]  ( .D(n101), .CLK(CLK), .Q(PRGA_IN[2]) );
  DFFPOSX1 \PRGA_IN_reg[1]  ( .D(n102), .CLK(CLK), .Q(PRGA_IN[1]) );
  DFFPOSX1 \PRGA_IN_reg[0]  ( .D(n103), .CLK(CLK), .Q(PRGA_IN[0]) );
  INVX2 U3 ( .A(n41), .Y(n28) );
  INVX2 U4 ( .A(RST), .Y(n1) );
  OR2X2 U5 ( .A(n39), .B(RST), .Y(n29) );
  AND2X2 U6 ( .A(n39), .B(n1), .Y(n44) );
  OAI21X1 U7 ( .A(n2), .B(n3), .C(n4), .Y(nextState[2]) );
  MUX2X1 U8 ( .B(n5), .A(n6), .S(state[0]), .Y(n4) );
  NOR2X1 U9 ( .A(state[2]), .B(n7), .Y(n6) );
  AND2X1 U10 ( .A(state[2]), .B(n8), .Y(n5) );
  OAI21X1 U11 ( .A(NEXT_BYTE), .B(n9), .C(state[1]), .Y(n8) );
  AND2X1 U12 ( .A(n10), .B(NEXT_BYTE), .Y(n2) );
  OAI21X1 U13 ( .A(state[2]), .B(n11), .C(n12), .Y(nextState[1]) );
  OAI21X1 U14 ( .A(n13), .B(n14), .C(n15), .Y(n12) );
  INVX1 U15 ( .A(n3), .Y(n14) );
  OAI21X1 U16 ( .A(state[2]), .B(n16), .C(n17), .Y(nextState[0]) );
  AOI22X1 U17 ( .A(n18), .B(n19), .C(NEXT_BYTE), .D(n20), .Y(n17) );
  OAI21X1 U18 ( .A(n10), .B(n3), .C(n21), .Y(n20) );
  INVX1 U19 ( .A(n13), .Y(n21) );
  NOR2X1 U20 ( .A(n16), .B(n9), .Y(n13) );
  NOR2X1 U21 ( .A(n22), .B(N39), .Y(n9) );
  NAND3X1 U22 ( .A(state[0]), .B(n7), .C(state[2]), .Y(n3) );
  AND2X1 U23 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n10) );
  OAI21X1 U24 ( .A(n23), .B(n15), .C(n24), .Y(n19) );
  INVX1 U25 ( .A(NEXT_BYTE), .Y(n15) );
  AOI21X1 U26 ( .A(EOP), .B(n22), .C(N39), .Y(n23) );
  NAND2X1 U27 ( .A(n25), .B(n26), .Y(n22) );
  NOR2X1 U28 ( .A(BYTE_COUNT[3]), .B(BYTE_COUNT[2]), .Y(n26) );
  NOR2X1 U29 ( .A(BYTE_COUNT[1]), .B(BYTE_COUNT[0]), .Y(n25) );
  NOR2X1 U30 ( .A(state[1]), .B(state[0]), .Y(n18) );
  INVX1 U31 ( .A(n27), .Y(n68) );
  AOI22X1 U32 ( .A(n28), .B(DATA[7]), .C(n29), .D(tempData[7]), .Y(n27) );
  INVX1 U33 ( .A(n30), .Y(n69) );
  AOI22X1 U34 ( .A(n28), .B(DATA[6]), .C(n29), .D(tempData[6]), .Y(n30) );
  INVX1 U35 ( .A(n31), .Y(n70) );
  AOI22X1 U36 ( .A(n28), .B(DATA[5]), .C(n29), .D(tempData[5]), .Y(n31) );
  INVX1 U37 ( .A(n32), .Y(n71) );
  AOI22X1 U38 ( .A(n28), .B(DATA[4]), .C(n29), .D(tempData[4]), .Y(n32) );
  INVX1 U39 ( .A(n33), .Y(n72) );
  AOI22X1 U40 ( .A(n28), .B(DATA[3]), .C(n29), .D(tempData[3]), .Y(n33) );
  INVX1 U41 ( .A(n34), .Y(n73) );
  AOI22X1 U42 ( .A(n28), .B(DATA[2]), .C(n29), .D(tempData[2]), .Y(n34) );
  INVX1 U43 ( .A(n35), .Y(n74) );
  AOI22X1 U44 ( .A(n28), .B(DATA[1]), .C(n29), .D(tempData[1]), .Y(n35) );
  INVX1 U45 ( .A(n36), .Y(n75) );
  AOI22X1 U46 ( .A(n28), .B(DATA[0]), .C(n29), .D(tempData[0]), .Y(n36) );
  INVX1 U47 ( .A(n37), .Y(n86) );
  AOI22X1 U48 ( .A(OPCODE[1]), .B(n28), .C(n29), .D(tempOpcode[1]), .Y(n37) );
  INVX1 U49 ( .A(n38), .Y(n88) );
  AOI22X1 U50 ( .A(OPCODE[0]), .B(n28), .C(n29), .D(tempOpcode[0]), .Y(n38) );
  OAI21X1 U51 ( .A(n1), .B(n40), .C(n41), .Y(n92) );
  INVX1 U52 ( .A(B_READY), .Y(n40) );
  OAI21X1 U53 ( .A(n1), .B(n42), .C(n43), .Y(n93) );
  AOI22X1 U54 ( .A(n28), .B(OPCODE[1]), .C(n44), .D(tempOpcode[1]), .Y(n43) );
  INVX1 U55 ( .A(PRGA_OPCODE[1]), .Y(n42) );
  OAI21X1 U56 ( .A(n1), .B(n45), .C(n46), .Y(n94) );
  AOI22X1 U57 ( .A(n28), .B(OPCODE[0]), .C(n44), .D(tempOpcode[0]), .Y(n46) );
  INVX1 U58 ( .A(PRGA_OPCODE[0]), .Y(n45) );
  MUX2X1 U59 ( .B(n47), .A(n48), .S(RST), .Y(n95) );
  INVX1 U60 ( .A(R_ENABLE), .Y(n48) );
  NAND3X1 U61 ( .A(n7), .B(n24), .C(state[0]), .Y(n47) );
  OAI21X1 U62 ( .A(n1), .B(n49), .C(n50), .Y(n96) );
  AOI22X1 U63 ( .A(DATA[7]), .B(n28), .C(n44), .D(tempData[7]), .Y(n50) );
  INVX1 U64 ( .A(PRGA_IN[7]), .Y(n49) );
  OAI21X1 U65 ( .A(n1), .B(n51), .C(n52), .Y(n97) );
  AOI22X1 U66 ( .A(DATA[6]), .B(n28), .C(n44), .D(tempData[6]), .Y(n52) );
  INVX1 U67 ( .A(PRGA_IN[6]), .Y(n51) );
  OAI21X1 U68 ( .A(n1), .B(n53), .C(n54), .Y(n98) );
  AOI22X1 U69 ( .A(DATA[5]), .B(n28), .C(n44), .D(tempData[5]), .Y(n54) );
  INVX1 U70 ( .A(PRGA_IN[5]), .Y(n53) );
  OAI21X1 U71 ( .A(n1), .B(n55), .C(n56), .Y(n99) );
  AOI22X1 U72 ( .A(DATA[4]), .B(n28), .C(n44), .D(tempData[4]), .Y(n56) );
  INVX1 U73 ( .A(PRGA_IN[4]), .Y(n55) );
  OAI21X1 U74 ( .A(n1), .B(n57), .C(n58), .Y(n100) );
  AOI22X1 U75 ( .A(DATA[3]), .B(n28), .C(n44), .D(tempData[3]), .Y(n58) );
  INVX1 U76 ( .A(PRGA_IN[3]), .Y(n57) );
  OAI21X1 U77 ( .A(n1), .B(n59), .C(n60), .Y(n101) );
  AOI22X1 U78 ( .A(DATA[2]), .B(n28), .C(n44), .D(tempData[2]), .Y(n60) );
  INVX1 U79 ( .A(PRGA_IN[2]), .Y(n59) );
  OAI21X1 U80 ( .A(n1), .B(n61), .C(n62), .Y(n102) );
  AOI22X1 U81 ( .A(DATA[1]), .B(n28), .C(n44), .D(tempData[1]), .Y(n62) );
  INVX1 U82 ( .A(PRGA_IN[1]), .Y(n61) );
  OAI21X1 U83 ( .A(n1), .B(n63), .C(n64), .Y(n103) );
  AOI22X1 U84 ( .A(DATA[0]), .B(n28), .C(n44), .D(tempData[0]), .Y(n64) );
  NAND2X1 U85 ( .A(n11), .B(state[2]), .Y(n39) );
  INVX1 U86 ( .A(n65), .Y(n11) );
  OAI21X1 U87 ( .A(state[1]), .B(n66), .C(n16), .Y(n65) );
  NAND2X1 U88 ( .A(state[1]), .B(n66), .Y(n16) );
  NAND3X1 U89 ( .A(n66), .B(n7), .C(n67), .Y(n41) );
  NOR2X1 U90 ( .A(RST), .B(n24), .Y(n67) );
  INVX1 U91 ( .A(state[2]), .Y(n24) );
  INVX1 U92 ( .A(state[1]), .Y(n7) );
  INVX1 U93 ( .A(state[0]), .Y(n66) );
  INVX1 U94 ( .A(PRGA_IN[0]), .Y(n63) );
endmodule


module RFIFO_0 ( CLK, RST, W_ENABLE, R_ENABLE, RCV_DATA, RCV_OPCODE, DATA, 
        OUT_OPCODE, BYTE_COUNT, EMPTY, FULL );
  input [7:0] RCV_DATA;
  input [1:0] RCV_OPCODE;
  output [7:0] DATA;
  output [1:0] OUT_OPCODE;
  output [4:0] BYTE_COUNT;
  input CLK, RST, W_ENABLE, R_ENABLE;
  output EMPTY, FULL;
  wire   state, \opcode[0][1] , \opcode[0][0] , \opcode[1][1] , \opcode[1][0] ,
         \opcode[2][1] , \opcode[2][0] , \opcode[3][1] , \opcode[3][0] ,
         \opcode[4][1] , \opcode[4][0] , \opcode[5][1] , \opcode[5][0] ,
         \opcode[6][1] , \opcode[6][0] , \opcode[7][1] , \opcode[7][0] ,
         \opcode[8][1] , \opcode[8][0] , \opcode[9][1] , \opcode[9][0] ,
         \opcode[10][1] , \opcode[10][0] , \opcode[11][1] , \opcode[11][0] ,
         \opcode[12][1] , \opcode[12][0] , \opcode[13][1] , \opcode[13][0] ,
         \opcode[14][1] , \opcode[14][0] , \opcode[15][1] , \opcode[15][0] ,
         \opcode[16][1] , \opcode[16][0] , \opcode[17][1] , \opcode[17][0] ,
         \opcode[18][1] , \opcode[18][0] , \opcode[19][1] , \opcode[19][0] ,
         \opcode[20][1] , \opcode[20][0] , \opcode[21][1] , \opcode[21][0] ,
         \opcode[22][1] , \opcode[22][0] , \opcode[23][1] , \opcode[23][0] ,
         \opcode[24][1] , \opcode[24][0] , \opcode[25][1] , \opcode[25][0] ,
         \opcode[26][1] , \opcode[26][0] , \opcode[27][1] , \opcode[27][0] ,
         \opcode[28][1] , \opcode[28][0] , \opcode[29][1] , \opcode[29][0] ,
         \opcode[30][1] , \opcode[30][0] , \opcode[31][1] , \opcode[31][0] ,
         \memory[0][7] , \memory[0][6] , \memory[0][5] , \memory[0][4] ,
         \memory[0][3] , \memory[0][2] , \memory[0][1] , \memory[0][0] ,
         \memory[1][7] , \memory[1][6] , \memory[1][5] , \memory[1][4] ,
         \memory[1][3] , \memory[1][2] , \memory[1][1] , \memory[1][0] ,
         \memory[2][7] , \memory[2][6] , \memory[2][5] , \memory[2][4] ,
         \memory[2][3] , \memory[2][2] , \memory[2][1] , \memory[2][0] ,
         \memory[3][7] , \memory[3][6] , \memory[3][5] , \memory[3][4] ,
         \memory[3][3] , \memory[3][2] , \memory[3][1] , \memory[3][0] ,
         \memory[4][7] , \memory[4][6] , \memory[4][5] , \memory[4][4] ,
         \memory[4][3] , \memory[4][2] , \memory[4][1] , \memory[4][0] ,
         \memory[5][7] , \memory[5][6] , \memory[5][5] , \memory[5][4] ,
         \memory[5][3] , \memory[5][2] , \memory[5][1] , \memory[5][0] ,
         \memory[6][7] , \memory[6][6] , \memory[6][5] , \memory[6][4] ,
         \memory[6][3] , \memory[6][2] , \memory[6][1] , \memory[6][0] ,
         \memory[7][7] , \memory[7][6] , \memory[7][5] , \memory[7][4] ,
         \memory[7][3] , \memory[7][2] , \memory[7][1] , \memory[7][0] ,
         \memory[8][7] , \memory[8][6] , \memory[8][5] , \memory[8][4] ,
         \memory[8][3] , \memory[8][2] , \memory[8][1] , \memory[8][0] ,
         \memory[9][7] , \memory[9][6] , \memory[9][5] , \memory[9][4] ,
         \memory[9][3] , \memory[9][2] , \memory[9][1] , \memory[9][0] ,
         \memory[10][7] , \memory[10][6] , \memory[10][5] , \memory[10][4] ,
         \memory[10][3] , \memory[10][2] , \memory[10][1] , \memory[10][0] ,
         \memory[11][7] , \memory[11][6] , \memory[11][5] , \memory[11][4] ,
         \memory[11][3] , \memory[11][2] , \memory[11][1] , \memory[11][0] ,
         \memory[12][7] , \memory[12][6] , \memory[12][5] , \memory[12][4] ,
         \memory[12][3] , \memory[12][2] , \memory[12][1] , \memory[12][0] ,
         \memory[13][7] , \memory[13][6] , \memory[13][5] , \memory[13][4] ,
         \memory[13][3] , \memory[13][2] , \memory[13][1] , \memory[13][0] ,
         \memory[14][7] , \memory[14][6] , \memory[14][5] , \memory[14][4] ,
         \memory[14][3] , \memory[14][2] , \memory[14][1] , \memory[14][0] ,
         \memory[15][7] , \memory[15][6] , \memory[15][5] , \memory[15][4] ,
         \memory[15][3] , \memory[15][2] , \memory[15][1] , \memory[15][0] ,
         \memory[16][7] , \memory[16][6] , \memory[16][5] , \memory[16][4] ,
         \memory[16][3] , \memory[16][2] , \memory[16][1] , \memory[16][0] ,
         \memory[17][7] , \memory[17][6] , \memory[17][5] , \memory[17][4] ,
         \memory[17][3] , \memory[17][2] , \memory[17][1] , \memory[17][0] ,
         \memory[18][7] , \memory[18][6] , \memory[18][5] , \memory[18][4] ,
         \memory[18][3] , \memory[18][2] , \memory[18][1] , \memory[18][0] ,
         \memory[19][7] , \memory[19][6] , \memory[19][5] , \memory[19][4] ,
         \memory[19][3] , \memory[19][2] , \memory[19][1] , \memory[19][0] ,
         \memory[20][7] , \memory[20][6] , \memory[20][5] , \memory[20][4] ,
         \memory[20][3] , \memory[20][2] , \memory[20][1] , \memory[20][0] ,
         \memory[21][7] , \memory[21][6] , \memory[21][5] , \memory[21][4] ,
         \memory[21][3] , \memory[21][2] , \memory[21][1] , \memory[21][0] ,
         \memory[22][7] , \memory[22][6] , \memory[22][5] , \memory[22][4] ,
         \memory[22][3] , \memory[22][2] , \memory[22][1] , \memory[22][0] ,
         \memory[23][7] , \memory[23][6] , \memory[23][5] , \memory[23][4] ,
         \memory[23][3] , \memory[23][2] , \memory[23][1] , \memory[23][0] ,
         \memory[24][7] , \memory[24][6] , \memory[24][5] , \memory[24][4] ,
         \memory[24][3] , \memory[24][2] , \memory[24][1] , \memory[24][0] ,
         \memory[25][7] , \memory[25][6] , \memory[25][5] , \memory[25][4] ,
         \memory[25][3] , \memory[25][2] , \memory[25][1] , \memory[25][0] ,
         \memory[26][7] , \memory[26][6] , \memory[26][5] , \memory[26][4] ,
         \memory[26][3] , \memory[26][2] , \memory[26][1] , \memory[26][0] ,
         \memory[27][7] , \memory[27][6] , \memory[27][5] , \memory[27][4] ,
         \memory[27][3] , \memory[27][2] , \memory[27][1] , \memory[27][0] ,
         \memory[28][7] , \memory[28][6] , \memory[28][5] , \memory[28][4] ,
         \memory[28][3] , \memory[28][2] , \memory[28][1] , \memory[28][0] ,
         \memory[29][7] , \memory[29][6] , \memory[29][5] , \memory[29][4] ,
         \memory[29][3] , \memory[29][2] , \memory[29][1] , \memory[29][0] ,
         \memory[30][7] , \memory[30][6] , \memory[30][5] , \memory[30][4] ,
         \memory[30][3] , \memory[30][2] , \memory[30][1] , \memory[30][0] ,
         \memory[31][7] , \memory[31][6] , \memory[31][5] , \memory[31][4] ,
         \memory[31][3] , \memory[31][2] , \memory[31][1] , \memory[31][0] ,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n852, n861, n863, n865, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1607, n1608, n1610, n1612, n1614;
  wire   [4:0] readptr;
  wire   [4:0] writeptr;

  DFFSR state_reg ( .D(1'b1), .CLK(CLK), .R(n163), .S(1'b1), .Q(state) );
  DFFSR \readptr_reg[0]  ( .D(N343), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        readptr[0]) );
  DFFSR \readptr_reg[1]  ( .D(N344), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        readptr[1]) );
  DFFSR \readptr_reg[3]  ( .D(N346), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        readptr[3]) );
  DFFSR \writeptr_reg[3]  ( .D(n1608), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        writeptr[3]) );
  DFFSR \writeptr_reg[0]  ( .D(n1610), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        writeptr[0]) );
  DFFSR \writeptr_reg[1]  ( .D(n1612), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        writeptr[1]) );
  DFFSR \writeptr_reg[2]  ( .D(n1614), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        writeptr[2]) );
  DFFPOSX1 FULL_reg ( .D(n1431), .CLK(CLK), .Q(FULL) );
  DFFSR \BYTE_COUNT_reg[4]  ( .D(N342), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        BYTE_COUNT[4]) );
  DFFSR \BYTE_COUNT_reg[3]  ( .D(N341), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        BYTE_COUNT[3]) );
  DFFSR \BYTE_COUNT_reg[2]  ( .D(N340), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        BYTE_COUNT[2]) );
  DFFSR \BYTE_COUNT_reg[1]  ( .D(N339), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        BYTE_COUNT[1]) );
  DFFSR \BYTE_COUNT_reg[0]  ( .D(N338), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        BYTE_COUNT[0]) );
  DFFPOSX1 \memory_reg[0][7]  ( .D(n1406), .CLK(CLK), .Q(\memory[0][7] ) );
  DFFPOSX1 \memory_reg[0][6]  ( .D(n1405), .CLK(CLK), .Q(\memory[0][6] ) );
  DFFPOSX1 \memory_reg[0][5]  ( .D(n1404), .CLK(CLK), .Q(\memory[0][5] ) );
  DFFPOSX1 \memory_reg[0][4]  ( .D(n1403), .CLK(CLK), .Q(\memory[0][4] ) );
  DFFPOSX1 \memory_reg[0][3]  ( .D(n1402), .CLK(CLK), .Q(\memory[0][3] ) );
  DFFPOSX1 \memory_reg[0][2]  ( .D(n1401), .CLK(CLK), .Q(\memory[0][2] ) );
  DFFPOSX1 \memory_reg[0][1]  ( .D(n1400), .CLK(CLK), .Q(\memory[0][1] ) );
  DFFPOSX1 \memory_reg[0][0]  ( .D(n1399), .CLK(CLK), .Q(\memory[0][0] ) );
  DFFPOSX1 \memory_reg[1][7]  ( .D(n1414), .CLK(CLK), .Q(\memory[1][7] ) );
  DFFPOSX1 \memory_reg[1][6]  ( .D(n1413), .CLK(CLK), .Q(\memory[1][6] ) );
  DFFPOSX1 \memory_reg[1][5]  ( .D(n1412), .CLK(CLK), .Q(\memory[1][5] ) );
  DFFPOSX1 \memory_reg[1][4]  ( .D(n1411), .CLK(CLK), .Q(\memory[1][4] ) );
  DFFPOSX1 \memory_reg[1][3]  ( .D(n1410), .CLK(CLK), .Q(\memory[1][3] ) );
  DFFPOSX1 \memory_reg[1][2]  ( .D(n1409), .CLK(CLK), .Q(\memory[1][2] ) );
  DFFPOSX1 \memory_reg[1][1]  ( .D(n1408), .CLK(CLK), .Q(\memory[1][1] ) );
  DFFPOSX1 \memory_reg[1][0]  ( .D(n1407), .CLK(CLK), .Q(\memory[1][0] ) );
  DFFPOSX1 \memory_reg[2][7]  ( .D(n1422), .CLK(CLK), .Q(\memory[2][7] ) );
  DFFPOSX1 \memory_reg[2][6]  ( .D(n1421), .CLK(CLK), .Q(\memory[2][6] ) );
  DFFPOSX1 \memory_reg[2][5]  ( .D(n1420), .CLK(CLK), .Q(\memory[2][5] ) );
  DFFPOSX1 \memory_reg[2][4]  ( .D(n1419), .CLK(CLK), .Q(\memory[2][4] ) );
  DFFPOSX1 \memory_reg[2][3]  ( .D(n1418), .CLK(CLK), .Q(\memory[2][3] ) );
  DFFPOSX1 \memory_reg[2][2]  ( .D(n1417), .CLK(CLK), .Q(\memory[2][2] ) );
  DFFPOSX1 \memory_reg[2][1]  ( .D(n1416), .CLK(CLK), .Q(\memory[2][1] ) );
  DFFPOSX1 \memory_reg[2][0]  ( .D(n1415), .CLK(CLK), .Q(\memory[2][0] ) );
  DFFPOSX1 \memory_reg[3][7]  ( .D(n1430), .CLK(CLK), .Q(\memory[3][7] ) );
  DFFPOSX1 \memory_reg[3][6]  ( .D(n1429), .CLK(CLK), .Q(\memory[3][6] ) );
  DFFPOSX1 \memory_reg[3][5]  ( .D(n1428), .CLK(CLK), .Q(\memory[3][5] ) );
  DFFPOSX1 \memory_reg[3][4]  ( .D(n1427), .CLK(CLK), .Q(\memory[3][4] ) );
  DFFPOSX1 \memory_reg[3][3]  ( .D(n1426), .CLK(CLK), .Q(\memory[3][3] ) );
  DFFPOSX1 \memory_reg[3][2]  ( .D(n1425), .CLK(CLK), .Q(\memory[3][2] ) );
  DFFPOSX1 \memory_reg[3][1]  ( .D(n1424), .CLK(CLK), .Q(\memory[3][1] ) );
  DFFPOSX1 \memory_reg[3][0]  ( .D(n1423), .CLK(CLK), .Q(\memory[3][0] ) );
  DFFPOSX1 \memory_reg[4][7]  ( .D(n1602), .CLK(CLK), .Q(\memory[4][7] ) );
  DFFPOSX1 \memory_reg[4][6]  ( .D(n1601), .CLK(CLK), .Q(\memory[4][6] ) );
  DFFPOSX1 \memory_reg[4][5]  ( .D(n1600), .CLK(CLK), .Q(\memory[4][5] ) );
  DFFPOSX1 \memory_reg[4][4]  ( .D(n1599), .CLK(CLK), .Q(\memory[4][4] ) );
  DFFPOSX1 \memory_reg[4][3]  ( .D(n1598), .CLK(CLK), .Q(\memory[4][3] ) );
  DFFPOSX1 \memory_reg[4][2]  ( .D(n1597), .CLK(CLK), .Q(\memory[4][2] ) );
  DFFPOSX1 \memory_reg[4][1]  ( .D(n1596), .CLK(CLK), .Q(\memory[4][1] ) );
  DFFPOSX1 \memory_reg[4][0]  ( .D(n1595), .CLK(CLK), .Q(\memory[4][0] ) );
  DFFPOSX1 \memory_reg[5][7]  ( .D(n1592), .CLK(CLK), .Q(\memory[5][7] ) );
  DFFPOSX1 \memory_reg[5][6]  ( .D(n1591), .CLK(CLK), .Q(\memory[5][6] ) );
  DFFPOSX1 \memory_reg[5][5]  ( .D(n1590), .CLK(CLK), .Q(\memory[5][5] ) );
  DFFPOSX1 \memory_reg[5][4]  ( .D(n1589), .CLK(CLK), .Q(\memory[5][4] ) );
  DFFPOSX1 \memory_reg[5][3]  ( .D(n1588), .CLK(CLK), .Q(\memory[5][3] ) );
  DFFPOSX1 \memory_reg[5][2]  ( .D(n1587), .CLK(CLK), .Q(\memory[5][2] ) );
  DFFPOSX1 \memory_reg[5][1]  ( .D(n1586), .CLK(CLK), .Q(\memory[5][1] ) );
  DFFPOSX1 \memory_reg[5][0]  ( .D(n1585), .CLK(CLK), .Q(\memory[5][0] ) );
  DFFPOSX1 \memory_reg[6][7]  ( .D(n1582), .CLK(CLK), .Q(\memory[6][7] ) );
  DFFPOSX1 \memory_reg[6][6]  ( .D(n1581), .CLK(CLK), .Q(\memory[6][6] ) );
  DFFPOSX1 \memory_reg[6][5]  ( .D(n1580), .CLK(CLK), .Q(\memory[6][5] ) );
  DFFPOSX1 \memory_reg[6][4]  ( .D(n1579), .CLK(CLK), .Q(\memory[6][4] ) );
  DFFPOSX1 \memory_reg[6][3]  ( .D(n1578), .CLK(CLK), .Q(\memory[6][3] ) );
  DFFPOSX1 \memory_reg[6][2]  ( .D(n1577), .CLK(CLK), .Q(\memory[6][2] ) );
  DFFPOSX1 \memory_reg[6][1]  ( .D(n1576), .CLK(CLK), .Q(\memory[6][1] ) );
  DFFPOSX1 \memory_reg[6][0]  ( .D(n1575), .CLK(CLK), .Q(\memory[6][0] ) );
  DFFPOSX1 \memory_reg[7][7]  ( .D(n1572), .CLK(CLK), .Q(\memory[7][7] ) );
  DFFPOSX1 \memory_reg[7][6]  ( .D(n1571), .CLK(CLK), .Q(\memory[7][6] ) );
  DFFPOSX1 \memory_reg[7][5]  ( .D(n1570), .CLK(CLK), .Q(\memory[7][5] ) );
  DFFPOSX1 \memory_reg[7][4]  ( .D(n1569), .CLK(CLK), .Q(\memory[7][4] ) );
  DFFPOSX1 \memory_reg[7][3]  ( .D(n1568), .CLK(CLK), .Q(\memory[7][3] ) );
  DFFPOSX1 \memory_reg[7][2]  ( .D(n1567), .CLK(CLK), .Q(\memory[7][2] ) );
  DFFPOSX1 \memory_reg[7][1]  ( .D(n1566), .CLK(CLK), .Q(\memory[7][1] ) );
  DFFPOSX1 \memory_reg[7][0]  ( .D(n1565), .CLK(CLK), .Q(\memory[7][0] ) );
  DFFPOSX1 \memory_reg[8][7]  ( .D(n1433), .CLK(CLK), .Q(\memory[8][7] ) );
  DFFPOSX1 \memory_reg[8][6]  ( .D(n1434), .CLK(CLK), .Q(\memory[8][6] ) );
  DFFPOSX1 \memory_reg[8][5]  ( .D(n1435), .CLK(CLK), .Q(\memory[8][5] ) );
  DFFPOSX1 \memory_reg[8][4]  ( .D(n1436), .CLK(CLK), .Q(\memory[8][4] ) );
  DFFPOSX1 \memory_reg[8][3]  ( .D(n1437), .CLK(CLK), .Q(\memory[8][3] ) );
  DFFPOSX1 \memory_reg[8][2]  ( .D(n1438), .CLK(CLK), .Q(\memory[8][2] ) );
  DFFPOSX1 \memory_reg[8][1]  ( .D(n1439), .CLK(CLK), .Q(\memory[8][1] ) );
  DFFPOSX1 \memory_reg[8][0]  ( .D(n1440), .CLK(CLK), .Q(\memory[8][0] ) );
  DFFPOSX1 \memory_reg[9][7]  ( .D(n1441), .CLK(CLK), .Q(\memory[9][7] ) );
  DFFPOSX1 \memory_reg[9][6]  ( .D(n1442), .CLK(CLK), .Q(\memory[9][6] ) );
  DFFPOSX1 \memory_reg[9][5]  ( .D(n1443), .CLK(CLK), .Q(\memory[9][5] ) );
  DFFPOSX1 \memory_reg[9][4]  ( .D(n1444), .CLK(CLK), .Q(\memory[9][4] ) );
  DFFPOSX1 \memory_reg[9][3]  ( .D(n1445), .CLK(CLK), .Q(\memory[9][3] ) );
  DFFPOSX1 \memory_reg[9][2]  ( .D(n1446), .CLK(CLK), .Q(\memory[9][2] ) );
  DFFPOSX1 \memory_reg[9][1]  ( .D(n1447), .CLK(CLK), .Q(\memory[9][1] ) );
  DFFPOSX1 \memory_reg[9][0]  ( .D(n1448), .CLK(CLK), .Q(\memory[9][0] ) );
  DFFPOSX1 \memory_reg[10][7]  ( .D(n1449), .CLK(CLK), .Q(\memory[10][7] ) );
  DFFPOSX1 \memory_reg[10][6]  ( .D(n1450), .CLK(CLK), .Q(\memory[10][6] ) );
  DFFPOSX1 \memory_reg[10][5]  ( .D(n1451), .CLK(CLK), .Q(\memory[10][5] ) );
  DFFPOSX1 \memory_reg[10][4]  ( .D(n1452), .CLK(CLK), .Q(\memory[10][4] ) );
  DFFPOSX1 \memory_reg[10][3]  ( .D(n1453), .CLK(CLK), .Q(\memory[10][3] ) );
  DFFPOSX1 \memory_reg[10][2]  ( .D(n1454), .CLK(CLK), .Q(\memory[10][2] ) );
  DFFPOSX1 \memory_reg[10][1]  ( .D(n1455), .CLK(CLK), .Q(\memory[10][1] ) );
  DFFPOSX1 \memory_reg[10][0]  ( .D(n1456), .CLK(CLK), .Q(\memory[10][0] ) );
  DFFPOSX1 \memory_reg[11][7]  ( .D(n1457), .CLK(CLK), .Q(\memory[11][7] ) );
  DFFPOSX1 \memory_reg[11][6]  ( .D(n1458), .CLK(CLK), .Q(\memory[11][6] ) );
  DFFPOSX1 \memory_reg[11][5]  ( .D(n1459), .CLK(CLK), .Q(\memory[11][5] ) );
  DFFPOSX1 \memory_reg[11][4]  ( .D(n1460), .CLK(CLK), .Q(\memory[11][4] ) );
  DFFPOSX1 \memory_reg[11][3]  ( .D(n1461), .CLK(CLK), .Q(\memory[11][3] ) );
  DFFPOSX1 \memory_reg[11][2]  ( .D(n1462), .CLK(CLK), .Q(\memory[11][2] ) );
  DFFPOSX1 \memory_reg[11][1]  ( .D(n1463), .CLK(CLK), .Q(\memory[11][1] ) );
  DFFPOSX1 \memory_reg[11][0]  ( .D(n1464), .CLK(CLK), .Q(\memory[11][0] ) );
  DFFPOSX1 \memory_reg[12][7]  ( .D(n1391), .CLK(CLK), .Q(\memory[12][7] ) );
  DFFPOSX1 \memory_reg[12][6]  ( .D(n1392), .CLK(CLK), .Q(\memory[12][6] ) );
  DFFPOSX1 \memory_reg[12][5]  ( .D(n1393), .CLK(CLK), .Q(\memory[12][5] ) );
  DFFPOSX1 \memory_reg[12][4]  ( .D(n1394), .CLK(CLK), .Q(\memory[12][4] ) );
  DFFPOSX1 \memory_reg[12][3]  ( .D(n1395), .CLK(CLK), .Q(\memory[12][3] ) );
  DFFPOSX1 \memory_reg[12][2]  ( .D(n1396), .CLK(CLK), .Q(\memory[12][2] ) );
  DFFPOSX1 \memory_reg[12][1]  ( .D(n1397), .CLK(CLK), .Q(\memory[12][1] ) );
  DFFPOSX1 \memory_reg[12][0]  ( .D(n1398), .CLK(CLK), .Q(\memory[12][0] ) );
  DFFPOSX1 \memory_reg[13][7]  ( .D(n1383), .CLK(CLK), .Q(\memory[13][7] ) );
  DFFPOSX1 \memory_reg[13][6]  ( .D(n1384), .CLK(CLK), .Q(\memory[13][6] ) );
  DFFPOSX1 \memory_reg[13][5]  ( .D(n1385), .CLK(CLK), .Q(\memory[13][5] ) );
  DFFPOSX1 \memory_reg[13][4]  ( .D(n1386), .CLK(CLK), .Q(\memory[13][4] ) );
  DFFPOSX1 \memory_reg[13][3]  ( .D(n1387), .CLK(CLK), .Q(\memory[13][3] ) );
  DFFPOSX1 \memory_reg[13][2]  ( .D(n1388), .CLK(CLK), .Q(\memory[13][2] ) );
  DFFPOSX1 \memory_reg[13][1]  ( .D(n1389), .CLK(CLK), .Q(\memory[13][1] ) );
  DFFPOSX1 \memory_reg[13][0]  ( .D(n1390), .CLK(CLK), .Q(\memory[13][0] ) );
  DFFPOSX1 \memory_reg[14][7]  ( .D(n1375), .CLK(CLK), .Q(\memory[14][7] ) );
  DFFPOSX1 \memory_reg[14][6]  ( .D(n1376), .CLK(CLK), .Q(\memory[14][6] ) );
  DFFPOSX1 \memory_reg[14][5]  ( .D(n1377), .CLK(CLK), .Q(\memory[14][5] ) );
  DFFPOSX1 \memory_reg[14][4]  ( .D(n1378), .CLK(CLK), .Q(\memory[14][4] ) );
  DFFPOSX1 \memory_reg[14][3]  ( .D(n1379), .CLK(CLK), .Q(\memory[14][3] ) );
  DFFPOSX1 \memory_reg[14][2]  ( .D(n1380), .CLK(CLK), .Q(\memory[14][2] ) );
  DFFPOSX1 \memory_reg[14][1]  ( .D(n1381), .CLK(CLK), .Q(\memory[14][1] ) );
  DFFPOSX1 \memory_reg[14][0]  ( .D(n1382), .CLK(CLK), .Q(\memory[14][0] ) );
  DFFPOSX1 \memory_reg[15][7]  ( .D(n1367), .CLK(CLK), .Q(\memory[15][7] ) );
  DFFPOSX1 \memory_reg[15][6]  ( .D(n1368), .CLK(CLK), .Q(\memory[15][6] ) );
  DFFPOSX1 \memory_reg[15][5]  ( .D(n1369), .CLK(CLK), .Q(\memory[15][5] ) );
  DFFPOSX1 \memory_reg[15][4]  ( .D(n1370), .CLK(CLK), .Q(\memory[15][4] ) );
  DFFPOSX1 \memory_reg[15][3]  ( .D(n1371), .CLK(CLK), .Q(\memory[15][3] ) );
  DFFPOSX1 \memory_reg[15][2]  ( .D(n1372), .CLK(CLK), .Q(\memory[15][2] ) );
  DFFPOSX1 \memory_reg[15][1]  ( .D(n1373), .CLK(CLK), .Q(\memory[15][1] ) );
  DFFPOSX1 \memory_reg[15][0]  ( .D(n1374), .CLK(CLK), .Q(\memory[15][0] ) );
  DFFPOSX1 \memory_reg[16][7]  ( .D(n1465), .CLK(CLK), .Q(\memory[16][7] ) );
  DFFPOSX1 \memory_reg[16][6]  ( .D(n1466), .CLK(CLK), .Q(\memory[16][6] ) );
  DFFPOSX1 \memory_reg[16][5]  ( .D(n1467), .CLK(CLK), .Q(\memory[16][5] ) );
  DFFPOSX1 \memory_reg[16][4]  ( .D(n1468), .CLK(CLK), .Q(\memory[16][4] ) );
  DFFPOSX1 \memory_reg[16][3]  ( .D(n1469), .CLK(CLK), .Q(\memory[16][3] ) );
  DFFPOSX1 \memory_reg[16][2]  ( .D(n1470), .CLK(CLK), .Q(\memory[16][2] ) );
  DFFPOSX1 \memory_reg[16][1]  ( .D(n1471), .CLK(CLK), .Q(\memory[16][1] ) );
  DFFPOSX1 \memory_reg[16][0]  ( .D(n1472), .CLK(CLK), .Q(\memory[16][0] ) );
  DFFPOSX1 \memory_reg[17][7]  ( .D(n1473), .CLK(CLK), .Q(\memory[17][7] ) );
  DFFPOSX1 \memory_reg[17][6]  ( .D(n1474), .CLK(CLK), .Q(\memory[17][6] ) );
  DFFPOSX1 \memory_reg[17][5]  ( .D(n1475), .CLK(CLK), .Q(\memory[17][5] ) );
  DFFPOSX1 \memory_reg[17][4]  ( .D(n1476), .CLK(CLK), .Q(\memory[17][4] ) );
  DFFPOSX1 \memory_reg[17][3]  ( .D(n1477), .CLK(CLK), .Q(\memory[17][3] ) );
  DFFPOSX1 \memory_reg[17][2]  ( .D(n1478), .CLK(CLK), .Q(\memory[17][2] ) );
  DFFPOSX1 \memory_reg[17][1]  ( .D(n1479), .CLK(CLK), .Q(\memory[17][1] ) );
  DFFPOSX1 \memory_reg[17][0]  ( .D(n1480), .CLK(CLK), .Q(\memory[17][0] ) );
  DFFPOSX1 \memory_reg[18][7]  ( .D(n1481), .CLK(CLK), .Q(\memory[18][7] ) );
  DFFPOSX1 \memory_reg[18][6]  ( .D(n1482), .CLK(CLK), .Q(\memory[18][6] ) );
  DFFPOSX1 \memory_reg[18][5]  ( .D(n1483), .CLK(CLK), .Q(\memory[18][5] ) );
  DFFPOSX1 \memory_reg[18][4]  ( .D(n1484), .CLK(CLK), .Q(\memory[18][4] ) );
  DFFPOSX1 \memory_reg[18][3]  ( .D(n1485), .CLK(CLK), .Q(\memory[18][3] ) );
  DFFPOSX1 \memory_reg[18][2]  ( .D(n1486), .CLK(CLK), .Q(\memory[18][2] ) );
  DFFPOSX1 \memory_reg[18][1]  ( .D(n1487), .CLK(CLK), .Q(\memory[18][1] ) );
  DFFPOSX1 \memory_reg[18][0]  ( .D(n1488), .CLK(CLK), .Q(\memory[18][0] ) );
  DFFPOSX1 \memory_reg[19][7]  ( .D(n1489), .CLK(CLK), .Q(\memory[19][7] ) );
  DFFPOSX1 \memory_reg[19][6]  ( .D(n1490), .CLK(CLK), .Q(\memory[19][6] ) );
  DFFPOSX1 \memory_reg[19][5]  ( .D(n1491), .CLK(CLK), .Q(\memory[19][5] ) );
  DFFPOSX1 \memory_reg[19][4]  ( .D(n1492), .CLK(CLK), .Q(\memory[19][4] ) );
  DFFPOSX1 \memory_reg[19][3]  ( .D(n1493), .CLK(CLK), .Q(\memory[19][3] ) );
  DFFPOSX1 \memory_reg[19][2]  ( .D(n1494), .CLK(CLK), .Q(\memory[19][2] ) );
  DFFPOSX1 \memory_reg[19][1]  ( .D(n1495), .CLK(CLK), .Q(\memory[19][1] ) );
  DFFPOSX1 \memory_reg[19][0]  ( .D(n1496), .CLK(CLK), .Q(\memory[19][0] ) );
  DFFPOSX1 \memory_reg[20][7]  ( .D(n1359), .CLK(CLK), .Q(\memory[20][7] ) );
  DFFPOSX1 \memory_reg[20][6]  ( .D(n1360), .CLK(CLK), .Q(\memory[20][6] ) );
  DFFPOSX1 \memory_reg[20][5]  ( .D(n1361), .CLK(CLK), .Q(\memory[20][5] ) );
  DFFPOSX1 \memory_reg[20][4]  ( .D(n1362), .CLK(CLK), .Q(\memory[20][4] ) );
  DFFPOSX1 \memory_reg[20][3]  ( .D(n1363), .CLK(CLK), .Q(\memory[20][3] ) );
  DFFPOSX1 \memory_reg[20][2]  ( .D(n1364), .CLK(CLK), .Q(\memory[20][2] ) );
  DFFPOSX1 \memory_reg[20][1]  ( .D(n1365), .CLK(CLK), .Q(\memory[20][1] ) );
  DFFPOSX1 \memory_reg[20][0]  ( .D(n1366), .CLK(CLK), .Q(\memory[20][0] ) );
  DFFPOSX1 \memory_reg[21][7]  ( .D(n1351), .CLK(CLK), .Q(\memory[21][7] ) );
  DFFPOSX1 \memory_reg[21][6]  ( .D(n1352), .CLK(CLK), .Q(\memory[21][6] ) );
  DFFPOSX1 \memory_reg[21][5]  ( .D(n1353), .CLK(CLK), .Q(\memory[21][5] ) );
  DFFPOSX1 \memory_reg[21][4]  ( .D(n1354), .CLK(CLK), .Q(\memory[21][4] ) );
  DFFPOSX1 \memory_reg[21][3]  ( .D(n1355), .CLK(CLK), .Q(\memory[21][3] ) );
  DFFPOSX1 \memory_reg[21][2]  ( .D(n1356), .CLK(CLK), .Q(\memory[21][2] ) );
  DFFPOSX1 \memory_reg[21][1]  ( .D(n1357), .CLK(CLK), .Q(\memory[21][1] ) );
  DFFPOSX1 \memory_reg[21][0]  ( .D(n1358), .CLK(CLK), .Q(\memory[21][0] ) );
  DFFPOSX1 \memory_reg[22][7]  ( .D(n1343), .CLK(CLK), .Q(\memory[22][7] ) );
  DFFPOSX1 \memory_reg[22][6]  ( .D(n1344), .CLK(CLK), .Q(\memory[22][6] ) );
  DFFPOSX1 \memory_reg[22][5]  ( .D(n1345), .CLK(CLK), .Q(\memory[22][5] ) );
  DFFPOSX1 \memory_reg[22][4]  ( .D(n1346), .CLK(CLK), .Q(\memory[22][4] ) );
  DFFPOSX1 \memory_reg[22][3]  ( .D(n1347), .CLK(CLK), .Q(\memory[22][3] ) );
  DFFPOSX1 \memory_reg[22][2]  ( .D(n1348), .CLK(CLK), .Q(\memory[22][2] ) );
  DFFPOSX1 \memory_reg[22][1]  ( .D(n1349), .CLK(CLK), .Q(\memory[22][1] ) );
  DFFPOSX1 \memory_reg[22][0]  ( .D(n1350), .CLK(CLK), .Q(\memory[22][0] ) );
  DFFPOSX1 \memory_reg[23][7]  ( .D(n1335), .CLK(CLK), .Q(\memory[23][7] ) );
  DFFPOSX1 \memory_reg[23][6]  ( .D(n1336), .CLK(CLK), .Q(\memory[23][6] ) );
  DFFPOSX1 \memory_reg[23][5]  ( .D(n1337), .CLK(CLK), .Q(\memory[23][5] ) );
  DFFPOSX1 \memory_reg[23][4]  ( .D(n1338), .CLK(CLK), .Q(\memory[23][4] ) );
  DFFPOSX1 \memory_reg[23][3]  ( .D(n1339), .CLK(CLK), .Q(\memory[23][3] ) );
  DFFPOSX1 \memory_reg[23][2]  ( .D(n1340), .CLK(CLK), .Q(\memory[23][2] ) );
  DFFPOSX1 \memory_reg[23][1]  ( .D(n1341), .CLK(CLK), .Q(\memory[23][1] ) );
  DFFPOSX1 \memory_reg[23][0]  ( .D(n1342), .CLK(CLK), .Q(\memory[23][0] ) );
  DFFPOSX1 \memory_reg[24][7]  ( .D(n1327), .CLK(CLK), .Q(\memory[24][7] ) );
  DFFPOSX1 \memory_reg[24][6]  ( .D(n1328), .CLK(CLK), .Q(\memory[24][6] ) );
  DFFPOSX1 \memory_reg[24][5]  ( .D(n1329), .CLK(CLK), .Q(\memory[24][5] ) );
  DFFPOSX1 \memory_reg[24][4]  ( .D(n1330), .CLK(CLK), .Q(\memory[24][4] ) );
  DFFPOSX1 \memory_reg[24][3]  ( .D(n1331), .CLK(CLK), .Q(\memory[24][3] ) );
  DFFPOSX1 \memory_reg[24][2]  ( .D(n1332), .CLK(CLK), .Q(\memory[24][2] ) );
  DFFPOSX1 \memory_reg[24][1]  ( .D(n1333), .CLK(CLK), .Q(\memory[24][1] ) );
  DFFPOSX1 \memory_reg[24][0]  ( .D(n1334), .CLK(CLK), .Q(\memory[24][0] ) );
  DFFPOSX1 \memory_reg[25][7]  ( .D(n1319), .CLK(CLK), .Q(\memory[25][7] ) );
  DFFPOSX1 \memory_reg[25][6]  ( .D(n1320), .CLK(CLK), .Q(\memory[25][6] ) );
  DFFPOSX1 \memory_reg[25][5]  ( .D(n1321), .CLK(CLK), .Q(\memory[25][5] ) );
  DFFPOSX1 \memory_reg[25][4]  ( .D(n1322), .CLK(CLK), .Q(\memory[25][4] ) );
  DFFPOSX1 \memory_reg[25][3]  ( .D(n1323), .CLK(CLK), .Q(\memory[25][3] ) );
  DFFPOSX1 \memory_reg[25][2]  ( .D(n1324), .CLK(CLK), .Q(\memory[25][2] ) );
  DFFPOSX1 \memory_reg[25][1]  ( .D(n1325), .CLK(CLK), .Q(\memory[25][1] ) );
  DFFPOSX1 \memory_reg[25][0]  ( .D(n1326), .CLK(CLK), .Q(\memory[25][0] ) );
  DFFPOSX1 \memory_reg[26][7]  ( .D(n1311), .CLK(CLK), .Q(\memory[26][7] ) );
  DFFPOSX1 \memory_reg[26][6]  ( .D(n1312), .CLK(CLK), .Q(\memory[26][6] ) );
  DFFPOSX1 \memory_reg[26][5]  ( .D(n1313), .CLK(CLK), .Q(\memory[26][5] ) );
  DFFPOSX1 \memory_reg[26][4]  ( .D(n1314), .CLK(CLK), .Q(\memory[26][4] ) );
  DFFPOSX1 \memory_reg[26][3]  ( .D(n1315), .CLK(CLK), .Q(\memory[26][3] ) );
  DFFPOSX1 \memory_reg[26][2]  ( .D(n1316), .CLK(CLK), .Q(\memory[26][2] ) );
  DFFPOSX1 \memory_reg[26][1]  ( .D(n1317), .CLK(CLK), .Q(\memory[26][1] ) );
  DFFPOSX1 \memory_reg[26][0]  ( .D(n1318), .CLK(CLK), .Q(\memory[26][0] ) );
  DFFPOSX1 \memory_reg[27][7]  ( .D(n1303), .CLK(CLK), .Q(\memory[27][7] ) );
  DFFPOSX1 \memory_reg[27][6]  ( .D(n1304), .CLK(CLK), .Q(\memory[27][6] ) );
  DFFPOSX1 \memory_reg[27][5]  ( .D(n1305), .CLK(CLK), .Q(\memory[27][5] ) );
  DFFPOSX1 \memory_reg[27][4]  ( .D(n1306), .CLK(CLK), .Q(\memory[27][4] ) );
  DFFPOSX1 \memory_reg[27][3]  ( .D(n1307), .CLK(CLK), .Q(\memory[27][3] ) );
  DFFPOSX1 \memory_reg[27][2]  ( .D(n1308), .CLK(CLK), .Q(\memory[27][2] ) );
  DFFPOSX1 \memory_reg[27][1]  ( .D(n1309), .CLK(CLK), .Q(\memory[27][1] ) );
  DFFPOSX1 \memory_reg[27][0]  ( .D(n1310), .CLK(CLK), .Q(\memory[27][0] ) );
  DFFPOSX1 \memory_reg[28][7]  ( .D(n1497), .CLK(CLK), .Q(\memory[28][7] ) );
  DFFPOSX1 \memory_reg[28][6]  ( .D(n1498), .CLK(CLK), .Q(\memory[28][6] ) );
  DFFPOSX1 \memory_reg[28][5]  ( .D(n1499), .CLK(CLK), .Q(\memory[28][5] ) );
  DFFPOSX1 \memory_reg[28][4]  ( .D(n1500), .CLK(CLK), .Q(\memory[28][4] ) );
  DFFPOSX1 \memory_reg[28][3]  ( .D(n1501), .CLK(CLK), .Q(\memory[28][3] ) );
  DFFPOSX1 \memory_reg[28][2]  ( .D(n1502), .CLK(CLK), .Q(\memory[28][2] ) );
  DFFPOSX1 \memory_reg[28][1]  ( .D(n1503), .CLK(CLK), .Q(\memory[28][1] ) );
  DFFPOSX1 \memory_reg[28][0]  ( .D(n1504), .CLK(CLK), .Q(\memory[28][0] ) );
  DFFPOSX1 \memory_reg[29][7]  ( .D(n1505), .CLK(CLK), .Q(\memory[29][7] ) );
  DFFPOSX1 \memory_reg[29][6]  ( .D(n1506), .CLK(CLK), .Q(\memory[29][6] ) );
  DFFPOSX1 \memory_reg[29][5]  ( .D(n1507), .CLK(CLK), .Q(\memory[29][5] ) );
  DFFPOSX1 \memory_reg[29][4]  ( .D(n1508), .CLK(CLK), .Q(\memory[29][4] ) );
  DFFPOSX1 \memory_reg[29][3]  ( .D(n1509), .CLK(CLK), .Q(\memory[29][3] ) );
  DFFPOSX1 \memory_reg[29][2]  ( .D(n1510), .CLK(CLK), .Q(\memory[29][2] ) );
  DFFPOSX1 \memory_reg[29][1]  ( .D(n1511), .CLK(CLK), .Q(\memory[29][1] ) );
  DFFPOSX1 \memory_reg[29][0]  ( .D(n1512), .CLK(CLK), .Q(\memory[29][0] ) );
  DFFPOSX1 \memory_reg[30][7]  ( .D(n1513), .CLK(CLK), .Q(\memory[30][7] ) );
  DFFPOSX1 \memory_reg[30][6]  ( .D(n1514), .CLK(CLK), .Q(\memory[30][6] ) );
  DFFPOSX1 \memory_reg[30][5]  ( .D(n1515), .CLK(CLK), .Q(\memory[30][5] ) );
  DFFPOSX1 \memory_reg[30][4]  ( .D(n1516), .CLK(CLK), .Q(\memory[30][4] ) );
  DFFPOSX1 \memory_reg[30][3]  ( .D(n1517), .CLK(CLK), .Q(\memory[30][3] ) );
  DFFPOSX1 \memory_reg[30][2]  ( .D(n1518), .CLK(CLK), .Q(\memory[30][2] ) );
  DFFPOSX1 \memory_reg[30][1]  ( .D(n1519), .CLK(CLK), .Q(\memory[30][1] ) );
  DFFPOSX1 \memory_reg[30][0]  ( .D(n1520), .CLK(CLK), .Q(\memory[30][0] ) );
  DFFPOSX1 \memory_reg[31][7]  ( .D(n1521), .CLK(CLK), .Q(\memory[31][7] ) );
  DFFPOSX1 \memory_reg[31][6]  ( .D(n1522), .CLK(CLK), .Q(\memory[31][6] ) );
  DFFPOSX1 \memory_reg[31][5]  ( .D(n1523), .CLK(CLK), .Q(\memory[31][5] ) );
  DFFPOSX1 \memory_reg[31][4]  ( .D(n1524), .CLK(CLK), .Q(\memory[31][4] ) );
  DFFPOSX1 \memory_reg[31][3]  ( .D(n1525), .CLK(CLK), .Q(\memory[31][3] ) );
  DFFPOSX1 \memory_reg[31][2]  ( .D(n1526), .CLK(CLK), .Q(\memory[31][2] ) );
  DFFPOSX1 \memory_reg[31][1]  ( .D(n1527), .CLK(CLK), .Q(\memory[31][1] ) );
  DFFPOSX1 \memory_reg[31][0]  ( .D(n1528), .CLK(CLK), .Q(\memory[31][0] ) );
  DFFPOSX1 \opcode_reg[0][1]  ( .D(n1296), .CLK(CLK), .Q(\opcode[0][1] ) );
  DFFPOSX1 \opcode_reg[0][0]  ( .D(n1295), .CLK(CLK), .Q(\opcode[0][0] ) );
  DFFPOSX1 \opcode_reg[1][1]  ( .D(n1298), .CLK(CLK), .Q(\opcode[1][1] ) );
  DFFPOSX1 \opcode_reg[1][0]  ( .D(n1297), .CLK(CLK), .Q(\opcode[1][0] ) );
  DFFPOSX1 \opcode_reg[2][1]  ( .D(n1300), .CLK(CLK), .Q(\opcode[2][1] ) );
  DFFPOSX1 \opcode_reg[2][0]  ( .D(n1299), .CLK(CLK), .Q(\opcode[2][0] ) );
  DFFPOSX1 \opcode_reg[3][1]  ( .D(n1302), .CLK(CLK), .Q(\opcode[3][1] ) );
  DFFPOSX1 \opcode_reg[3][0]  ( .D(n1301), .CLK(CLK), .Q(\opcode[3][0] ) );
  DFFPOSX1 \opcode_reg[4][1]  ( .D(n1594), .CLK(CLK), .Q(\opcode[4][1] ) );
  DFFPOSX1 \opcode_reg[4][0]  ( .D(n1593), .CLK(CLK), .Q(\opcode[4][0] ) );
  DFFPOSX1 \opcode_reg[5][1]  ( .D(n1584), .CLK(CLK), .Q(\opcode[5][1] ) );
  DFFPOSX1 \opcode_reg[5][0]  ( .D(n1583), .CLK(CLK), .Q(\opcode[5][0] ) );
  DFFPOSX1 \opcode_reg[6][1]  ( .D(n1574), .CLK(CLK), .Q(\opcode[6][1] ) );
  DFFPOSX1 \opcode_reg[6][0]  ( .D(n1573), .CLK(CLK), .Q(\opcode[6][0] ) );
  DFFPOSX1 \opcode_reg[7][1]  ( .D(n1564), .CLK(CLK), .Q(\opcode[7][1] ) );
  DFFPOSX1 \opcode_reg[7][0]  ( .D(n1563), .CLK(CLK), .Q(\opcode[7][0] ) );
  DFFPOSX1 \opcode_reg[8][1]  ( .D(n1529), .CLK(CLK), .Q(\opcode[8][1] ) );
  DFFPOSX1 \opcode_reg[8][0]  ( .D(n1530), .CLK(CLK), .Q(\opcode[8][0] ) );
  DFFPOSX1 \opcode_reg[9][1]  ( .D(n1531), .CLK(CLK), .Q(\opcode[9][1] ) );
  DFFPOSX1 \opcode_reg[9][0]  ( .D(n1532), .CLK(CLK), .Q(\opcode[9][0] ) );
  DFFPOSX1 \opcode_reg[10][1]  ( .D(n1533), .CLK(CLK), .Q(\opcode[10][1] ) );
  DFFPOSX1 \opcode_reg[10][0]  ( .D(n1534), .CLK(CLK), .Q(\opcode[10][0] ) );
  DFFPOSX1 \opcode_reg[11][1]  ( .D(n1535), .CLK(CLK), .Q(\opcode[11][1] ) );
  DFFPOSX1 \opcode_reg[11][0]  ( .D(n1536), .CLK(CLK), .Q(\opcode[11][0] ) );
  DFFPOSX1 \opcode_reg[12][1]  ( .D(n1293), .CLK(CLK), .Q(\opcode[12][1] ) );
  DFFPOSX1 \opcode_reg[12][0]  ( .D(n1294), .CLK(CLK), .Q(\opcode[12][0] ) );
  DFFPOSX1 \opcode_reg[13][1]  ( .D(n1291), .CLK(CLK), .Q(\opcode[13][1] ) );
  DFFPOSX1 \opcode_reg[13][0]  ( .D(n1292), .CLK(CLK), .Q(\opcode[13][0] ) );
  DFFPOSX1 \opcode_reg[14][1]  ( .D(n1289), .CLK(CLK), .Q(\opcode[14][1] ) );
  DFFPOSX1 \opcode_reg[14][0]  ( .D(n1290), .CLK(CLK), .Q(\opcode[14][0] ) );
  DFFPOSX1 \opcode_reg[15][1]  ( .D(n1287), .CLK(CLK), .Q(\opcode[15][1] ) );
  DFFPOSX1 \opcode_reg[15][0]  ( .D(n1288), .CLK(CLK), .Q(\opcode[15][0] ) );
  DFFPOSX1 \opcode_reg[16][1]  ( .D(n1537), .CLK(CLK), .Q(\opcode[16][1] ) );
  DFFPOSX1 \opcode_reg[16][0]  ( .D(n1538), .CLK(CLK), .Q(\opcode[16][0] ) );
  DFFPOSX1 \opcode_reg[17][1]  ( .D(n1539), .CLK(CLK), .Q(\opcode[17][1] ) );
  DFFPOSX1 \opcode_reg[17][0]  ( .D(n1540), .CLK(CLK), .Q(\opcode[17][0] ) );
  DFFPOSX1 \opcode_reg[18][1]  ( .D(n1541), .CLK(CLK), .Q(\opcode[18][1] ) );
  DFFPOSX1 \opcode_reg[18][0]  ( .D(n1542), .CLK(CLK), .Q(\opcode[18][0] ) );
  DFFPOSX1 \opcode_reg[19][1]  ( .D(n1543), .CLK(CLK), .Q(\opcode[19][1] ) );
  DFFPOSX1 \opcode_reg[19][0]  ( .D(n1544), .CLK(CLK), .Q(\opcode[19][0] ) );
  DFFPOSX1 \opcode_reg[20][1]  ( .D(n1285), .CLK(CLK), .Q(\opcode[20][1] ) );
  DFFPOSX1 \opcode_reg[20][0]  ( .D(n1286), .CLK(CLK), .Q(\opcode[20][0] ) );
  DFFPOSX1 \opcode_reg[21][1]  ( .D(n1283), .CLK(CLK), .Q(\opcode[21][1] ) );
  DFFPOSX1 \opcode_reg[21][0]  ( .D(n1284), .CLK(CLK), .Q(\opcode[21][0] ) );
  DFFPOSX1 \opcode_reg[22][1]  ( .D(n1281), .CLK(CLK), .Q(\opcode[22][1] ) );
  DFFPOSX1 \opcode_reg[22][0]  ( .D(n1282), .CLK(CLK), .Q(\opcode[22][0] ) );
  DFFPOSX1 \opcode_reg[23][1]  ( .D(n1279), .CLK(CLK), .Q(\opcode[23][1] ) );
  DFFPOSX1 \opcode_reg[23][0]  ( .D(n1280), .CLK(CLK), .Q(\opcode[23][0] ) );
  DFFPOSX1 \opcode_reg[24][1]  ( .D(n1277), .CLK(CLK), .Q(\opcode[24][1] ) );
  DFFPOSX1 \opcode_reg[24][0]  ( .D(n1278), .CLK(CLK), .Q(\opcode[24][0] ) );
  DFFPOSX1 \opcode_reg[25][1]  ( .D(n1275), .CLK(CLK), .Q(\opcode[25][1] ) );
  DFFPOSX1 \opcode_reg[25][0]  ( .D(n1276), .CLK(CLK), .Q(\opcode[25][0] ) );
  DFFPOSX1 \opcode_reg[26][1]  ( .D(n1273), .CLK(CLK), .Q(\opcode[26][1] ) );
  DFFPOSX1 \opcode_reg[26][0]  ( .D(n1274), .CLK(CLK), .Q(\opcode[26][0] ) );
  DFFPOSX1 \opcode_reg[27][1]  ( .D(n1271), .CLK(CLK), .Q(\opcode[27][1] ) );
  DFFPOSX1 \opcode_reg[27][0]  ( .D(n1272), .CLK(CLK), .Q(\opcode[27][0] ) );
  DFFPOSX1 \opcode_reg[28][1]  ( .D(n1545), .CLK(CLK), .Q(\opcode[28][1] ) );
  DFFPOSX1 \opcode_reg[28][0]  ( .D(n1546), .CLK(CLK), .Q(\opcode[28][0] ) );
  DFFPOSX1 \opcode_reg[29][1]  ( .D(n1547), .CLK(CLK), .Q(\opcode[29][1] ) );
  DFFPOSX1 \opcode_reg[29][0]  ( .D(n1548), .CLK(CLK), .Q(\opcode[29][0] ) );
  DFFPOSX1 \opcode_reg[30][1]  ( .D(n1549), .CLK(CLK), .Q(\opcode[30][1] ) );
  DFFPOSX1 \opcode_reg[30][0]  ( .D(n1550), .CLK(CLK), .Q(\opcode[30][0] ) );
  DFFPOSX1 \opcode_reg[31][1]  ( .D(n1551), .CLK(CLK), .Q(\opcode[31][1] ) );
  DFFPOSX1 \opcode_reg[31][0]  ( .D(n1552), .CLK(CLK), .Q(\opcode[31][0] ) );
  DFFPOSX1 \DATA_reg[7]  ( .D(n1553), .CLK(CLK), .Q(DATA[7]) );
  DFFPOSX1 \DATA_reg[6]  ( .D(n1554), .CLK(CLK), .Q(DATA[6]) );
  DFFPOSX1 \DATA_reg[5]  ( .D(n1555), .CLK(CLK), .Q(DATA[5]) );
  DFFPOSX1 \DATA_reg[4]  ( .D(n1556), .CLK(CLK), .Q(DATA[4]) );
  DFFPOSX1 \DATA_reg[3]  ( .D(n1557), .CLK(CLK), .Q(DATA[3]) );
  DFFPOSX1 \DATA_reg[2]  ( .D(n1558), .CLK(CLK), .Q(DATA[2]) );
  DFFPOSX1 \DATA_reg[1]  ( .D(n1559), .CLK(CLK), .Q(DATA[1]) );
  DFFPOSX1 \DATA_reg[0]  ( .D(n1560), .CLK(CLK), .Q(DATA[0]) );
  DFFPOSX1 \OUT_OPCODE_reg[1]  ( .D(n1561), .CLK(CLK), .Q(OUT_OPCODE[1]) );
  DFFPOSX1 \OUT_OPCODE_reg[0]  ( .D(n1562), .CLK(CLK), .Q(OUT_OPCODE[0]) );
  DFFPOSX1 EMPTY_reg ( .D(n1432), .CLK(CLK), .Q(EMPTY) );
  DFFSR \readptr_reg[2]  ( .D(N345), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        readptr[2]) );
  DFFSR \readptr_reg[4]  ( .D(N347), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        readptr[4]) );
  DFFSR \writeptr_reg[4]  ( .D(n1607), .CLK(CLK), .R(n163), .S(1'b1), .Q(
        writeptr[4]) );
  INVX2 U3 ( .A(n17), .Y(n127) );
  INVX2 U4 ( .A(writeptr[0]), .Y(n132) );
  INVX1 U5 ( .A(n88), .Y(n40) );
  XOR2X1 U6 ( .A(n46), .B(n134), .Y(n575) );
  INVX2 U7 ( .A(n46), .Y(n131) );
  XNOR2X1 U8 ( .A(n101), .B(n135), .Y(n82) );
  INVX4 U9 ( .A(n135), .Y(n136) );
  INVX2 U10 ( .A(n534), .Y(n542) );
  NAND2X1 U11 ( .A(RCV_OPCODE[1]), .B(RCV_OPCODE[0]), .Y(n1) );
  NAND2X1 U12 ( .A(RCV_OPCODE[1]), .B(RCV_OPCODE[0]), .Y(n2) );
  INVX2 U13 ( .A(n1), .Y(n3) );
  NAND2X1 U14 ( .A(n2), .B(n230), .Y(n4) );
  NAND2X1 U15 ( .A(n1), .B(n241), .Y(n5) );
  AND2X2 U16 ( .A(n209), .B(n218), .Y(n6) );
  INVX1 U17 ( .A(n331), .Y(n115) );
  AND2X2 U18 ( .A(n1237), .B(n1247), .Y(n7) );
  AND2X2 U19 ( .A(n1267), .B(n1237), .Y(n8) );
  AND2X1 U20 ( .A(n1258), .B(n1237), .Y(n9) );
  AND2X2 U21 ( .A(n1267), .B(n86), .Y(n10) );
  AND2X1 U22 ( .A(n1237), .B(n1248), .Y(n11) );
  AND2X1 U23 ( .A(n1238), .B(n1237), .Y(n12) );
  AND2X1 U24 ( .A(n1238), .B(n86), .Y(n13) );
  AND2X1 U25 ( .A(n1248), .B(n86), .Y(n14) );
  AND2X1 U26 ( .A(n1259), .B(n86), .Y(n15) );
  AND2X2 U27 ( .A(n1259), .B(n1237), .Y(n16) );
  AND2X2 U28 ( .A(n1268), .B(n1237), .Y(n17) );
  AND2X2 U29 ( .A(n1268), .B(n86), .Y(n18) );
  INVX1 U30 ( .A(RCV_DATA[5]), .Y(n540) );
  INVX1 U31 ( .A(RCV_DATA[0]), .Y(n535) );
  INVX1 U32 ( .A(RCV_DATA[2]), .Y(n537) );
  INVX1 U33 ( .A(RCV_DATA[3]), .Y(n538) );
  INVX1 U34 ( .A(RCV_DATA[4]), .Y(n539) );
  NAND2X1 U38 ( .A(n227), .B(n161), .Y(n22) );
  NAND2X1 U39 ( .A(n251), .B(n161), .Y(n23) );
  NAND3X1 U40 ( .A(n66), .B(n64), .C(n191), .Y(n24) );
  INVX1 U41 ( .A(RCV_DATA[1]), .Y(n536) );
  NAND2X1 U42 ( .A(readptr[0]), .B(n219), .Y(n25) );
  INVX2 U43 ( .A(n134), .Y(n219) );
  NAND2X1 U44 ( .A(n293), .B(n161), .Y(n26) );
  INVX2 U45 ( .A(n247), .Y(n249) );
  NAND2X1 U46 ( .A(n276), .B(n160), .Y(n27) );
  INVX1 U47 ( .A(RCV_DATA[6]), .Y(n541) );
  INVX1 U48 ( .A(n575), .Y(n576) );
  OR2X1 U49 ( .A(n132), .B(n129), .Y(n28) );
  XNOR2X1 U50 ( .A(n569), .B(n51), .Y(n64) );
  INVX2 U51 ( .A(n618), .Y(n51) );
  BUFX2 U52 ( .A(n67), .Y(n29) );
  NAND2X1 U53 ( .A(n261), .B(n160), .Y(n30) );
  NAND3X1 U54 ( .A(n70), .B(n134), .C(n130), .Y(n31) );
  INVX2 U55 ( .A(n322), .Y(n323) );
  NAND2X1 U56 ( .A(n160), .B(n296), .Y(n32) );
  NAND2X1 U57 ( .A(n265), .B(n161), .Y(n33) );
  NOR2X1 U58 ( .A(n614), .B(n57), .Y(n34) );
  INVX1 U59 ( .A(n34), .Y(n612) );
  NAND2X1 U60 ( .A(n193), .B(n160), .Y(n35) );
  NAND2X1 U61 ( .A(n160), .B(n220), .Y(n36) );
  NAND2X1 U62 ( .A(n161), .B(n210), .Y(n37) );
  NAND2X1 U63 ( .A(n160), .B(n246), .Y(n38) );
  NAND2X1 U64 ( .A(n161), .B(n254), .Y(n39) );
  INVX8 U65 ( .A(n128), .Y(n70) );
  INVX2 U66 ( .A(n297), .Y(n298) );
  AND2X2 U67 ( .A(n40), .B(n41), .Y(n166) );
  INVX1 U68 ( .A(n41), .Y(n543) );
  INVX2 U69 ( .A(n266), .Y(n268) );
  MUX2X1 U70 ( .B(n116), .A(n321), .S(n3), .Y(n287) );
  INVX4 U71 ( .A(n480), .Y(n481) );
  INVX4 U72 ( .A(n448), .Y(n456) );
  AND2X2 U73 ( .A(n545), .B(n164), .Y(n41) );
  NAND2X1 U74 ( .A(n83), .B(W_ENABLE), .Y(n42) );
  INVX8 U75 ( .A(n162), .Y(n161) );
  BUFX4 U76 ( .A(readptr[2]), .Y(n43) );
  INVX1 U77 ( .A(n189), .Y(n44) );
  INVX2 U78 ( .A(n44), .Y(n45) );
  INVX4 U79 ( .A(n488), .Y(n496) );
  INVX4 U80 ( .A(n528), .Y(n529) );
  INVX4 U81 ( .A(n518), .Y(n526) );
  INVX4 U82 ( .A(n530), .Y(n531) );
  INVX1 U83 ( .A(writeptr[1]), .Y(n46) );
  INVX8 U84 ( .A(n132), .Y(n134) );
  INVX4 U85 ( .A(n508), .Y(n516) );
  INVX4 U86 ( .A(n532), .Y(n533) );
  INVX1 U87 ( .A(RCV_OPCODE[1]), .Y(n341) );
  AND2X2 U88 ( .A(n49), .B(n618), .Y(n86) );
  AND2X2 U89 ( .A(n49), .B(n43), .Y(n87) );
  OR2X2 U90 ( .A(n68), .B(n42), .Y(n47) );
  BUFX2 U91 ( .A(n592), .Y(n48) );
  BUFX4 U92 ( .A(readptr[1]), .Y(n49) );
  INVX4 U93 ( .A(n57), .Y(n50) );
  INVX2 U94 ( .A(readptr[0]), .Y(n57) );
  INVX2 U95 ( .A(n115), .Y(n116) );
  INVX4 U96 ( .A(n568), .Y(n162) );
  BUFX2 U97 ( .A(writeptr[4]), .Y(n52) );
  INVX1 U98 ( .A(n31), .Y(n117) );
  INVX2 U99 ( .A(n620), .Y(n53) );
  INVX2 U100 ( .A(readptr[4]), .Y(n620) );
  NAND2X1 U101 ( .A(n116), .B(n45), .Y(n54) );
  NAND2X1 U102 ( .A(W_ENABLE), .B(n83), .Y(n55) );
  BUFX2 U103 ( .A(n29), .Y(n56) );
  INVX1 U104 ( .A(readptr[0]), .Y(n617) );
  INVX2 U105 ( .A(n226), .Y(n58) );
  INVX4 U106 ( .A(n58), .Y(n59) );
  INVX2 U107 ( .A(n260), .Y(n60) );
  INVX4 U108 ( .A(n60), .Y(n61) );
  AND2X2 U109 ( .A(n52), .B(n264), .Y(n89) );
  AND2X2 U110 ( .A(n52), .B(n73), .Y(n90) );
  INVX1 U111 ( .A(writeptr[4]), .Y(n591) );
  INVX4 U112 ( .A(n498), .Y(n506) );
  NAND2X1 U113 ( .A(n160), .B(n290), .Y(n62) );
  NOR2X1 U114 ( .A(n129), .B(n132), .Y(n63) );
  INVX2 U115 ( .A(writeptr[1]), .Y(n129) );
  INVX1 U116 ( .A(n64), .Y(n561) );
  NAND2X1 U117 ( .A(n161), .B(n281), .Y(n65) );
  BUFX4 U118 ( .A(n305), .Y(n91) );
  BUFX4 U119 ( .A(n305), .Y(n92) );
  BUFX4 U120 ( .A(n236), .Y(n94) );
  BUFX4 U121 ( .A(n336), .Y(n96) );
  BUFX4 U122 ( .A(n271), .Y(n98) );
  INVX4 U123 ( .A(n32), .Y(n487) );
  INVX1 U124 ( .A(n67), .Y(n579) );
  INVX4 U125 ( .A(n30), .Y(n437) );
  INVX4 U126 ( .A(n23), .Y(n431) );
  INVX4 U127 ( .A(n390), .Y(n398) );
  INVX4 U128 ( .A(n22), .Y(n389) );
  NOR2X1 U129 ( .A(n41), .B(n190), .Y(n66) );
  INVX4 U130 ( .A(n382), .Y(n383) );
  INVX4 U131 ( .A(n70), .Y(n218) );
  INVX4 U132 ( .A(n35), .Y(n350) );
  INVX4 U133 ( .A(n38), .Y(n428) );
  INVX4 U134 ( .A(n37), .Y(n380) );
  INVX4 U135 ( .A(n39), .Y(n433) );
  INVX4 U136 ( .A(n36), .Y(n385) );
  INVX4 U137 ( .A(n434), .Y(n435) );
  INVX4 U138 ( .A(n386), .Y(n387) );
  INVX4 U139 ( .A(n410), .Y(n418) );
  INVX4 U140 ( .A(n362), .Y(n370) );
  INVX4 U141 ( .A(n400), .Y(n408) );
  INVX4 U142 ( .A(n352), .Y(n360) );
  INVX4 U143 ( .A(n65), .Y(n476) );
  INVX2 U144 ( .A(n24), .Y(n68) );
  INVX4 U145 ( .A(n27), .Y(n466) );
  INVX4 U146 ( .A(n26), .Y(n485) );
  INVX4 U147 ( .A(n62), .Y(n483) );
  INVX4 U148 ( .A(n33), .Y(n446) );
  AND2X2 U149 ( .A(n24), .B(W_ENABLE), .Y(n67) );
  OR2X1 U150 ( .A(n316), .B(n55), .Y(n69) );
  OR2X2 U151 ( .A(n68), .B(n71), .Y(n478) );
  NAND2X1 U152 ( .A(n83), .B(W_ENABLE), .Y(n71) );
  INVX1 U153 ( .A(n478), .Y(n479) );
  INVX8 U154 ( .A(n162), .Y(n160) );
  INVX2 U155 ( .A(n14), .Y(n105) );
  INVX2 U156 ( .A(n341), .Y(n143) );
  INVX2 U157 ( .A(n11), .Y(n123) );
  INVX2 U158 ( .A(n9), .Y(n124) );
  INVX1 U159 ( .A(n802), .Y(n106) );
  INVX2 U160 ( .A(n13), .Y(n102) );
  INVX2 U161 ( .A(n15), .Y(n108) );
  INVX2 U162 ( .A(n139), .Y(n137) );
  INVX2 U163 ( .A(n139), .Y(n138) );
  INVX2 U164 ( .A(n339), .Y(n139) );
  INVX2 U165 ( .A(n143), .Y(n140) );
  INVX2 U166 ( .A(n143), .Y(n141) );
  BUFX2 U167 ( .A(n336), .Y(n95) );
  INVX2 U168 ( .A(n143), .Y(n142) );
  AND2X2 U169 ( .A(RCV_OPCODE[0]), .B(RCV_OPCODE[1]), .Y(n72) );
  BUFX2 U170 ( .A(n271), .Y(n97) );
  BUFX2 U171 ( .A(n236), .Y(n93) );
  INVX2 U172 ( .A(n6), .Y(n118) );
  NOR2X1 U173 ( .A(RST), .B(n100), .Y(n73) );
  INVX2 U174 ( .A(RST), .Y(n163) );
  AND2X2 U175 ( .A(n1268), .B(n87), .Y(n74) );
  AND2X2 U176 ( .A(n1238), .B(n87), .Y(n75) );
  AND2X2 U177 ( .A(n1259), .B(n87), .Y(n76) );
  AND2X2 U178 ( .A(n1248), .B(n87), .Y(n77) );
  AND2X2 U179 ( .A(n1267), .B(n87), .Y(n78) );
  AND2X2 U180 ( .A(n1236), .B(n87), .Y(n79) );
  AND2X2 U181 ( .A(n1247), .B(n87), .Y(n80) );
  AND2X2 U182 ( .A(n1258), .B(n87), .Y(n81) );
  XOR2X1 U183 ( .A(n586), .B(n82), .Y(n562) );
  XNOR2X1 U184 ( .A(n592), .B(n558), .Y(n563) );
  INVX1 U185 ( .A(n219), .Y(n133) );
  INVX2 U186 ( .A(n7), .Y(n122) );
  INVX4 U187 ( .A(n8), .Y(n126) );
  INVX2 U188 ( .A(n119), .Y(n120) );
  INVX1 U189 ( .A(n793), .Y(n119) );
  INVX4 U190 ( .A(n16), .Y(n125) );
  INVX2 U191 ( .A(n12), .Y(n121) );
  INVX4 U192 ( .A(n10), .Y(n112) );
  INVX2 U193 ( .A(n103), .Y(n104) );
  INVX1 U194 ( .A(n794), .Y(n103) );
  INVX2 U195 ( .A(n106), .Y(n107) );
  INVX2 U196 ( .A(n109), .Y(n110) );
  INVX1 U197 ( .A(n812), .Y(n109) );
  INVX4 U198 ( .A(n18), .Y(n111) );
  INVX4 U199 ( .A(n129), .Y(n130) );
  AND2X2 U200 ( .A(n264), .B(n591), .Y(n83) );
  AND2X2 U201 ( .A(n73), .B(n591), .Y(n84) );
  INVX2 U202 ( .A(n85), .Y(n113) );
  INVX2 U203 ( .A(n85), .Y(n114) );
  INVX2 U204 ( .A(n145), .Y(n144) );
  INVX2 U205 ( .A(n147), .Y(n146) );
  INVX2 U206 ( .A(n149), .Y(n148) );
  INVX2 U207 ( .A(n151), .Y(n150) );
  INVX2 U208 ( .A(n153), .Y(n152) );
  INVX2 U209 ( .A(n157), .Y(n156) );
  INVX2 U210 ( .A(RCV_DATA[7]), .Y(n158) );
  INVX2 U211 ( .A(RCV_DATA[7]), .Y(n159) );
  INVX2 U212 ( .A(n155), .Y(n154) );
  OR2X2 U213 ( .A(n614), .B(n168), .Y(n85) );
  XOR2X1 U214 ( .A(n130), .B(n49), .Y(n88) );
  INVX2 U215 ( .A(readptr[3]), .Y(n135) );
  INVX2 U216 ( .A(n538), .Y(n151) );
  INVX2 U217 ( .A(n540), .Y(n155) );
  INVX2 U218 ( .A(n535), .Y(n145) );
  INVX2 U219 ( .A(n536), .Y(n147) );
  INVX2 U220 ( .A(n537), .Y(n149) );
  INVX2 U221 ( .A(n539), .Y(n153) );
  INVX2 U222 ( .A(n541), .Y(n157) );
  INVX2 U223 ( .A(writeptr[3]), .Y(n99) );
  INVX2 U224 ( .A(n99), .Y(n100) );
  INVX2 U225 ( .A(n99), .Y(n101) );
  INVX1 U226 ( .A(n100), .Y(n587) );
  INVX2 U227 ( .A(writeptr[2]), .Y(n128) );
  AND2X2 U228 ( .A(n1238), .B(n1239), .Y(n796) );
  AND2X2 U229 ( .A(n1236), .B(n1239), .Y(n795) );
  AND2X2 U230 ( .A(n1239), .B(n1248), .Y(n804) );
  AND2X2 U231 ( .A(n1239), .B(n1247), .Y(n803) );
  AND2X2 U232 ( .A(n1259), .B(n1239), .Y(n814) );
  AND2X2 U233 ( .A(n1258), .B(n1239), .Y(n813) );
  AND2X2 U234 ( .A(n1268), .B(n1239), .Y(n821) );
  AND2X2 U235 ( .A(n1267), .B(n1239), .Y(n820) );
  INVX2 U236 ( .A(\memory[16][7] ), .Y(n735) );
  INVX2 U237 ( .A(\memory[17][7] ), .Y(n743) );
  INVX2 U238 ( .A(\memory[18][7] ), .Y(n751) );
  INVX2 U239 ( .A(readptr[2]), .Y(n618) );
  INVX2 U240 ( .A(\memory[19][7] ), .Y(n759) );
  NAND2X1 U241 ( .A(n1236), .B(n86), .Y(n794) );
  INVX2 U242 ( .A(\memory[24][7] ), .Y(n661) );
  INVX2 U243 ( .A(\memory[25][7] ), .Y(n653) );
  INVX2 U244 ( .A(\memory[26][7] ), .Y(n645) );
  INVX2 U245 ( .A(\memory[27][7] ), .Y(n637) );
  NAND2X1 U246 ( .A(n1247), .B(n86), .Y(n802) );
  INVX2 U247 ( .A(\memory[3][7] ), .Y(n700) );
  INVX2 U248 ( .A(\memory[2][7] ), .Y(n692) );
  NAND2X1 U249 ( .A(n1258), .B(n86), .Y(n812) );
  INVX2 U250 ( .A(\memory[1][7] ), .Y(n684) );
  INVX2 U251 ( .A(\memory[0][7] ), .Y(n676) );
  INVX2 U252 ( .A(\memory[8][7] ), .Y(n703) );
  INVX2 U253 ( .A(\memory[9][7] ), .Y(n711) );
  INVX2 U254 ( .A(\memory[10][7] ), .Y(n719) );
  INVX2 U255 ( .A(\memory[11][7] ), .Y(n727) );
  INVX2 U256 ( .A(\memory[16][6] ), .Y(n736) );
  INVX2 U257 ( .A(\memory[17][6] ), .Y(n744) );
  INVX2 U258 ( .A(\memory[18][6] ), .Y(n752) );
  INVX2 U259 ( .A(\memory[19][6] ), .Y(n760) );
  INVX2 U260 ( .A(\memory[24][6] ), .Y(n662) );
  INVX2 U261 ( .A(\memory[25][6] ), .Y(n654) );
  INVX2 U262 ( .A(\memory[26][6] ), .Y(n646) );
  INVX2 U263 ( .A(\memory[27][6] ), .Y(n638) );
  INVX2 U264 ( .A(\memory[3][6] ), .Y(n699) );
  INVX2 U265 ( .A(\memory[2][6] ), .Y(n691) );
  INVX2 U266 ( .A(\memory[1][6] ), .Y(n683) );
  INVX2 U267 ( .A(\memory[0][6] ), .Y(n675) );
  INVX2 U268 ( .A(\memory[8][6] ), .Y(n704) );
  INVX2 U269 ( .A(\memory[9][6] ), .Y(n712) );
  INVX2 U270 ( .A(\memory[10][6] ), .Y(n720) );
  INVX2 U271 ( .A(\memory[11][6] ), .Y(n728) );
  INVX2 U272 ( .A(\memory[16][5] ), .Y(n737) );
  INVX2 U273 ( .A(\memory[17][5] ), .Y(n745) );
  INVX2 U274 ( .A(\memory[18][5] ), .Y(n753) );
  INVX2 U275 ( .A(\memory[19][5] ), .Y(n761) );
  INVX2 U276 ( .A(\memory[24][5] ), .Y(n663) );
  INVX2 U277 ( .A(\memory[25][5] ), .Y(n655) );
  INVX2 U278 ( .A(\memory[26][5] ), .Y(n647) );
  INVX2 U279 ( .A(\memory[27][5] ), .Y(n639) );
  INVX2 U280 ( .A(\memory[3][5] ), .Y(n698) );
  INVX2 U281 ( .A(\memory[2][5] ), .Y(n690) );
  INVX2 U282 ( .A(\memory[1][5] ), .Y(n682) );
  INVX2 U283 ( .A(\memory[0][5] ), .Y(n674) );
  INVX2 U284 ( .A(\memory[8][5] ), .Y(n705) );
  INVX2 U285 ( .A(\memory[9][5] ), .Y(n713) );
  INVX2 U286 ( .A(\memory[10][5] ), .Y(n721) );
  INVX2 U287 ( .A(\memory[11][5] ), .Y(n729) );
  INVX2 U288 ( .A(\memory[16][4] ), .Y(n738) );
  INVX2 U289 ( .A(\memory[17][4] ), .Y(n746) );
  INVX2 U290 ( .A(\memory[18][4] ), .Y(n754) );
  INVX2 U291 ( .A(\memory[19][4] ), .Y(n762) );
  INVX2 U292 ( .A(\memory[24][4] ), .Y(n664) );
  INVX2 U293 ( .A(\memory[25][4] ), .Y(n656) );
  INVX2 U294 ( .A(\memory[26][4] ), .Y(n648) );
  INVX2 U295 ( .A(\memory[27][4] ), .Y(n640) );
  INVX2 U296 ( .A(\memory[3][4] ), .Y(n697) );
  INVX2 U297 ( .A(\memory[2][4] ), .Y(n689) );
  INVX2 U298 ( .A(\memory[1][4] ), .Y(n681) );
  INVX2 U299 ( .A(\memory[0][4] ), .Y(n673) );
  INVX2 U300 ( .A(\memory[8][4] ), .Y(n706) );
  INVX2 U301 ( .A(\memory[9][4] ), .Y(n714) );
  INVX2 U302 ( .A(\memory[10][4] ), .Y(n722) );
  INVX2 U303 ( .A(\memory[11][4] ), .Y(n730) );
  INVX2 U304 ( .A(\memory[16][3] ), .Y(n739) );
  INVX2 U305 ( .A(\memory[17][3] ), .Y(n747) );
  INVX2 U306 ( .A(\memory[18][3] ), .Y(n755) );
  INVX2 U307 ( .A(\memory[19][3] ), .Y(n763) );
  INVX2 U308 ( .A(\memory[24][3] ), .Y(n665) );
  INVX2 U309 ( .A(\memory[25][3] ), .Y(n657) );
  INVX2 U310 ( .A(\memory[26][3] ), .Y(n649) );
  INVX2 U311 ( .A(\memory[27][3] ), .Y(n641) );
  INVX2 U312 ( .A(\memory[3][3] ), .Y(n696) );
  INVX2 U313 ( .A(\memory[2][3] ), .Y(n688) );
  INVX2 U314 ( .A(\memory[1][3] ), .Y(n680) );
  INVX2 U315 ( .A(\memory[0][3] ), .Y(n672) );
  INVX2 U316 ( .A(\memory[8][3] ), .Y(n707) );
  INVX2 U317 ( .A(\memory[9][3] ), .Y(n715) );
  INVX2 U318 ( .A(\memory[10][3] ), .Y(n723) );
  INVX2 U319 ( .A(\memory[11][3] ), .Y(n731) );
  INVX2 U320 ( .A(\memory[16][2] ), .Y(n740) );
  INVX2 U321 ( .A(\memory[17][2] ), .Y(n748) );
  INVX2 U322 ( .A(\memory[18][2] ), .Y(n756) );
  INVX2 U323 ( .A(\memory[19][2] ), .Y(n764) );
  INVX2 U324 ( .A(\memory[24][2] ), .Y(n666) );
  INVX2 U325 ( .A(\memory[25][2] ), .Y(n658) );
  INVX2 U326 ( .A(\memory[26][2] ), .Y(n650) );
  INVX2 U327 ( .A(\memory[27][2] ), .Y(n642) );
  INVX2 U328 ( .A(\memory[3][2] ), .Y(n695) );
  INVX2 U329 ( .A(\memory[2][2] ), .Y(n687) );
  INVX2 U330 ( .A(\memory[1][2] ), .Y(n679) );
  INVX2 U331 ( .A(\memory[0][2] ), .Y(n671) );
  INVX2 U332 ( .A(\memory[8][2] ), .Y(n708) );
  INVX2 U333 ( .A(\memory[9][2] ), .Y(n716) );
  INVX2 U334 ( .A(\memory[10][2] ), .Y(n724) );
  INVX2 U335 ( .A(\memory[11][2] ), .Y(n732) );
  INVX2 U336 ( .A(\memory[16][1] ), .Y(n741) );
  INVX2 U337 ( .A(\memory[17][1] ), .Y(n749) );
  INVX2 U338 ( .A(\memory[18][1] ), .Y(n757) );
  INVX2 U339 ( .A(\memory[19][1] ), .Y(n765) );
  INVX2 U340 ( .A(\memory[24][1] ), .Y(n667) );
  INVX2 U341 ( .A(\memory[25][1] ), .Y(n659) );
  INVX2 U342 ( .A(\memory[26][1] ), .Y(n651) );
  INVX2 U343 ( .A(\memory[27][1] ), .Y(n643) );
  INVX2 U344 ( .A(\memory[3][1] ), .Y(n694) );
  INVX2 U345 ( .A(\memory[2][1] ), .Y(n686) );
  INVX2 U346 ( .A(\memory[1][1] ), .Y(n678) );
  INVX2 U347 ( .A(\memory[0][1] ), .Y(n670) );
  INVX2 U348 ( .A(\memory[8][1] ), .Y(n709) );
  INVX2 U349 ( .A(\memory[9][1] ), .Y(n717) );
  INVX2 U350 ( .A(\memory[10][1] ), .Y(n725) );
  INVX2 U351 ( .A(\memory[11][1] ), .Y(n733) );
  INVX2 U352 ( .A(\memory[16][0] ), .Y(n742) );
  INVX2 U353 ( .A(\memory[17][0] ), .Y(n750) );
  INVX2 U354 ( .A(\memory[18][0] ), .Y(n758) );
  INVX2 U355 ( .A(\memory[19][0] ), .Y(n766) );
  INVX2 U356 ( .A(\memory[24][0] ), .Y(n668) );
  INVX2 U357 ( .A(\memory[25][0] ), .Y(n660) );
  INVX2 U358 ( .A(\memory[26][0] ), .Y(n652) );
  INVX2 U359 ( .A(\memory[27][0] ), .Y(n644) );
  INVX2 U360 ( .A(\memory[3][0] ), .Y(n693) );
  INVX2 U361 ( .A(\memory[2][0] ), .Y(n685) );
  INVX2 U362 ( .A(\memory[1][0] ), .Y(n677) );
  INVX2 U363 ( .A(\memory[0][0] ), .Y(n669) );
  INVX2 U364 ( .A(\memory[8][0] ), .Y(n710) );
  INVX2 U365 ( .A(\memory[9][0] ), .Y(n718) );
  INVX2 U366 ( .A(\memory[10][0] ), .Y(n726) );
  INVX2 U367 ( .A(\memory[11][0] ), .Y(n734) );
  INVX2 U368 ( .A(\opcode[16][1] ), .Y(n775) );
  INVX2 U369 ( .A(\opcode[17][1] ), .Y(n777) );
  INVX2 U370 ( .A(\opcode[18][1] ), .Y(n779) );
  INVX2 U371 ( .A(\opcode[19][1] ), .Y(n781) );
  INVX2 U372 ( .A(\opcode[24][1] ), .Y(n627) );
  INVX2 U373 ( .A(\opcode[25][1] ), .Y(n625) );
  INVX2 U374 ( .A(\opcode[26][1] ), .Y(n623) );
  INVX2 U375 ( .A(\opcode[27][1] ), .Y(n621) );
  INVX2 U376 ( .A(\opcode[3][1] ), .Y(n636) );
  INVX2 U377 ( .A(\opcode[2][1] ), .Y(n634) );
  INVX2 U378 ( .A(\opcode[1][1] ), .Y(n632) );
  INVX2 U379 ( .A(\opcode[0][1] ), .Y(n630) );
  INVX2 U380 ( .A(\opcode[8][1] ), .Y(n767) );
  INVX2 U381 ( .A(\opcode[9][1] ), .Y(n769) );
  INVX2 U382 ( .A(\opcode[10][1] ), .Y(n771) );
  INVX2 U383 ( .A(\opcode[11][1] ), .Y(n773) );
  INVX2 U384 ( .A(\opcode[16][0] ), .Y(n776) );
  INVX2 U385 ( .A(\opcode[17][0] ), .Y(n778) );
  INVX2 U386 ( .A(\opcode[18][0] ), .Y(n780) );
  INVX2 U387 ( .A(\opcode[19][0] ), .Y(n782) );
  INVX2 U388 ( .A(n136), .Y(n619) );
  INVX2 U389 ( .A(\opcode[24][0] ), .Y(n628) );
  INVX2 U390 ( .A(\opcode[25][0] ), .Y(n626) );
  INVX2 U391 ( .A(\opcode[26][0] ), .Y(n624) );
  INVX2 U392 ( .A(\opcode[27][0] ), .Y(n622) );
  INVX2 U393 ( .A(\opcode[3][0] ), .Y(n635) );
  INVX2 U394 ( .A(\opcode[2][0] ), .Y(n633) );
  INVX2 U395 ( .A(\opcode[1][0] ), .Y(n631) );
  INVX2 U396 ( .A(\opcode[0][0] ), .Y(n629) );
  INVX2 U397 ( .A(\opcode[8][0] ), .Y(n768) );
  INVX2 U398 ( .A(\opcode[9][0] ), .Y(n770) );
  INVX2 U399 ( .A(\opcode[10][0] ), .Y(n772) );
  INVX2 U400 ( .A(\opcode[11][0] ), .Y(n774) );
  NAND2X1 U401 ( .A(readptr[0]), .B(n219), .Y(n545) );
  NAND2X1 U402 ( .A(n134), .B(n617), .Y(n164) );
  XNOR2X1 U403 ( .A(n70), .B(n43), .Y(n548) );
  XNOR2X1 U404 ( .A(n101), .B(n136), .Y(n553) );
  XNOR2X1 U405 ( .A(writeptr[4]), .B(readptr[4]), .Y(n558) );
  AND2X2 U406 ( .A(n553), .B(n558), .Y(n165) );
  NAND3X1 U407 ( .A(n166), .B(n548), .C(n165), .Y(n167) );
  MUX2X1 U408 ( .B(n167), .A(n702), .S(RST), .Y(n1432) );
  INVX2 U409 ( .A(OUT_OPCODE[0]), .Y(n170) );
  INVX2 U410 ( .A(n1226), .Y(n169) );
  NAND2X1 U411 ( .A(R_ENABLE), .B(n167), .Y(n614) );
  NAND2X1 U412 ( .A(n163), .B(state), .Y(n168) );
  MUX2X1 U413 ( .B(n170), .A(n169), .S(n113), .Y(n1562) );
  INVX2 U414 ( .A(OUT_OPCODE[1]), .Y(n172) );
  INVX2 U415 ( .A(n1199), .Y(n171) );
  MUX2X1 U416 ( .B(n172), .A(n171), .S(n114), .Y(n1561) );
  INVX2 U417 ( .A(DATA[0]), .Y(n174) );
  INVX2 U418 ( .A(n1172), .Y(n173) );
  MUX2X1 U419 ( .B(n174), .A(n173), .S(n113), .Y(n1560) );
  INVX2 U420 ( .A(DATA[1]), .Y(n176) );
  INVX2 U421 ( .A(n1015), .Y(n175) );
  MUX2X1 U422 ( .B(n176), .A(n175), .S(n114), .Y(n1559) );
  INVX2 U423 ( .A(DATA[2]), .Y(n178) );
  INVX2 U424 ( .A(n988), .Y(n177) );
  MUX2X1 U425 ( .B(n178), .A(n177), .S(n113), .Y(n1558) );
  INVX2 U426 ( .A(DATA[3]), .Y(n180) );
  INVX2 U427 ( .A(n961), .Y(n179) );
  MUX2X1 U428 ( .B(n180), .A(n179), .S(n114), .Y(n1557) );
  INVX2 U429 ( .A(DATA[4]), .Y(n182) );
  INVX2 U430 ( .A(n934), .Y(n181) );
  MUX2X1 U431 ( .B(n182), .A(n181), .S(n113), .Y(n1556) );
  INVX2 U432 ( .A(DATA[5]), .Y(n184) );
  INVX2 U433 ( .A(n863), .Y(n183) );
  MUX2X1 U434 ( .B(n184), .A(n183), .S(n114), .Y(n1555) );
  INVX2 U435 ( .A(DATA[6]), .Y(n186) );
  INVX2 U436 ( .A(n822), .Y(n185) );
  MUX2X1 U437 ( .B(n186), .A(n185), .S(n113), .Y(n1554) );
  INVX2 U438 ( .A(DATA[7]), .Y(n188) );
  INVX2 U439 ( .A(n783), .Y(n187) );
  MUX2X1 U440 ( .B(n188), .A(n187), .S(n114), .Y(n1553) );
  INVX2 U441 ( .A(RCV_OPCODE[0]), .Y(n339) );
  INVX2 U442 ( .A(\opcode[31][0] ), .Y(n195) );
  INVX2 U443 ( .A(n130), .Y(n203) );
  NAND3X1 U444 ( .A(n134), .B(n218), .C(n203), .Y(n328) );
  NAND3X1 U445 ( .A(n134), .B(n218), .C(n131), .Y(n331) );
  NAND2X1 U446 ( .A(n70), .B(n28), .Y(n189) );
  NAND2X1 U447 ( .A(n331), .B(n189), .Y(n569) );
  NAND3X1 U448 ( .A(n70), .B(n134), .C(n130), .Y(n586) );
  INVX2 U449 ( .A(n562), .Y(n190) );
  NOR2X1 U450 ( .A(n41), .B(n190), .Y(n192) );
  INVX2 U451 ( .A(n49), .Y(n611) );
  XNOR2X1 U452 ( .A(n575), .B(n611), .Y(n565) );
  NAND3X1 U453 ( .A(n100), .B(n63), .C(n70), .Y(n592) );
  AND2X2 U454 ( .A(n565), .B(n563), .Y(n191) );
  NAND3X1 U455 ( .A(n192), .B(n64), .C(n191), .Y(n299) );
  NAND3X1 U456 ( .A(n72), .B(n67), .C(n84), .Y(n336) );
  NAND2X1 U457 ( .A(n100), .B(n163), .Y(n286) );
  INVX2 U458 ( .A(n286), .Y(n264) );
  NAND3X1 U459 ( .A(n89), .B(W_ENABLE), .C(n299), .Y(n226) );
  NOR2X1 U460 ( .A(n31), .B(n59), .Y(n193) );
  NAND2X1 U461 ( .A(RCV_OPCODE[1]), .B(RCV_OPCODE[0]), .Y(n568) );
  NAND2X1 U462 ( .A(n193), .B(n160), .Y(n342) );
  OAI21X1 U463 ( .A(n328), .B(n95), .C(n342), .Y(n194) );
  INVX2 U464 ( .A(n194), .Y(n196) );
  MUX2X1 U465 ( .B(n137), .A(n195), .S(n196), .Y(n1552) );
  INVX2 U466 ( .A(\opcode[31][1] ), .Y(n197) );
  MUX2X1 U467 ( .B(n140), .A(n197), .S(n196), .Y(n1551) );
  INVX2 U468 ( .A(\opcode[30][0] ), .Y(n200) );
  OR2X2 U469 ( .A(n130), .B(n134), .Y(n577) );
  INVX2 U470 ( .A(n577), .Y(n209) );
  NAND3X1 U471 ( .A(n70), .B(n130), .C(n219), .Y(n316) );
  NOR2X1 U472 ( .A(n316), .B(n59), .Y(n198) );
  NAND2X1 U473 ( .A(n161), .B(n198), .Y(n352) );
  OAI21X1 U474 ( .A(n118), .B(n96), .C(n352), .Y(n199) );
  INVX2 U475 ( .A(n199), .Y(n201) );
  MUX2X1 U476 ( .B(n138), .A(n200), .S(n201), .Y(n1550) );
  INVX2 U477 ( .A(\opcode[30][1] ), .Y(n202) );
  MUX2X1 U478 ( .B(n142), .A(n202), .S(n201), .Y(n1549) );
  INVX2 U479 ( .A(\opcode[29][0] ), .Y(n206) );
  NAND3X1 U480 ( .A(n72), .B(n67), .C(n89), .Y(n236) );
  NAND3X1 U481 ( .A(n70), .B(n134), .C(n203), .Y(n321) );
  NOR2X1 U482 ( .A(n321), .B(n59), .Y(n204) );
  NAND2X1 U483 ( .A(n1), .B(n204), .Y(n362) );
  OAI21X1 U484 ( .A(n31), .B(n94), .C(n362), .Y(n205) );
  INVX2 U485 ( .A(n205), .Y(n207) );
  MUX2X1 U486 ( .B(n339), .A(n206), .S(n207), .Y(n1548) );
  INVX2 U487 ( .A(\opcode[29][1] ), .Y(n208) );
  MUX2X1 U488 ( .B(n142), .A(n208), .S(n207), .Y(n1547) );
  INVX2 U489 ( .A(\opcode[28][0] ), .Y(n212) );
  NAND2X1 U490 ( .A(n209), .B(n70), .Y(n325) );
  NOR2X1 U491 ( .A(n325), .B(n59), .Y(n210) );
  NAND2X1 U492 ( .A(n161), .B(n210), .Y(n372) );
  OAI21X1 U493 ( .A(n316), .B(n94), .C(n372), .Y(n211) );
  INVX2 U494 ( .A(n211), .Y(n213) );
  MUX2X1 U495 ( .B(n339), .A(n212), .S(n213), .Y(n1546) );
  INVX2 U496 ( .A(\opcode[28][1] ), .Y(n214) );
  MUX2X1 U497 ( .B(n142), .A(n214), .S(n213), .Y(n1545) );
  NOR2X1 U498 ( .A(n116), .B(n59), .Y(n215) );
  NAND2X1 U499 ( .A(n215), .B(n2), .Y(n382) );
  OAI21X1 U500 ( .A(n321), .B(n93), .C(n382), .Y(n216) );
  INVX2 U501 ( .A(n216), .Y(n217) );
  MUX2X1 U502 ( .B(n339), .A(n622), .S(n217), .Y(n1272) );
  MUX2X1 U503 ( .B(n142), .A(n621), .S(n217), .Y(n1271) );
  NAND3X1 U504 ( .A(n131), .B(n219), .C(n218), .Y(n337) );
  NOR2X1 U505 ( .A(n337), .B(n59), .Y(n220) );
  NAND2X1 U506 ( .A(n160), .B(n220), .Y(n384) );
  OAI21X1 U507 ( .A(n325), .B(n93), .C(n384), .Y(n221) );
  INVX2 U508 ( .A(n221), .Y(n222) );
  MUX2X1 U509 ( .B(n339), .A(n624), .S(n222), .Y(n1274) );
  MUX2X1 U510 ( .B(n142), .A(n623), .S(n222), .Y(n1273) );
  NOR2X1 U511 ( .A(n328), .B(n59), .Y(n223) );
  NAND2X1 U512 ( .A(n223), .B(n160), .Y(n386) );
  OAI21X1 U513 ( .A(n116), .B(n94), .C(n386), .Y(n224) );
  INVX2 U514 ( .A(n224), .Y(n225) );
  MUX2X1 U515 ( .B(n339), .A(n626), .S(n225), .Y(n1276) );
  MUX2X1 U516 ( .B(n142), .A(n625), .S(n225), .Y(n1275) );
  NOR2X1 U517 ( .A(n118), .B(n59), .Y(n227) );
  NAND2X1 U518 ( .A(n227), .B(n160), .Y(n388) );
  OAI21X1 U519 ( .A(n337), .B(n94), .C(n388), .Y(n228) );
  INVX2 U520 ( .A(n228), .Y(n229) );
  MUX2X1 U521 ( .B(n339), .A(n628), .S(n229), .Y(n1278) );
  MUX2X1 U522 ( .B(n142), .A(n627), .S(n229), .Y(n1277) );
  INVX2 U523 ( .A(\opcode[23][0] ), .Y(n232) );
  NAND3X1 U524 ( .A(n90), .B(W_ENABLE), .C(n299), .Y(n260) );
  NOR2X1 U525 ( .A(n31), .B(n61), .Y(n230) );
  NAND2X1 U526 ( .A(n2), .B(n230), .Y(n390) );
  OAI21X1 U527 ( .A(n328), .B(n93), .C(n4), .Y(n231) );
  INVX2 U528 ( .A(n231), .Y(n233) );
  MUX2X1 U529 ( .B(n138), .A(n232), .S(n233), .Y(n1280) );
  INVX2 U530 ( .A(\opcode[23][1] ), .Y(n234) );
  MUX2X1 U531 ( .B(n141), .A(n234), .S(n233), .Y(n1279) );
  INVX2 U532 ( .A(\opcode[22][0] ), .Y(n238) );
  NOR2X1 U533 ( .A(n316), .B(n61), .Y(n235) );
  NAND2X1 U534 ( .A(n160), .B(n235), .Y(n400) );
  OAI21X1 U535 ( .A(n118), .B(n94), .C(n400), .Y(n237) );
  INVX2 U536 ( .A(n237), .Y(n239) );
  MUX2X1 U537 ( .B(n138), .A(n238), .S(n239), .Y(n1282) );
  INVX2 U538 ( .A(\opcode[22][1] ), .Y(n240) );
  MUX2X1 U539 ( .B(n141), .A(n240), .S(n239), .Y(n1281) );
  INVX2 U540 ( .A(\opcode[21][0] ), .Y(n243) );
  NAND3X1 U541 ( .A(n72), .B(n67), .C(n90), .Y(n271) );
  NOR2X1 U542 ( .A(n321), .B(n61), .Y(n241) );
  NAND2X1 U543 ( .A(n161), .B(n241), .Y(n410) );
  OAI21X1 U544 ( .A(n31), .B(n97), .C(n5), .Y(n242) );
  INVX2 U545 ( .A(n242), .Y(n244) );
  MUX2X1 U546 ( .B(n138), .A(n243), .S(n244), .Y(n1284) );
  INVX2 U547 ( .A(\opcode[21][1] ), .Y(n245) );
  MUX2X1 U548 ( .B(n141), .A(n245), .S(n244), .Y(n1283) );
  INVX2 U549 ( .A(\opcode[20][0] ), .Y(n248) );
  NOR2X1 U550 ( .A(n325), .B(n61), .Y(n246) );
  NAND2X1 U551 ( .A(n160), .B(n246), .Y(n420) );
  OAI21X1 U552 ( .A(n316), .B(n97), .C(n420), .Y(n247) );
  MUX2X1 U553 ( .B(n138), .A(n248), .S(n249), .Y(n1286) );
  INVX2 U554 ( .A(\opcode[20][1] ), .Y(n250) );
  MUX2X1 U555 ( .B(n141), .A(n250), .S(n249), .Y(n1285) );
  NOR2X1 U556 ( .A(n116), .B(n61), .Y(n251) );
  NAND2X1 U557 ( .A(n251), .B(n161), .Y(n430) );
  OAI21X1 U558 ( .A(n321), .B(n97), .C(n430), .Y(n252) );
  INVX2 U559 ( .A(n252), .Y(n253) );
  MUX2X1 U560 ( .B(n138), .A(n782), .S(n253), .Y(n1544) );
  MUX2X1 U561 ( .B(n141), .A(n781), .S(n253), .Y(n1543) );
  NOR2X1 U562 ( .A(n337), .B(n61), .Y(n254) );
  NAND2X1 U563 ( .A(n160), .B(n254), .Y(n432) );
  OAI21X1 U564 ( .A(n325), .B(n98), .C(n432), .Y(n255) );
  INVX2 U565 ( .A(n255), .Y(n256) );
  MUX2X1 U566 ( .B(n138), .A(n780), .S(n256), .Y(n1542) );
  MUX2X1 U567 ( .B(n141), .A(n779), .S(n256), .Y(n1541) );
  NOR2X1 U568 ( .A(n328), .B(n61), .Y(n257) );
  NAND2X1 U569 ( .A(n161), .B(n257), .Y(n434) );
  OAI21X1 U570 ( .A(n116), .B(n98), .C(n434), .Y(n258) );
  INVX2 U571 ( .A(n258), .Y(n259) );
  MUX2X1 U572 ( .B(n138), .A(n778), .S(n259), .Y(n1540) );
  MUX2X1 U573 ( .B(n141), .A(n777), .S(n259), .Y(n1539) );
  NOR2X1 U574 ( .A(n118), .B(n61), .Y(n261) );
  NAND2X1 U575 ( .A(n261), .B(n160), .Y(n436) );
  OAI21X1 U576 ( .A(n337), .B(n98), .C(n436), .Y(n262) );
  INVX2 U577 ( .A(n262), .Y(n263) );
  MUX2X1 U578 ( .B(n138), .A(n776), .S(n263), .Y(n1538) );
  MUX2X1 U579 ( .B(n141), .A(n775), .S(n263), .Y(n1537) );
  INVX2 U580 ( .A(\opcode[15][0] ), .Y(n267) );
  NOR2X1 U581 ( .A(n31), .B(n478), .Y(n265) );
  NAND2X1 U582 ( .A(n161), .B(n265), .Y(n438) );
  OAI21X1 U583 ( .A(n328), .B(n98), .C(n438), .Y(n266) );
  MUX2X1 U584 ( .B(n138), .A(n267), .S(n268), .Y(n1288) );
  INVX2 U585 ( .A(\opcode[15][1] ), .Y(n269) );
  MUX2X1 U586 ( .B(n141), .A(n269), .S(n268), .Y(n1287) );
  INVX2 U587 ( .A(\opcode[14][0] ), .Y(n273) );
  NOR2X1 U588 ( .A(n68), .B(n69), .Y(n270) );
  NAND2X1 U589 ( .A(n270), .B(n161), .Y(n448) );
  OAI21X1 U590 ( .A(n118), .B(n98), .C(n448), .Y(n272) );
  INVX2 U591 ( .A(n272), .Y(n274) );
  MUX2X1 U592 ( .B(n138), .A(n273), .S(n274), .Y(n1290) );
  INVX2 U593 ( .A(\opcode[14][1] ), .Y(n275) );
  MUX2X1 U594 ( .B(n141), .A(n275), .S(n274), .Y(n1289) );
  INVX2 U595 ( .A(\opcode[13][0] ), .Y(n278) );
  NAND3X1 U596 ( .A(n72), .B(n67), .C(n83), .Y(n305) );
  NOR2X1 U597 ( .A(n321), .B(n47), .Y(n276) );
  NAND2X1 U598 ( .A(n276), .B(n161), .Y(n458) );
  OAI21X1 U599 ( .A(n31), .B(n92), .C(n458), .Y(n277) );
  INVX2 U600 ( .A(n277), .Y(n279) );
  MUX2X1 U601 ( .B(n138), .A(n278), .S(n279), .Y(n1292) );
  INVX2 U602 ( .A(\opcode[13][1] ), .Y(n280) );
  MUX2X1 U603 ( .B(n141), .A(n280), .S(n279), .Y(n1291) );
  INVX2 U604 ( .A(\opcode[12][0] ), .Y(n283) );
  NOR2X1 U605 ( .A(n325), .B(n47), .Y(n281) );
  NAND2X1 U606 ( .A(n281), .B(n161), .Y(n468) );
  OAI21X1 U607 ( .A(n316), .B(n91), .C(n468), .Y(n282) );
  INVX2 U608 ( .A(n282), .Y(n284) );
  MUX2X1 U609 ( .B(n137), .A(n283), .S(n284), .Y(n1294) );
  INVX2 U610 ( .A(\opcode[12][1] ), .Y(n285) );
  MUX2X1 U611 ( .B(n140), .A(n285), .S(n284), .Y(n1293) );
  NOR3X1 U612 ( .A(n52), .B(n579), .C(n286), .Y(n288) );
  AND2X2 U613 ( .A(n288), .B(n287), .Y(n289) );
  MUX2X1 U614 ( .B(n774), .A(n137), .S(n289), .Y(n1536) );
  MUX2X1 U615 ( .B(n773), .A(n142), .S(n289), .Y(n1535) );
  NOR2X1 U616 ( .A(n337), .B(n478), .Y(n290) );
  NAND2X1 U617 ( .A(n290), .B(n161), .Y(n482) );
  OAI21X1 U618 ( .A(n325), .B(n92), .C(n482), .Y(n291) );
  INVX2 U619 ( .A(n291), .Y(n292) );
  MUX2X1 U620 ( .B(n137), .A(n772), .S(n292), .Y(n1534) );
  MUX2X1 U621 ( .B(n140), .A(n771), .S(n292), .Y(n1533) );
  NOR2X1 U622 ( .A(n328), .B(n47), .Y(n293) );
  NAND2X1 U623 ( .A(n293), .B(n160), .Y(n484) );
  OAI21X1 U624 ( .A(n116), .B(n92), .C(n484), .Y(n294) );
  INVX2 U625 ( .A(n294), .Y(n295) );
  MUX2X1 U626 ( .B(n137), .A(n770), .S(n295), .Y(n1532) );
  MUX2X1 U627 ( .B(n140), .A(n769), .S(n295), .Y(n1531) );
  NOR2X1 U628 ( .A(n478), .B(n118), .Y(n296) );
  NAND2X1 U629 ( .A(n161), .B(n296), .Y(n486) );
  OAI21X1 U630 ( .A(n337), .B(n91), .C(n486), .Y(n297) );
  MUX2X1 U631 ( .B(n137), .A(n768), .S(n298), .Y(n1530) );
  MUX2X1 U632 ( .B(n140), .A(n767), .S(n298), .Y(n1529) );
  INVX2 U633 ( .A(\opcode[7][0] ), .Y(n301) );
  NAND3X1 U634 ( .A(n84), .B(n24), .C(W_ENABLE), .Y(n334) );
  INVX2 U635 ( .A(n334), .Y(n329) );
  NAND3X1 U636 ( .A(n117), .B(n329), .C(n2), .Y(n488) );
  OAI21X1 U637 ( .A(n328), .B(n91), .C(n488), .Y(n300) );
  INVX2 U638 ( .A(n300), .Y(n302) );
  MUX2X1 U639 ( .B(n137), .A(n301), .S(n302), .Y(n1563) );
  INVX2 U640 ( .A(\opcode[7][1] ), .Y(n303) );
  MUX2X1 U641 ( .B(n140), .A(n303), .S(n302), .Y(n1564) );
  INVX2 U642 ( .A(\opcode[6][0] ), .Y(n307) );
  INVX2 U643 ( .A(n316), .Y(n304) );
  NAND3X1 U644 ( .A(n304), .B(n329), .C(n2), .Y(n498) );
  OAI21X1 U645 ( .A(n118), .B(n92), .C(n498), .Y(n306) );
  INVX2 U646 ( .A(n306), .Y(n308) );
  MUX2X1 U647 ( .B(n137), .A(n307), .S(n308), .Y(n1573) );
  INVX2 U648 ( .A(\opcode[6][1] ), .Y(n309) );
  MUX2X1 U649 ( .B(n140), .A(n309), .S(n308), .Y(n1574) );
  INVX2 U650 ( .A(\opcode[5][0] ), .Y(n312) );
  INVX2 U651 ( .A(n321), .Y(n310) );
  NAND3X1 U652 ( .A(n310), .B(n329), .C(n2), .Y(n508) );
  OAI21X1 U653 ( .A(n31), .B(n95), .C(n508), .Y(n311) );
  INVX2 U654 ( .A(n311), .Y(n313) );
  MUX2X1 U655 ( .B(n137), .A(n312), .S(n313), .Y(n1583) );
  INVX2 U656 ( .A(\opcode[5][1] ), .Y(n314) );
  MUX2X1 U657 ( .B(n140), .A(n314), .S(n313), .Y(n1584) );
  INVX2 U658 ( .A(\opcode[4][0] ), .Y(n318) );
  INVX2 U659 ( .A(n325), .Y(n315) );
  NAND3X1 U660 ( .A(n315), .B(n329), .C(n2), .Y(n518) );
  OAI21X1 U661 ( .A(n316), .B(n95), .C(n518), .Y(n317) );
  INVX2 U662 ( .A(n317), .Y(n319) );
  MUX2X1 U663 ( .B(n137), .A(n318), .S(n319), .Y(n1593) );
  INVX2 U664 ( .A(\opcode[4][1] ), .Y(n320) );
  MUX2X1 U665 ( .B(n140), .A(n320), .S(n319), .Y(n1594) );
  NAND3X1 U666 ( .A(n115), .B(n329), .C(n2), .Y(n528) );
  OAI21X1 U667 ( .A(n321), .B(n96), .C(n528), .Y(n322) );
  MUX2X1 U668 ( .B(n137), .A(n635), .S(n323), .Y(n1301) );
  MUX2X1 U669 ( .B(n140), .A(n636), .S(n323), .Y(n1302) );
  INVX2 U670 ( .A(n337), .Y(n324) );
  NAND3X1 U671 ( .A(n324), .B(n329), .C(n2), .Y(n530) );
  OAI21X1 U672 ( .A(n325), .B(n96), .C(n530), .Y(n326) );
  INVX2 U673 ( .A(n326), .Y(n327) );
  MUX2X1 U674 ( .B(n137), .A(n633), .S(n327), .Y(n1299) );
  MUX2X1 U675 ( .B(n140), .A(n634), .S(n327), .Y(n1300) );
  INVX2 U676 ( .A(n328), .Y(n330) );
  NAND3X1 U677 ( .A(n330), .B(n329), .C(n160), .Y(n532) );
  OAI21X1 U678 ( .A(n116), .B(n96), .C(n532), .Y(n332) );
  INVX2 U679 ( .A(n332), .Y(n333) );
  MUX2X1 U680 ( .B(n137), .A(n631), .S(n333), .Y(n1297) );
  MUX2X1 U681 ( .B(n140), .A(n632), .S(n333), .Y(n1298) );
  NOR2X1 U682 ( .A(n118), .B(n334), .Y(n335) );
  NAND2X1 U683 ( .A(n335), .B(n2), .Y(n534) );
  OAI21X1 U684 ( .A(n337), .B(n96), .C(n534), .Y(n338) );
  INVX2 U685 ( .A(n338), .Y(n340) );
  MUX2X1 U686 ( .B(n138), .A(n629), .S(n340), .Y(n1295) );
  MUX2X1 U687 ( .B(n141), .A(n630), .S(n340), .Y(n1296) );
  INVX2 U688 ( .A(\memory[31][0] ), .Y(n343) );
  MUX2X1 U689 ( .B(n343), .A(n144), .S(n350), .Y(n1528) );
  INVX2 U690 ( .A(\memory[31][1] ), .Y(n344) );
  MUX2X1 U691 ( .B(n344), .A(n146), .S(n350), .Y(n1527) );
  INVX2 U692 ( .A(\memory[31][2] ), .Y(n345) );
  MUX2X1 U693 ( .B(n345), .A(n148), .S(n350), .Y(n1526) );
  INVX2 U694 ( .A(\memory[31][3] ), .Y(n346) );
  MUX2X1 U695 ( .B(n346), .A(n150), .S(n350), .Y(n1525) );
  INVX2 U696 ( .A(\memory[31][4] ), .Y(n347) );
  MUX2X1 U697 ( .B(n347), .A(n152), .S(n350), .Y(n1524) );
  INVX2 U698 ( .A(\memory[31][5] ), .Y(n348) );
  MUX2X1 U699 ( .B(n348), .A(n154), .S(n350), .Y(n1523) );
  INVX2 U700 ( .A(\memory[31][6] ), .Y(n349) );
  MUX2X1 U701 ( .B(n349), .A(n156), .S(n350), .Y(n1522) );
  INVX2 U702 ( .A(\memory[31][7] ), .Y(n351) );
  MUX2X1 U703 ( .B(n351), .A(n158), .S(n350), .Y(n1521) );
  INVX2 U704 ( .A(\memory[30][0] ), .Y(n353) );
  MUX2X1 U705 ( .B(n353), .A(n144), .S(n360), .Y(n1520) );
  INVX2 U706 ( .A(\memory[30][1] ), .Y(n354) );
  MUX2X1 U707 ( .B(n354), .A(n146), .S(n360), .Y(n1519) );
  INVX2 U708 ( .A(\memory[30][2] ), .Y(n355) );
  MUX2X1 U709 ( .B(n355), .A(n148), .S(n360), .Y(n1518) );
  INVX2 U710 ( .A(\memory[30][3] ), .Y(n356) );
  MUX2X1 U711 ( .B(n356), .A(n150), .S(n360), .Y(n1517) );
  INVX2 U712 ( .A(\memory[30][4] ), .Y(n357) );
  MUX2X1 U713 ( .B(n357), .A(n152), .S(n360), .Y(n1516) );
  INVX2 U714 ( .A(\memory[30][5] ), .Y(n358) );
  MUX2X1 U715 ( .B(n358), .A(n154), .S(n360), .Y(n1515) );
  INVX2 U716 ( .A(\memory[30][6] ), .Y(n359) );
  MUX2X1 U717 ( .B(n359), .A(n156), .S(n360), .Y(n1514) );
  INVX2 U718 ( .A(\memory[30][7] ), .Y(n361) );
  MUX2X1 U719 ( .B(n361), .A(n158), .S(n360), .Y(n1513) );
  INVX2 U720 ( .A(\memory[29][0] ), .Y(n363) );
  MUX2X1 U721 ( .B(n363), .A(n144), .S(n370), .Y(n1512) );
  INVX2 U722 ( .A(\memory[29][1] ), .Y(n364) );
  MUX2X1 U723 ( .B(n364), .A(n146), .S(n370), .Y(n1511) );
  INVX2 U724 ( .A(\memory[29][2] ), .Y(n365) );
  MUX2X1 U725 ( .B(n365), .A(n148), .S(n370), .Y(n1510) );
  INVX2 U726 ( .A(\memory[29][3] ), .Y(n366) );
  MUX2X1 U727 ( .B(n366), .A(n150), .S(n370), .Y(n1509) );
  INVX2 U728 ( .A(\memory[29][4] ), .Y(n367) );
  MUX2X1 U729 ( .B(n367), .A(n152), .S(n370), .Y(n1508) );
  INVX2 U730 ( .A(\memory[29][5] ), .Y(n368) );
  MUX2X1 U731 ( .B(n368), .A(n154), .S(n370), .Y(n1507) );
  INVX2 U732 ( .A(\memory[29][6] ), .Y(n369) );
  MUX2X1 U733 ( .B(n369), .A(n156), .S(n370), .Y(n1506) );
  INVX2 U734 ( .A(\memory[29][7] ), .Y(n371) );
  MUX2X1 U735 ( .B(n371), .A(n158), .S(n370), .Y(n1505) );
  INVX2 U736 ( .A(\memory[28][0] ), .Y(n373) );
  MUX2X1 U737 ( .B(n373), .A(n144), .S(n380), .Y(n1504) );
  INVX2 U738 ( .A(\memory[28][1] ), .Y(n374) );
  MUX2X1 U739 ( .B(n374), .A(n146), .S(n380), .Y(n1503) );
  INVX2 U740 ( .A(\memory[28][2] ), .Y(n375) );
  MUX2X1 U741 ( .B(n375), .A(n148), .S(n380), .Y(n1502) );
  INVX2 U742 ( .A(\memory[28][3] ), .Y(n376) );
  MUX2X1 U743 ( .B(n376), .A(n150), .S(n380), .Y(n1501) );
  INVX2 U744 ( .A(\memory[28][4] ), .Y(n377) );
  MUX2X1 U745 ( .B(n377), .A(n152), .S(n380), .Y(n1500) );
  INVX2 U746 ( .A(\memory[28][5] ), .Y(n378) );
  MUX2X1 U747 ( .B(n378), .A(n154), .S(n380), .Y(n1499) );
  INVX2 U748 ( .A(\memory[28][6] ), .Y(n379) );
  MUX2X1 U749 ( .B(n379), .A(n156), .S(n380), .Y(n1498) );
  INVX2 U750 ( .A(\memory[28][7] ), .Y(n381) );
  MUX2X1 U751 ( .B(n381), .A(n158), .S(n380), .Y(n1497) );
  MUX2X1 U752 ( .B(n644), .A(n144), .S(n383), .Y(n1310) );
  MUX2X1 U753 ( .B(n643), .A(n146), .S(n383), .Y(n1309) );
  MUX2X1 U754 ( .B(n642), .A(n148), .S(n383), .Y(n1308) );
  MUX2X1 U755 ( .B(n641), .A(n150), .S(n383), .Y(n1307) );
  MUX2X1 U756 ( .B(n640), .A(n152), .S(n383), .Y(n1306) );
  MUX2X1 U757 ( .B(n639), .A(n154), .S(n383), .Y(n1305) );
  MUX2X1 U758 ( .B(n638), .A(n156), .S(n383), .Y(n1304) );
  MUX2X1 U759 ( .B(n637), .A(n158), .S(n383), .Y(n1303) );
  MUX2X1 U760 ( .B(n652), .A(n144), .S(n385), .Y(n1318) );
  MUX2X1 U761 ( .B(n651), .A(n146), .S(n385), .Y(n1317) );
  MUX2X1 U762 ( .B(n650), .A(n148), .S(n385), .Y(n1316) );
  MUX2X1 U763 ( .B(n649), .A(n150), .S(n385), .Y(n1315) );
  MUX2X1 U764 ( .B(n648), .A(n152), .S(n385), .Y(n1314) );
  MUX2X1 U765 ( .B(n647), .A(n154), .S(n385), .Y(n1313) );
  MUX2X1 U766 ( .B(n646), .A(n156), .S(n385), .Y(n1312) );
  MUX2X1 U767 ( .B(n645), .A(n158), .S(n385), .Y(n1311) );
  MUX2X1 U768 ( .B(n660), .A(n144), .S(n387), .Y(n1326) );
  MUX2X1 U769 ( .B(n659), .A(n146), .S(n387), .Y(n1325) );
  MUX2X1 U770 ( .B(n658), .A(n148), .S(n387), .Y(n1324) );
  MUX2X1 U771 ( .B(n657), .A(n150), .S(n387), .Y(n1323) );
  MUX2X1 U772 ( .B(n656), .A(n152), .S(n387), .Y(n1322) );
  MUX2X1 U773 ( .B(n655), .A(n154), .S(n387), .Y(n1321) );
  MUX2X1 U774 ( .B(n654), .A(n156), .S(n387), .Y(n1320) );
  MUX2X1 U775 ( .B(n653), .A(n158), .S(n387), .Y(n1319) );
  MUX2X1 U776 ( .B(n668), .A(n144), .S(n389), .Y(n1334) );
  MUX2X1 U777 ( .B(n667), .A(n146), .S(n389), .Y(n1333) );
  MUX2X1 U778 ( .B(n666), .A(n148), .S(n389), .Y(n1332) );
  MUX2X1 U779 ( .B(n665), .A(n150), .S(n389), .Y(n1331) );
  MUX2X1 U780 ( .B(n664), .A(n152), .S(n389), .Y(n1330) );
  MUX2X1 U781 ( .B(n663), .A(n540), .S(n389), .Y(n1329) );
  MUX2X1 U782 ( .B(n662), .A(n156), .S(n389), .Y(n1328) );
  MUX2X1 U783 ( .B(n661), .A(n158), .S(n389), .Y(n1327) );
  INVX2 U784 ( .A(\memory[23][0] ), .Y(n391) );
  MUX2X1 U785 ( .B(n391), .A(n144), .S(n398), .Y(n1342) );
  INVX2 U786 ( .A(\memory[23][1] ), .Y(n392) );
  MUX2X1 U787 ( .B(n392), .A(n146), .S(n398), .Y(n1341) );
  INVX2 U788 ( .A(\memory[23][2] ), .Y(n393) );
  MUX2X1 U789 ( .B(n393), .A(n148), .S(n398), .Y(n1340) );
  INVX2 U790 ( .A(\memory[23][3] ), .Y(n394) );
  MUX2X1 U791 ( .B(n394), .A(n150), .S(n398), .Y(n1339) );
  INVX2 U792 ( .A(\memory[23][4] ), .Y(n395) );
  MUX2X1 U793 ( .B(n395), .A(n152), .S(n398), .Y(n1338) );
  INVX2 U794 ( .A(\memory[23][5] ), .Y(n396) );
  MUX2X1 U795 ( .B(n396), .A(n540), .S(n398), .Y(n1337) );
  INVX2 U796 ( .A(\memory[23][6] ), .Y(n397) );
  MUX2X1 U797 ( .B(n397), .A(n156), .S(n398), .Y(n1336) );
  INVX2 U798 ( .A(\memory[23][7] ), .Y(n399) );
  MUX2X1 U799 ( .B(n399), .A(n158), .S(n398), .Y(n1335) );
  INVX2 U800 ( .A(\memory[22][0] ), .Y(n401) );
  MUX2X1 U801 ( .B(n401), .A(n144), .S(n408), .Y(n1350) );
  INVX2 U802 ( .A(\memory[22][1] ), .Y(n402) );
  MUX2X1 U803 ( .B(n402), .A(n146), .S(n408), .Y(n1349) );
  INVX2 U804 ( .A(\memory[22][2] ), .Y(n403) );
  MUX2X1 U805 ( .B(n403), .A(n148), .S(n408), .Y(n1348) );
  INVX2 U806 ( .A(\memory[22][3] ), .Y(n404) );
  MUX2X1 U807 ( .B(n404), .A(n150), .S(n408), .Y(n1347) );
  INVX2 U808 ( .A(\memory[22][4] ), .Y(n405) );
  MUX2X1 U809 ( .B(n405), .A(n152), .S(n408), .Y(n1346) );
  INVX2 U810 ( .A(\memory[22][5] ), .Y(n406) );
  MUX2X1 U811 ( .B(n406), .A(n540), .S(n408), .Y(n1345) );
  INVX2 U812 ( .A(\memory[22][6] ), .Y(n407) );
  MUX2X1 U813 ( .B(n407), .A(n156), .S(n408), .Y(n1344) );
  INVX2 U814 ( .A(\memory[22][7] ), .Y(n409) );
  MUX2X1 U815 ( .B(n409), .A(n158), .S(n408), .Y(n1343) );
  INVX2 U816 ( .A(\memory[21][0] ), .Y(n411) );
  MUX2X1 U817 ( .B(n411), .A(n144), .S(n418), .Y(n1358) );
  INVX2 U818 ( .A(\memory[21][1] ), .Y(n412) );
  MUX2X1 U819 ( .B(n412), .A(n146), .S(n418), .Y(n1357) );
  INVX2 U820 ( .A(\memory[21][2] ), .Y(n413) );
  MUX2X1 U821 ( .B(n413), .A(n148), .S(n418), .Y(n1356) );
  INVX2 U822 ( .A(\memory[21][3] ), .Y(n414) );
  MUX2X1 U823 ( .B(n414), .A(n150), .S(n418), .Y(n1355) );
  INVX2 U824 ( .A(\memory[21][4] ), .Y(n415) );
  MUX2X1 U825 ( .B(n415), .A(n152), .S(n418), .Y(n1354) );
  INVX2 U826 ( .A(\memory[21][5] ), .Y(n416) );
  MUX2X1 U827 ( .B(n416), .A(n540), .S(n418), .Y(n1353) );
  INVX2 U828 ( .A(\memory[21][6] ), .Y(n417) );
  MUX2X1 U829 ( .B(n417), .A(n156), .S(n418), .Y(n1352) );
  INVX2 U830 ( .A(\memory[21][7] ), .Y(n419) );
  MUX2X1 U831 ( .B(n419), .A(n158), .S(n418), .Y(n1351) );
  INVX2 U832 ( .A(\memory[20][0] ), .Y(n421) );
  MUX2X1 U833 ( .B(n421), .A(n144), .S(n428), .Y(n1366) );
  INVX2 U834 ( .A(\memory[20][1] ), .Y(n422) );
  MUX2X1 U835 ( .B(n422), .A(n146), .S(n428), .Y(n1365) );
  INVX2 U836 ( .A(\memory[20][2] ), .Y(n423) );
  MUX2X1 U837 ( .B(n423), .A(n148), .S(n428), .Y(n1364) );
  INVX2 U838 ( .A(\memory[20][3] ), .Y(n424) );
  MUX2X1 U839 ( .B(n424), .A(n150), .S(n428), .Y(n1363) );
  INVX2 U840 ( .A(\memory[20][4] ), .Y(n425) );
  MUX2X1 U841 ( .B(n425), .A(n152), .S(n428), .Y(n1362) );
  INVX2 U842 ( .A(\memory[20][5] ), .Y(n426) );
  MUX2X1 U843 ( .B(n426), .A(n154), .S(n428), .Y(n1361) );
  INVX2 U844 ( .A(\memory[20][6] ), .Y(n427) );
  MUX2X1 U845 ( .B(n427), .A(n156), .S(n428), .Y(n1360) );
  INVX2 U846 ( .A(\memory[20][7] ), .Y(n429) );
  MUX2X1 U847 ( .B(n429), .A(n158), .S(n428), .Y(n1359) );
  MUX2X1 U848 ( .B(n766), .A(n144), .S(n431), .Y(n1496) );
  MUX2X1 U849 ( .B(n765), .A(n146), .S(n431), .Y(n1495) );
  MUX2X1 U850 ( .B(n764), .A(n148), .S(n431), .Y(n1494) );
  MUX2X1 U851 ( .B(n763), .A(n150), .S(n431), .Y(n1493) );
  MUX2X1 U852 ( .B(n762), .A(n152), .S(n431), .Y(n1492) );
  MUX2X1 U853 ( .B(n761), .A(n540), .S(n431), .Y(n1491) );
  MUX2X1 U854 ( .B(n760), .A(n156), .S(n431), .Y(n1490) );
  MUX2X1 U855 ( .B(n759), .A(n159), .S(n431), .Y(n1489) );
  MUX2X1 U856 ( .B(n758), .A(n144), .S(n433), .Y(n1488) );
  MUX2X1 U857 ( .B(n757), .A(n146), .S(n433), .Y(n1487) );
  MUX2X1 U858 ( .B(n756), .A(n148), .S(n433), .Y(n1486) );
  MUX2X1 U859 ( .B(n755), .A(n150), .S(n433), .Y(n1485) );
  MUX2X1 U860 ( .B(n754), .A(n152), .S(n433), .Y(n1484) );
  MUX2X1 U861 ( .B(n753), .A(n540), .S(n433), .Y(n1483) );
  MUX2X1 U862 ( .B(n752), .A(n156), .S(n433), .Y(n1482) );
  MUX2X1 U863 ( .B(n751), .A(n159), .S(n433), .Y(n1481) );
  MUX2X1 U864 ( .B(n750), .A(n144), .S(n435), .Y(n1480) );
  MUX2X1 U865 ( .B(n749), .A(n146), .S(n435), .Y(n1479) );
  MUX2X1 U866 ( .B(n748), .A(n148), .S(n435), .Y(n1478) );
  MUX2X1 U867 ( .B(n747), .A(n150), .S(n435), .Y(n1477) );
  MUX2X1 U868 ( .B(n746), .A(n152), .S(n435), .Y(n1476) );
  MUX2X1 U869 ( .B(n745), .A(n540), .S(n435), .Y(n1475) );
  MUX2X1 U870 ( .B(n744), .A(n156), .S(n435), .Y(n1474) );
  MUX2X1 U871 ( .B(n743), .A(n159), .S(n435), .Y(n1473) );
  MUX2X1 U872 ( .B(n742), .A(n144), .S(n437), .Y(n1472) );
  MUX2X1 U873 ( .B(n741), .A(n146), .S(n437), .Y(n1471) );
  MUX2X1 U874 ( .B(n740), .A(n148), .S(n437), .Y(n1470) );
  MUX2X1 U875 ( .B(n739), .A(n150), .S(n437), .Y(n1469) );
  MUX2X1 U876 ( .B(n738), .A(n152), .S(n437), .Y(n1468) );
  MUX2X1 U877 ( .B(n737), .A(n540), .S(n437), .Y(n1467) );
  MUX2X1 U878 ( .B(n736), .A(n156), .S(n437), .Y(n1466) );
  MUX2X1 U879 ( .B(n735), .A(n159), .S(n437), .Y(n1465) );
  INVX2 U880 ( .A(\memory[15][0] ), .Y(n439) );
  MUX2X1 U881 ( .B(n439), .A(n144), .S(n446), .Y(n1374) );
  INVX2 U882 ( .A(\memory[15][1] ), .Y(n440) );
  MUX2X1 U883 ( .B(n440), .A(n146), .S(n446), .Y(n1373) );
  INVX2 U884 ( .A(\memory[15][2] ), .Y(n441) );
  MUX2X1 U885 ( .B(n441), .A(n148), .S(n446), .Y(n1372) );
  INVX2 U886 ( .A(\memory[15][3] ), .Y(n442) );
  MUX2X1 U887 ( .B(n442), .A(n150), .S(n446), .Y(n1371) );
  INVX2 U888 ( .A(\memory[15][4] ), .Y(n443) );
  MUX2X1 U889 ( .B(n443), .A(n152), .S(n446), .Y(n1370) );
  INVX2 U890 ( .A(\memory[15][5] ), .Y(n444) );
  MUX2X1 U891 ( .B(n444), .A(n540), .S(n446), .Y(n1369) );
  INVX2 U892 ( .A(\memory[15][6] ), .Y(n445) );
  MUX2X1 U893 ( .B(n445), .A(n156), .S(n446), .Y(n1368) );
  INVX2 U894 ( .A(\memory[15][7] ), .Y(n447) );
  MUX2X1 U895 ( .B(n447), .A(n159), .S(n446), .Y(n1367) );
  INVX2 U896 ( .A(\memory[14][0] ), .Y(n449) );
  MUX2X1 U897 ( .B(n449), .A(n144), .S(n456), .Y(n1382) );
  INVX2 U898 ( .A(\memory[14][1] ), .Y(n450) );
  MUX2X1 U899 ( .B(n450), .A(n536), .S(n456), .Y(n1381) );
  INVX2 U900 ( .A(\memory[14][2] ), .Y(n451) );
  MUX2X1 U901 ( .B(n451), .A(n148), .S(n456), .Y(n1380) );
  INVX2 U902 ( .A(\memory[14][3] ), .Y(n452) );
  MUX2X1 U903 ( .B(n452), .A(n150), .S(n456), .Y(n1379) );
  INVX2 U904 ( .A(\memory[14][4] ), .Y(n453) );
  MUX2X1 U905 ( .B(n453), .A(n152), .S(n456), .Y(n1378) );
  INVX2 U906 ( .A(\memory[14][5] ), .Y(n454) );
  MUX2X1 U907 ( .B(n454), .A(n540), .S(n456), .Y(n1377) );
  INVX2 U908 ( .A(\memory[14][6] ), .Y(n455) );
  MUX2X1 U909 ( .B(n455), .A(n541), .S(n456), .Y(n1376) );
  INVX2 U910 ( .A(\memory[14][7] ), .Y(n457) );
  MUX2X1 U911 ( .B(n457), .A(n159), .S(n456), .Y(n1375) );
  INVX2 U912 ( .A(\memory[13][0] ), .Y(n459) );
  MUX2X1 U913 ( .B(n459), .A(n144), .S(n466), .Y(n1390) );
  INVX2 U914 ( .A(\memory[13][1] ), .Y(n460) );
  MUX2X1 U915 ( .B(n460), .A(n536), .S(n466), .Y(n1389) );
  INVX2 U916 ( .A(\memory[13][2] ), .Y(n461) );
  MUX2X1 U917 ( .B(n461), .A(n148), .S(n466), .Y(n1388) );
  INVX2 U918 ( .A(\memory[13][3] ), .Y(n462) );
  MUX2X1 U919 ( .B(n462), .A(n150), .S(n466), .Y(n1387) );
  INVX2 U920 ( .A(\memory[13][4] ), .Y(n463) );
  MUX2X1 U921 ( .B(n463), .A(n152), .S(n466), .Y(n1386) );
  INVX2 U922 ( .A(\memory[13][5] ), .Y(n464) );
  MUX2X1 U923 ( .B(n464), .A(n540), .S(n466), .Y(n1385) );
  INVX2 U924 ( .A(\memory[13][6] ), .Y(n465) );
  MUX2X1 U925 ( .B(n465), .A(n541), .S(n466), .Y(n1384) );
  INVX2 U926 ( .A(\memory[13][7] ), .Y(n467) );
  MUX2X1 U927 ( .B(n467), .A(n159), .S(n466), .Y(n1383) );
  INVX2 U928 ( .A(\memory[12][0] ), .Y(n469) );
  MUX2X1 U929 ( .B(n469), .A(n535), .S(n476), .Y(n1398) );
  INVX2 U930 ( .A(\memory[12][1] ), .Y(n470) );
  MUX2X1 U931 ( .B(n470), .A(n536), .S(n476), .Y(n1397) );
  INVX2 U932 ( .A(\memory[12][2] ), .Y(n471) );
  MUX2X1 U933 ( .B(n471), .A(n537), .S(n476), .Y(n1396) );
  INVX2 U934 ( .A(\memory[12][3] ), .Y(n472) );
  MUX2X1 U935 ( .B(n472), .A(n538), .S(n476), .Y(n1395) );
  INVX2 U936 ( .A(\memory[12][4] ), .Y(n473) );
  MUX2X1 U937 ( .B(n473), .A(n539), .S(n476), .Y(n1394) );
  INVX2 U938 ( .A(\memory[12][5] ), .Y(n474) );
  MUX2X1 U939 ( .B(n474), .A(n154), .S(n476), .Y(n1393) );
  INVX2 U940 ( .A(\memory[12][6] ), .Y(n475) );
  MUX2X1 U941 ( .B(n475), .A(n541), .S(n476), .Y(n1392) );
  INVX2 U942 ( .A(\memory[12][7] ), .Y(n477) );
  MUX2X1 U943 ( .B(n477), .A(n159), .S(n476), .Y(n1391) );
  NAND3X1 U944 ( .A(n115), .B(n160), .C(n479), .Y(n480) );
  MUX2X1 U945 ( .B(n734), .A(n535), .S(n481), .Y(n1464) );
  MUX2X1 U946 ( .B(n733), .A(n536), .S(n481), .Y(n1463) );
  MUX2X1 U947 ( .B(n732), .A(n537), .S(n481), .Y(n1462) );
  MUX2X1 U948 ( .B(n731), .A(n538), .S(n481), .Y(n1461) );
  MUX2X1 U949 ( .B(n730), .A(n539), .S(n481), .Y(n1460) );
  MUX2X1 U950 ( .B(n729), .A(n154), .S(n481), .Y(n1459) );
  MUX2X1 U951 ( .B(n728), .A(n541), .S(n481), .Y(n1458) );
  MUX2X1 U952 ( .B(n727), .A(n159), .S(n481), .Y(n1457) );
  MUX2X1 U953 ( .B(n726), .A(n535), .S(n483), .Y(n1456) );
  MUX2X1 U954 ( .B(n725), .A(n536), .S(n483), .Y(n1455) );
  MUX2X1 U955 ( .B(n724), .A(n537), .S(n483), .Y(n1454) );
  MUX2X1 U956 ( .B(n723), .A(n538), .S(n483), .Y(n1453) );
  MUX2X1 U957 ( .B(n722), .A(n539), .S(n483), .Y(n1452) );
  MUX2X1 U958 ( .B(n721), .A(n154), .S(n483), .Y(n1451) );
  MUX2X1 U959 ( .B(n720), .A(n541), .S(n483), .Y(n1450) );
  MUX2X1 U960 ( .B(n719), .A(n159), .S(n483), .Y(n1449) );
  MUX2X1 U961 ( .B(n718), .A(n144), .S(n485), .Y(n1448) );
  MUX2X1 U962 ( .B(n717), .A(n536), .S(n485), .Y(n1447) );
  MUX2X1 U963 ( .B(n716), .A(n148), .S(n485), .Y(n1446) );
  MUX2X1 U964 ( .B(n715), .A(n150), .S(n485), .Y(n1445) );
  MUX2X1 U965 ( .B(n714), .A(n152), .S(n485), .Y(n1444) );
  MUX2X1 U966 ( .B(n713), .A(n154), .S(n485), .Y(n1443) );
  MUX2X1 U967 ( .B(n712), .A(n541), .S(n485), .Y(n1442) );
  MUX2X1 U968 ( .B(n711), .A(n159), .S(n485), .Y(n1441) );
  MUX2X1 U969 ( .B(n710), .A(n144), .S(n487), .Y(n1440) );
  MUX2X1 U970 ( .B(n709), .A(n536), .S(n487), .Y(n1439) );
  MUX2X1 U971 ( .B(n708), .A(n148), .S(n487), .Y(n1438) );
  MUX2X1 U972 ( .B(n707), .A(n150), .S(n487), .Y(n1437) );
  MUX2X1 U973 ( .B(n706), .A(n152), .S(n487), .Y(n1436) );
  MUX2X1 U974 ( .B(n705), .A(n154), .S(n487), .Y(n1435) );
  MUX2X1 U975 ( .B(n704), .A(n541), .S(n487), .Y(n1434) );
  MUX2X1 U976 ( .B(n703), .A(n159), .S(n487), .Y(n1433) );
  INVX2 U977 ( .A(\memory[7][0] ), .Y(n489) );
  MUX2X1 U978 ( .B(n489), .A(n535), .S(n496), .Y(n1565) );
  INVX2 U979 ( .A(\memory[7][1] ), .Y(n490) );
  MUX2X1 U980 ( .B(n490), .A(n536), .S(n496), .Y(n1566) );
  INVX2 U981 ( .A(\memory[7][2] ), .Y(n491) );
  MUX2X1 U982 ( .B(n491), .A(n537), .S(n496), .Y(n1567) );
  INVX2 U983 ( .A(\memory[7][3] ), .Y(n492) );
  MUX2X1 U984 ( .B(n492), .A(n538), .S(n496), .Y(n1568) );
  INVX2 U985 ( .A(\memory[7][4] ), .Y(n493) );
  MUX2X1 U986 ( .B(n493), .A(n539), .S(n496), .Y(n1569) );
  INVX2 U987 ( .A(\memory[7][5] ), .Y(n494) );
  MUX2X1 U988 ( .B(n494), .A(n154), .S(n496), .Y(n1570) );
  INVX2 U989 ( .A(\memory[7][6] ), .Y(n495) );
  MUX2X1 U990 ( .B(n495), .A(n541), .S(n496), .Y(n1571) );
  INVX2 U991 ( .A(\memory[7][7] ), .Y(n497) );
  MUX2X1 U992 ( .B(n497), .A(n159), .S(n496), .Y(n1572) );
  INVX2 U993 ( .A(\memory[6][0] ), .Y(n499) );
  MUX2X1 U994 ( .B(n499), .A(n535), .S(n506), .Y(n1575) );
  INVX2 U995 ( .A(\memory[6][1] ), .Y(n500) );
  MUX2X1 U996 ( .B(n500), .A(n536), .S(n506), .Y(n1576) );
  INVX2 U997 ( .A(\memory[6][2] ), .Y(n501) );
  MUX2X1 U998 ( .B(n501), .A(n537), .S(n506), .Y(n1577) );
  INVX2 U999 ( .A(\memory[6][3] ), .Y(n502) );
  MUX2X1 U1000 ( .B(n502), .A(n538), .S(n506), .Y(n1578) );
  INVX2 U1001 ( .A(\memory[6][4] ), .Y(n503) );
  MUX2X1 U1002 ( .B(n503), .A(n539), .S(n506), .Y(n1579) );
  INVX2 U1003 ( .A(\memory[6][5] ), .Y(n504) );
  MUX2X1 U1004 ( .B(n504), .A(n154), .S(n506), .Y(n1580) );
  INVX2 U1005 ( .A(\memory[6][6] ), .Y(n505) );
  MUX2X1 U1006 ( .B(n505), .A(n541), .S(n506), .Y(n1581) );
  INVX2 U1007 ( .A(\memory[6][7] ), .Y(n507) );
  MUX2X1 U1008 ( .B(n507), .A(n158), .S(n506), .Y(n1582) );
  INVX2 U1009 ( .A(\memory[5][0] ), .Y(n509) );
  MUX2X1 U1010 ( .B(n509), .A(n535), .S(n516), .Y(n1585) );
  INVX2 U1011 ( .A(\memory[5][1] ), .Y(n510) );
  MUX2X1 U1012 ( .B(n510), .A(n536), .S(n516), .Y(n1586) );
  INVX2 U1013 ( .A(\memory[5][2] ), .Y(n511) );
  MUX2X1 U1014 ( .B(n511), .A(n537), .S(n516), .Y(n1587) );
  INVX2 U1015 ( .A(\memory[5][3] ), .Y(n512) );
  MUX2X1 U1016 ( .B(n512), .A(n538), .S(n516), .Y(n1588) );
  INVX2 U1017 ( .A(\memory[5][4] ), .Y(n513) );
  MUX2X1 U1018 ( .B(n513), .A(n539), .S(n516), .Y(n1589) );
  INVX2 U1019 ( .A(\memory[5][5] ), .Y(n514) );
  MUX2X1 U1020 ( .B(n514), .A(n154), .S(n516), .Y(n1590) );
  INVX2 U1021 ( .A(\memory[5][6] ), .Y(n515) );
  MUX2X1 U1022 ( .B(n515), .A(n541), .S(n516), .Y(n1591) );
  INVX2 U1023 ( .A(\memory[5][7] ), .Y(n517) );
  MUX2X1 U1024 ( .B(n517), .A(n159), .S(n516), .Y(n1592) );
  INVX2 U1025 ( .A(\memory[4][0] ), .Y(n519) );
  MUX2X1 U1026 ( .B(n519), .A(n535), .S(n526), .Y(n1595) );
  INVX2 U1027 ( .A(\memory[4][1] ), .Y(n520) );
  MUX2X1 U1028 ( .B(n520), .A(n536), .S(n526), .Y(n1596) );
  INVX2 U1029 ( .A(\memory[4][2] ), .Y(n521) );
  MUX2X1 U1030 ( .B(n521), .A(n537), .S(n526), .Y(n1597) );
  INVX2 U1031 ( .A(\memory[4][3] ), .Y(n522) );
  MUX2X1 U1032 ( .B(n522), .A(n538), .S(n526), .Y(n1598) );
  INVX2 U1033 ( .A(\memory[4][4] ), .Y(n523) );
  MUX2X1 U1034 ( .B(n523), .A(n539), .S(n526), .Y(n1599) );
  INVX2 U1035 ( .A(\memory[4][5] ), .Y(n524) );
  MUX2X1 U1036 ( .B(n524), .A(n154), .S(n526), .Y(n1600) );
  INVX2 U1037 ( .A(\memory[4][6] ), .Y(n525) );
  MUX2X1 U1038 ( .B(n525), .A(n541), .S(n526), .Y(n1601) );
  INVX2 U1039 ( .A(\memory[4][7] ), .Y(n527) );
  MUX2X1 U1040 ( .B(n527), .A(n158), .S(n526), .Y(n1602) );
  MUX2X1 U1041 ( .B(n693), .A(n535), .S(n529), .Y(n1423) );
  MUX2X1 U1042 ( .B(n694), .A(n146), .S(n529), .Y(n1424) );
  MUX2X1 U1043 ( .B(n695), .A(n537), .S(n529), .Y(n1425) );
  MUX2X1 U1044 ( .B(n696), .A(n538), .S(n529), .Y(n1426) );
  MUX2X1 U1045 ( .B(n697), .A(n539), .S(n529), .Y(n1427) );
  MUX2X1 U1046 ( .B(n698), .A(n154), .S(n529), .Y(n1428) );
  MUX2X1 U1047 ( .B(n699), .A(n156), .S(n529), .Y(n1429) );
  MUX2X1 U1048 ( .B(n700), .A(n159), .S(n529), .Y(n1430) );
  MUX2X1 U1049 ( .B(n685), .A(n535), .S(n531), .Y(n1415) );
  MUX2X1 U1050 ( .B(n686), .A(n146), .S(n531), .Y(n1416) );
  MUX2X1 U1051 ( .B(n687), .A(n537), .S(n531), .Y(n1417) );
  MUX2X1 U1052 ( .B(n688), .A(n538), .S(n531), .Y(n1418) );
  MUX2X1 U1053 ( .B(n689), .A(n539), .S(n531), .Y(n1419) );
  MUX2X1 U1054 ( .B(n690), .A(n154), .S(n531), .Y(n1420) );
  MUX2X1 U1055 ( .B(n691), .A(n156), .S(n531), .Y(n1421) );
  MUX2X1 U1056 ( .B(n692), .A(n158), .S(n531), .Y(n1422) );
  MUX2X1 U1057 ( .B(n677), .A(n535), .S(n533), .Y(n1407) );
  MUX2X1 U1058 ( .B(n678), .A(n146), .S(n533), .Y(n1408) );
  MUX2X1 U1059 ( .B(n679), .A(n537), .S(n533), .Y(n1409) );
  MUX2X1 U1060 ( .B(n680), .A(n538), .S(n533), .Y(n1410) );
  MUX2X1 U1061 ( .B(n681), .A(n539), .S(n533), .Y(n1411) );
  MUX2X1 U1062 ( .B(n682), .A(n154), .S(n533), .Y(n1412) );
  MUX2X1 U1063 ( .B(n683), .A(n156), .S(n533), .Y(n1413) );
  MUX2X1 U1064 ( .B(n684), .A(n159), .S(n533), .Y(n1414) );
  MUX2X1 U1065 ( .B(n669), .A(n535), .S(n542), .Y(n1399) );
  MUX2X1 U1066 ( .B(n670), .A(n146), .S(n542), .Y(n1400) );
  MUX2X1 U1067 ( .B(n671), .A(n537), .S(n542), .Y(n1401) );
  MUX2X1 U1068 ( .B(n672), .A(n538), .S(n542), .Y(n1402) );
  MUX2X1 U1069 ( .B(n673), .A(n539), .S(n542), .Y(n1403) );
  MUX2X1 U1070 ( .B(n674), .A(n154), .S(n542), .Y(n1404) );
  MUX2X1 U1071 ( .B(n675), .A(n156), .S(n542), .Y(n1405) );
  MUX2X1 U1072 ( .B(n676), .A(n158), .S(n542), .Y(n1406) );
  AND2X2 U1073 ( .A(state), .B(n543), .Y(N338) );
  XOR2X1 U1074 ( .A(n25), .B(n88), .Y(n544) );
  INVX2 U1075 ( .A(state), .Y(n615) );
  NOR2X1 U1076 ( .A(n544), .B(n615), .Y(N339) );
  NAND2X1 U1077 ( .A(n130), .B(n611), .Y(n547) );
  OAI21X1 U1078 ( .A(n131), .B(n611), .C(n25), .Y(n546) );
  AND2X2 U1079 ( .A(n547), .B(n546), .Y(n552) );
  XNOR2X1 U1080 ( .A(n552), .B(n548), .Y(n549) );
  AND2X2 U1081 ( .A(state), .B(n549), .Y(N340) );
  NOR2X1 U1082 ( .A(n70), .B(n618), .Y(n551) );
  NAND2X1 U1083 ( .A(n70), .B(n618), .Y(n550) );
  OAI21X1 U1084 ( .A(n552), .B(n551), .C(n550), .Y(n556) );
  XNOR2X1 U1085 ( .A(n556), .B(n553), .Y(n554) );
  NOR2X1 U1086 ( .A(n554), .B(n615), .Y(N341) );
  NAND2X1 U1087 ( .A(n136), .B(n587), .Y(n557) );
  NOR2X1 U1088 ( .A(n136), .B(n587), .Y(n555) );
  AOI21X1 U1089 ( .A(n557), .B(n556), .C(n555), .Y(n559) );
  XNOR2X1 U1090 ( .A(n559), .B(n558), .Y(n560) );
  AND2X2 U1091 ( .A(state), .B(n560), .Y(N342) );
  NOR2X1 U1092 ( .A(n41), .B(n561), .Y(n566) );
  AND2X2 U1093 ( .A(n563), .B(n562), .Y(n564) );
  NAND3X1 U1094 ( .A(n566), .B(n565), .C(n564), .Y(n567) );
  MUX2X1 U1095 ( .B(n567), .A(n701), .S(RST), .Y(n1431) );
  NAND2X1 U1096 ( .A(n56), .B(n161), .Y(n583) );
  INVX2 U1097 ( .A(n583), .Y(n594) );
  NAND2X1 U1098 ( .A(n594), .B(n54), .Y(n574) );
  NAND2X1 U1099 ( .A(n29), .B(n72), .Y(n585) );
  INVX2 U1100 ( .A(n585), .Y(n597) );
  NAND2X1 U1101 ( .A(n70), .B(n577), .Y(n570) );
  NAND2X1 U1102 ( .A(n570), .B(n118), .Y(n571) );
  NAND2X1 U1103 ( .A(n597), .B(n571), .Y(n573) );
  NAND2X1 U1104 ( .A(n70), .B(n579), .Y(n572) );
  NAND3X1 U1105 ( .A(n574), .B(n573), .C(n572), .Y(n1614) );
  NAND2X1 U1106 ( .A(n594), .B(n576), .Y(n582) );
  NAND2X1 U1107 ( .A(n577), .B(n28), .Y(n578) );
  NAND2X1 U1108 ( .A(n597), .B(n578), .Y(n581) );
  NAND2X1 U1109 ( .A(n131), .B(n579), .Y(n580) );
  NAND3X1 U1110 ( .A(n582), .B(n581), .C(n580), .Y(n1612) );
  AND2X2 U1111 ( .A(n585), .B(n583), .Y(n584) );
  MUX2X1 U1112 ( .B(n584), .A(n56), .S(n133), .Y(n1610) );
  OAI21X1 U1113 ( .A(n6), .B(n585), .C(n56), .Y(n596) );
  NAND2X1 U1114 ( .A(n100), .B(n596), .Y(n590) );
  NAND3X1 U1115 ( .A(n597), .B(n6), .C(n587), .Y(n595) );
  XOR2X1 U1116 ( .A(n587), .B(n31), .Y(n588) );
  NAND2X1 U1117 ( .A(n588), .B(n594), .Y(n589) );
  NAND3X1 U1118 ( .A(n590), .B(n595), .C(n589), .Y(n1608) );
  XOR2X1 U1119 ( .A(n48), .B(n591), .Y(n593) );
  NAND2X1 U1120 ( .A(n594), .B(n593), .Y(n603) );
  INVX2 U1121 ( .A(n595), .Y(n601) );
  INVX2 U1122 ( .A(n596), .Y(n599) );
  NAND2X1 U1123 ( .A(n597), .B(n101), .Y(n598) );
  NAND2X1 U1124 ( .A(n599), .B(n598), .Y(n600) );
  MUX2X1 U1125 ( .B(n601), .A(n600), .S(n52), .Y(n602) );
  NAND2X1 U1126 ( .A(n603), .B(n602), .Y(n1607) );
  NAND2X1 U1127 ( .A(n87), .B(n34), .Y(n607) );
  INVX2 U1128 ( .A(n607), .Y(n604) );
  NAND2X1 U1129 ( .A(n604), .B(n136), .Y(n605) );
  XNOR2X1 U1130 ( .A(n605), .B(n620), .Y(n606) );
  NOR2X1 U1131 ( .A(n615), .B(n606), .Y(N347) );
  XNOR2X1 U1132 ( .A(n607), .B(n619), .Y(n608) );
  NOR2X1 U1133 ( .A(n615), .B(n608), .Y(N346) );
  NAND2X1 U1134 ( .A(n86), .B(n34), .Y(n610) );
  OAI21X1 U1135 ( .A(n612), .B(n611), .C(n43), .Y(n609) );
  AOI21X1 U1136 ( .A(n610), .B(n609), .C(n615), .Y(N345) );
  XNOR2X1 U1137 ( .A(n612), .B(n611), .Y(n613) );
  NOR2X1 U1138 ( .A(n615), .B(n613), .Y(N344) );
  XNOR2X1 U1139 ( .A(n614), .B(n57), .Y(n616) );
  NOR2X1 U1140 ( .A(n616), .B(n615), .Y(N343) );
  INVX1 U1141 ( .A(FULL), .Y(n701) );
  INVX1 U1142 ( .A(EMPTY), .Y(n702) );
  NAND2X1 U1143 ( .A(n784), .B(n785), .Y(n783) );
  NOR2X1 U1144 ( .A(n786), .B(n787), .Y(n785) );
  NAND3X1 U1145 ( .A(n788), .B(n789), .C(n790), .Y(n787) );
  NOR2X1 U1146 ( .A(n791), .B(n792), .Y(n790) );
  OAI22X1 U1147 ( .A(n735), .B(n121), .C(n743), .D(n120), .Y(n792) );
  OAI22X1 U1148 ( .A(n751), .B(n102), .C(n759), .D(n104), .Y(n791) );
  AOI22X1 U1149 ( .A(n79), .B(\memory[23][7] ), .C(n75), .D(\memory[22][7] ), 
        .Y(n789) );
  AOI22X1 U1150 ( .A(n795), .B(\memory[21][7] ), .C(n796), .D(\memory[20][7] ), 
        .Y(n788) );
  NAND3X1 U1151 ( .A(n797), .B(n798), .C(n799), .Y(n786) );
  NOR2X1 U1152 ( .A(n800), .B(n801), .Y(n799) );
  OAI22X1 U1153 ( .A(n661), .B(n123), .C(n653), .D(n122), .Y(n801) );
  OAI22X1 U1154 ( .A(n645), .B(n105), .C(n637), .D(n107), .Y(n800) );
  AOI22X1 U1155 ( .A(n80), .B(\memory[31][7] ), .C(n77), .D(\memory[30][7] ), 
        .Y(n798) );
  AOI22X1 U1156 ( .A(n803), .B(\memory[29][7] ), .C(n804), .D(\memory[28][7] ), 
        .Y(n797) );
  NOR2X1 U1157 ( .A(n805), .B(n806), .Y(n784) );
  NAND3X1 U1158 ( .A(n807), .B(n808), .C(n809), .Y(n806) );
  NOR2X1 U1159 ( .A(n810), .B(n811), .Y(n809) );
  OAI22X1 U1160 ( .A(n700), .B(n108), .C(n692), .D(n110), .Y(n811) );
  OAI22X1 U1161 ( .A(n684), .B(n125), .C(n676), .D(n124), .Y(n810) );
  AOI22X1 U1162 ( .A(n813), .B(\memory[4][7] ), .C(n814), .D(\memory[5][7] ), 
        .Y(n808) );
  AOI22X1 U1163 ( .A(n81), .B(\memory[6][7] ), .C(n76), .D(\memory[7][7] ), 
        .Y(n807) );
  NAND3X1 U1164 ( .A(n815), .B(n816), .C(n817), .Y(n805) );
  NOR2X1 U1165 ( .A(n818), .B(n819), .Y(n817) );
  OAI22X1 U1166 ( .A(n703), .B(n127), .C(n711), .D(n126), .Y(n819) );
  OAI22X1 U1167 ( .A(n719), .B(n111), .C(n727), .D(n112), .Y(n818) );
  AOI22X1 U1168 ( .A(n78), .B(\memory[15][7] ), .C(n74), .D(\memory[14][7] ), 
        .Y(n816) );
  AOI22X1 U1169 ( .A(n820), .B(\memory[13][7] ), .C(n821), .D(\memory[12][7] ), 
        .Y(n815) );
  NAND2X1 U1170 ( .A(n823), .B(n824), .Y(n822) );
  NOR2X1 U1171 ( .A(n825), .B(n826), .Y(n824) );
  NAND3X1 U1172 ( .A(n827), .B(n828), .C(n829), .Y(n826) );
  NOR2X1 U1173 ( .A(n830), .B(n831), .Y(n829) );
  OAI22X1 U1174 ( .A(n736), .B(n121), .C(n744), .D(n120), .Y(n831) );
  OAI22X1 U1175 ( .A(n752), .B(n102), .C(n760), .D(n104), .Y(n830) );
  AOI22X1 U1176 ( .A(n79), .B(\memory[23][6] ), .C(n75), .D(\memory[22][6] ), 
        .Y(n828) );
  AOI22X1 U1177 ( .A(n795), .B(\memory[21][6] ), .C(n796), .D(\memory[20][6] ), 
        .Y(n827) );
  NAND3X1 U1178 ( .A(n832), .B(n833), .C(n834), .Y(n825) );
  NOR2X1 U1179 ( .A(n835), .B(n836), .Y(n834) );
  OAI22X1 U1180 ( .A(n662), .B(n123), .C(n654), .D(n122), .Y(n836) );
  OAI22X1 U1181 ( .A(n646), .B(n105), .C(n638), .D(n107), .Y(n835) );
  AOI22X1 U1182 ( .A(n80), .B(\memory[31][6] ), .C(n77), .D(\memory[30][6] ), 
        .Y(n833) );
  AOI22X1 U1183 ( .A(n803), .B(\memory[29][6] ), .C(n804), .D(\memory[28][6] ), 
        .Y(n832) );
  NOR2X1 U1184 ( .A(n837), .B(n838), .Y(n823) );
  NAND3X1 U1185 ( .A(n839), .B(n840), .C(n841), .Y(n838) );
  NOR2X1 U1186 ( .A(n842), .B(n843), .Y(n841) );
  OAI22X1 U1187 ( .A(n699), .B(n108), .C(n691), .D(n110), .Y(n843) );
  OAI22X1 U1188 ( .A(n683), .B(n125), .C(n675), .D(n124), .Y(n842) );
  AOI22X1 U1189 ( .A(n813), .B(\memory[4][6] ), .C(n814), .D(\memory[5][6] ), 
        .Y(n840) );
  AOI22X1 U1190 ( .A(n81), .B(\memory[6][6] ), .C(n76), .D(\memory[7][6] ), 
        .Y(n839) );
  NAND3X1 U1200 ( .A(n844), .B(n845), .C(n846), .Y(n837) );
  NOR2X1 U1201 ( .A(n852), .B(n861), .Y(n846) );
  OAI22X1 U1203 ( .A(n704), .B(n127), .C(n712), .D(n126), .Y(n861) );
  OAI22X1 U1207 ( .A(n720), .B(n111), .C(n728), .D(n112), .Y(n852) );
  AOI22X1 U1208 ( .A(n78), .B(\memory[15][6] ), .C(n74), .D(\memory[14][6] ), 
        .Y(n845) );
  AOI22X1 U1209 ( .A(n820), .B(\memory[13][6] ), .C(n821), .D(\memory[12][6] ), 
        .Y(n844) );
  NAND2X1 U1210 ( .A(n865), .B(n909), .Y(n863) );
  NOR2X1 U1211 ( .A(n910), .B(n911), .Y(n909) );
  NAND3X1 U1212 ( .A(n912), .B(n913), .C(n914), .Y(n911) );
  NOR2X1 U1213 ( .A(n915), .B(n916), .Y(n914) );
  OAI22X1 U1214 ( .A(n737), .B(n121), .C(n745), .D(n120), .Y(n916) );
  OAI22X1 U1215 ( .A(n753), .B(n102), .C(n761), .D(n104), .Y(n915) );
  AOI22X1 U1216 ( .A(n79), .B(\memory[23][5] ), .C(n75), .D(\memory[22][5] ), 
        .Y(n913) );
  AOI22X1 U1217 ( .A(n795), .B(\memory[21][5] ), .C(n796), .D(\memory[20][5] ), 
        .Y(n912) );
  NAND3X1 U1218 ( .A(n917), .B(n918), .C(n919), .Y(n910) );
  NOR2X1 U1219 ( .A(n920), .B(n921), .Y(n919) );
  OAI22X1 U1220 ( .A(n663), .B(n123), .C(n655), .D(n122), .Y(n921) );
  OAI22X1 U1221 ( .A(n647), .B(n105), .C(n639), .D(n107), .Y(n920) );
  AOI22X1 U1222 ( .A(n80), .B(\memory[31][5] ), .C(n77), .D(\memory[30][5] ), 
        .Y(n918) );
  AOI22X1 U1223 ( .A(n803), .B(\memory[29][5] ), .C(n804), .D(\memory[28][5] ), 
        .Y(n917) );
  NOR2X1 U1224 ( .A(n922), .B(n923), .Y(n865) );
  NAND3X1 U1225 ( .A(n924), .B(n925), .C(n926), .Y(n923) );
  NOR2X1 U1226 ( .A(n927), .B(n928), .Y(n926) );
  OAI22X1 U1227 ( .A(n698), .B(n108), .C(n690), .D(n110), .Y(n928) );
  OAI22X1 U1228 ( .A(n682), .B(n125), .C(n674), .D(n124), .Y(n927) );
  AOI22X1 U1229 ( .A(n813), .B(\memory[4][5] ), .C(n814), .D(\memory[5][5] ), 
        .Y(n925) );
  AOI22X1 U1230 ( .A(n81), .B(\memory[6][5] ), .C(n76), .D(\memory[7][5] ), 
        .Y(n924) );
  NAND3X1 U1231 ( .A(n929), .B(n930), .C(n931), .Y(n922) );
  NOR2X1 U1232 ( .A(n932), .B(n933), .Y(n931) );
  OAI22X1 U1233 ( .A(n705), .B(n127), .C(n713), .D(n126), .Y(n933) );
  OAI22X1 U1234 ( .A(n721), .B(n111), .C(n729), .D(n112), .Y(n932) );
  AOI22X1 U1235 ( .A(n78), .B(\memory[15][5] ), .C(n74), .D(\memory[14][5] ), 
        .Y(n930) );
  AOI22X1 U1236 ( .A(n820), .B(\memory[13][5] ), .C(n821), .D(\memory[12][5] ), 
        .Y(n929) );
  NAND2X1 U1237 ( .A(n935), .B(n936), .Y(n934) );
  NOR2X1 U1238 ( .A(n937), .B(n938), .Y(n936) );
  NAND3X1 U1239 ( .A(n939), .B(n940), .C(n941), .Y(n938) );
  NOR2X1 U1240 ( .A(n942), .B(n943), .Y(n941) );
  OAI22X1 U1241 ( .A(n738), .B(n121), .C(n746), .D(n120), .Y(n943) );
  OAI22X1 U1242 ( .A(n754), .B(n102), .C(n762), .D(n104), .Y(n942) );
  AOI22X1 U1243 ( .A(n79), .B(\memory[23][4] ), .C(n75), .D(\memory[22][4] ), 
        .Y(n940) );
  AOI22X1 U1244 ( .A(n795), .B(\memory[21][4] ), .C(n796), .D(\memory[20][4] ), 
        .Y(n939) );
  NAND3X1 U1245 ( .A(n944), .B(n945), .C(n946), .Y(n937) );
  NOR2X1 U1246 ( .A(n947), .B(n948), .Y(n946) );
  OAI22X1 U1247 ( .A(n664), .B(n123), .C(n656), .D(n122), .Y(n948) );
  OAI22X1 U1248 ( .A(n648), .B(n105), .C(n640), .D(n107), .Y(n947) );
  AOI22X1 U1249 ( .A(n80), .B(\memory[31][4] ), .C(n77), .D(\memory[30][4] ), 
        .Y(n945) );
  AOI22X1 U1250 ( .A(n803), .B(\memory[29][4] ), .C(n804), .D(\memory[28][4] ), 
        .Y(n944) );
  NOR2X1 U1251 ( .A(n949), .B(n950), .Y(n935) );
  NAND3X1 U1252 ( .A(n951), .B(n952), .C(n953), .Y(n950) );
  NOR2X1 U1253 ( .A(n954), .B(n955), .Y(n953) );
  OAI22X1 U1254 ( .A(n697), .B(n108), .C(n689), .D(n110), .Y(n955) );
  OAI22X1 U1255 ( .A(n681), .B(n125), .C(n673), .D(n124), .Y(n954) );
  AOI22X1 U1256 ( .A(n813), .B(\memory[4][4] ), .C(n814), .D(\memory[5][4] ), 
        .Y(n952) );
  AOI22X1 U1257 ( .A(n81), .B(\memory[6][4] ), .C(n76), .D(\memory[7][4] ), 
        .Y(n951) );
  NAND3X1 U1258 ( .A(n956), .B(n957), .C(n958), .Y(n949) );
  NOR2X1 U1259 ( .A(n959), .B(n960), .Y(n958) );
  OAI22X1 U1260 ( .A(n706), .B(n127), .C(n714), .D(n126), .Y(n960) );
  OAI22X1 U1261 ( .A(n722), .B(n111), .C(n730), .D(n112), .Y(n959) );
  AOI22X1 U1262 ( .A(n78), .B(\memory[15][4] ), .C(n74), .D(\memory[14][4] ), 
        .Y(n957) );
  AOI22X1 U1263 ( .A(n820), .B(\memory[13][4] ), .C(n821), .D(\memory[12][4] ), 
        .Y(n956) );
  NAND2X1 U1264 ( .A(n962), .B(n963), .Y(n961) );
  NOR2X1 U1265 ( .A(n964), .B(n965), .Y(n963) );
  NAND3X1 U1266 ( .A(n966), .B(n967), .C(n968), .Y(n965) );
  NOR2X1 U1267 ( .A(n969), .B(n970), .Y(n968) );
  OAI22X1 U1268 ( .A(n739), .B(n121), .C(n747), .D(n120), .Y(n970) );
  OAI22X1 U1269 ( .A(n755), .B(n102), .C(n763), .D(n104), .Y(n969) );
  AOI22X1 U1270 ( .A(n79), .B(\memory[23][3] ), .C(n75), .D(\memory[22][3] ), 
        .Y(n967) );
  AOI22X1 U1271 ( .A(n795), .B(\memory[21][3] ), .C(n796), .D(\memory[20][3] ), 
        .Y(n966) );
  NAND3X1 U1272 ( .A(n971), .B(n972), .C(n973), .Y(n964) );
  NOR2X1 U1273 ( .A(n974), .B(n975), .Y(n973) );
  OAI22X1 U1274 ( .A(n665), .B(n123), .C(n657), .D(n122), .Y(n975) );
  OAI22X1 U1275 ( .A(n649), .B(n105), .C(n641), .D(n107), .Y(n974) );
  AOI22X1 U1276 ( .A(n80), .B(\memory[31][3] ), .C(n77), .D(\memory[30][3] ), 
        .Y(n972) );
  AOI22X1 U1277 ( .A(n803), .B(\memory[29][3] ), .C(n804), .D(\memory[28][3] ), 
        .Y(n971) );
  NOR2X1 U1278 ( .A(n976), .B(n977), .Y(n962) );
  NAND3X1 U1279 ( .A(n978), .B(n979), .C(n980), .Y(n977) );
  NOR2X1 U1280 ( .A(n981), .B(n982), .Y(n980) );
  OAI22X1 U1281 ( .A(n696), .B(n108), .C(n688), .D(n110), .Y(n982) );
  OAI22X1 U1282 ( .A(n680), .B(n125), .C(n672), .D(n124), .Y(n981) );
  AOI22X1 U1283 ( .A(n813), .B(\memory[4][3] ), .C(n814), .D(\memory[5][3] ), 
        .Y(n979) );
  AOI22X1 U1284 ( .A(n81), .B(\memory[6][3] ), .C(n76), .D(\memory[7][3] ), 
        .Y(n978) );
  NAND3X1 U1285 ( .A(n983), .B(n984), .C(n985), .Y(n976) );
  NOR2X1 U1286 ( .A(n986), .B(n987), .Y(n985) );
  OAI22X1 U1287 ( .A(n707), .B(n127), .C(n715), .D(n126), .Y(n987) );
  OAI22X1 U1288 ( .A(n723), .B(n111), .C(n731), .D(n112), .Y(n986) );
  AOI22X1 U1289 ( .A(n78), .B(\memory[15][3] ), .C(n74), .D(\memory[14][3] ), 
        .Y(n984) );
  AOI22X1 U1290 ( .A(n820), .B(\memory[13][3] ), .C(n821), .D(\memory[12][3] ), 
        .Y(n983) );
  NAND2X1 U1291 ( .A(n989), .B(n990), .Y(n988) );
  NOR2X1 U1292 ( .A(n991), .B(n992), .Y(n990) );
  NAND3X1 U1293 ( .A(n993), .B(n994), .C(n995), .Y(n992) );
  NOR2X1 U1294 ( .A(n996), .B(n997), .Y(n995) );
  OAI22X1 U1295 ( .A(n740), .B(n121), .C(n748), .D(n120), .Y(n997) );
  OAI22X1 U1296 ( .A(n756), .B(n102), .C(n764), .D(n104), .Y(n996) );
  AOI22X1 U1297 ( .A(n79), .B(\memory[23][2] ), .C(n75), .D(\memory[22][2] ), 
        .Y(n994) );
  AOI22X1 U1298 ( .A(n795), .B(\memory[21][2] ), .C(n796), .D(\memory[20][2] ), 
        .Y(n993) );
  NAND3X1 U1299 ( .A(n998), .B(n999), .C(n1000), .Y(n991) );
  NOR2X1 U1300 ( .A(n1001), .B(n1002), .Y(n1000) );
  OAI22X1 U1301 ( .A(n666), .B(n123), .C(n658), .D(n122), .Y(n1002) );
  OAI22X1 U1302 ( .A(n650), .B(n105), .C(n642), .D(n107), .Y(n1001) );
  AOI22X1 U1303 ( .A(n80), .B(\memory[31][2] ), .C(n77), .D(\memory[30][2] ), 
        .Y(n999) );
  AOI22X1 U1304 ( .A(n803), .B(\memory[29][2] ), .C(n804), .D(\memory[28][2] ), 
        .Y(n998) );
  NOR2X1 U1305 ( .A(n1003), .B(n1004), .Y(n989) );
  NAND3X1 U1306 ( .A(n1005), .B(n1006), .C(n1007), .Y(n1004) );
  NOR2X1 U1307 ( .A(n1008), .B(n1009), .Y(n1007) );
  OAI22X1 U1308 ( .A(n695), .B(n108), .C(n687), .D(n110), .Y(n1009) );
  OAI22X1 U1309 ( .A(n679), .B(n125), .C(n671), .D(n124), .Y(n1008) );
  AOI22X1 U1310 ( .A(n813), .B(\memory[4][2] ), .C(n814), .D(\memory[5][2] ), 
        .Y(n1006) );
  AOI22X1 U1311 ( .A(n81), .B(\memory[6][2] ), .C(n76), .D(\memory[7][2] ), 
        .Y(n1005) );
  NAND3X1 U1312 ( .A(n1010), .B(n1011), .C(n1012), .Y(n1003) );
  NOR2X1 U1313 ( .A(n1013), .B(n1014), .Y(n1012) );
  OAI22X1 U1314 ( .A(n708), .B(n127), .C(n716), .D(n126), .Y(n1014) );
  OAI22X1 U1315 ( .A(n724), .B(n111), .C(n732), .D(n112), .Y(n1013) );
  AOI22X1 U1316 ( .A(n78), .B(\memory[15][2] ), .C(n74), .D(\memory[14][2] ), 
        .Y(n1011) );
  AOI22X1 U1317 ( .A(n820), .B(\memory[13][2] ), .C(n821), .D(\memory[12][2] ), 
        .Y(n1010) );
  NAND2X1 U1318 ( .A(n1016), .B(n1017), .Y(n1015) );
  NOR2X1 U1319 ( .A(n1018), .B(n1019), .Y(n1017) );
  NAND3X1 U1320 ( .A(n1020), .B(n1021), .C(n1022), .Y(n1019) );
  NOR2X1 U1321 ( .A(n1023), .B(n1024), .Y(n1022) );
  OAI22X1 U1322 ( .A(n741), .B(n121), .C(n749), .D(n120), .Y(n1024) );
  OAI22X1 U1323 ( .A(n757), .B(n102), .C(n765), .D(n104), .Y(n1023) );
  AOI22X1 U1324 ( .A(n79), .B(\memory[23][1] ), .C(n75), .D(\memory[22][1] ), 
        .Y(n1021) );
  AOI22X1 U1325 ( .A(n795), .B(\memory[21][1] ), .C(n796), .D(\memory[20][1] ), 
        .Y(n1020) );
  NAND3X1 U1326 ( .A(n1025), .B(n1026), .C(n1027), .Y(n1018) );
  NOR2X1 U1327 ( .A(n1028), .B(n1029), .Y(n1027) );
  OAI22X1 U1328 ( .A(n667), .B(n123), .C(n659), .D(n122), .Y(n1029) );
  OAI22X1 U1329 ( .A(n651), .B(n105), .C(n643), .D(n107), .Y(n1028) );
  AOI22X1 U1330 ( .A(n80), .B(\memory[31][1] ), .C(n77), .D(\memory[30][1] ), 
        .Y(n1026) );
  AOI22X1 U1331 ( .A(n803), .B(\memory[29][1] ), .C(n804), .D(\memory[28][1] ), 
        .Y(n1025) );
  NOR2X1 U1332 ( .A(n1064), .B(n1065), .Y(n1016) );
  NAND3X1 U1333 ( .A(n1066), .B(n1067), .C(n1068), .Y(n1065) );
  NOR2X1 U1334 ( .A(n1069), .B(n1070), .Y(n1068) );
  OAI22X1 U1335 ( .A(n694), .B(n108), .C(n686), .D(n110), .Y(n1070) );
  OAI22X1 U1336 ( .A(n678), .B(n125), .C(n670), .D(n124), .Y(n1069) );
  AOI22X1 U1337 ( .A(n813), .B(\memory[4][1] ), .C(n814), .D(\memory[5][1] ), 
        .Y(n1067) );
  AOI22X1 U1338 ( .A(n81), .B(\memory[6][1] ), .C(n76), .D(\memory[7][1] ), 
        .Y(n1066) );
  NAND3X1 U1339 ( .A(n1071), .B(n1168), .C(n1169), .Y(n1064) );
  NOR2X1 U1340 ( .A(n1170), .B(n1171), .Y(n1169) );
  OAI22X1 U1341 ( .A(n709), .B(n127), .C(n717), .D(n126), .Y(n1171) );
  OAI22X1 U1342 ( .A(n725), .B(n111), .C(n733), .D(n112), .Y(n1170) );
  AOI22X1 U1343 ( .A(n78), .B(\memory[15][1] ), .C(n74), .D(\memory[14][1] ), 
        .Y(n1168) );
  AOI22X1 U1344 ( .A(n820), .B(\memory[13][1] ), .C(n821), .D(\memory[12][1] ), 
        .Y(n1071) );
  NAND2X1 U1345 ( .A(n1173), .B(n1174), .Y(n1172) );
  NOR2X1 U1346 ( .A(n1175), .B(n1176), .Y(n1174) );
  NAND3X1 U1347 ( .A(n1177), .B(n1178), .C(n1179), .Y(n1176) );
  NOR2X1 U1348 ( .A(n1180), .B(n1181), .Y(n1179) );
  OAI22X1 U1349 ( .A(n742), .B(n121), .C(n750), .D(n120), .Y(n1181) );
  OAI22X1 U1350 ( .A(n758), .B(n102), .C(n766), .D(n104), .Y(n1180) );
  AOI22X1 U1351 ( .A(n79), .B(\memory[23][0] ), .C(n75), .D(\memory[22][0] ), 
        .Y(n1178) );
  AOI22X1 U1352 ( .A(n795), .B(\memory[21][0] ), .C(n796), .D(\memory[20][0] ), 
        .Y(n1177) );
  NAND3X1 U1353 ( .A(n1182), .B(n1183), .C(n1184), .Y(n1175) );
  NOR2X1 U1354 ( .A(n1185), .B(n1186), .Y(n1184) );
  OAI22X1 U1355 ( .A(n668), .B(n123), .C(n660), .D(n122), .Y(n1186) );
  OAI22X1 U1356 ( .A(n652), .B(n105), .C(n644), .D(n107), .Y(n1185) );
  AOI22X1 U1357 ( .A(n80), .B(\memory[31][0] ), .C(n77), .D(\memory[30][0] ), 
        .Y(n1183) );
  AOI22X1 U1358 ( .A(n803), .B(\memory[29][0] ), .C(n804), .D(\memory[28][0] ), 
        .Y(n1182) );
  NOR2X1 U1359 ( .A(n1187), .B(n1188), .Y(n1173) );
  NAND3X1 U1360 ( .A(n1189), .B(n1190), .C(n1191), .Y(n1188) );
  NOR2X1 U1361 ( .A(n1192), .B(n1193), .Y(n1191) );
  OAI22X1 U1362 ( .A(n693), .B(n108), .C(n685), .D(n110), .Y(n1193) );
  OAI22X1 U1363 ( .A(n677), .B(n125), .C(n669), .D(n124), .Y(n1192) );
  AOI22X1 U1364 ( .A(n813), .B(\memory[4][0] ), .C(n814), .D(\memory[5][0] ), 
        .Y(n1190) );
  AOI22X1 U1365 ( .A(n81), .B(\memory[6][0] ), .C(n76), .D(\memory[7][0] ), 
        .Y(n1189) );
  NAND3X1 U1366 ( .A(n1194), .B(n1195), .C(n1196), .Y(n1187) );
  NOR2X1 U1367 ( .A(n1197), .B(n1198), .Y(n1196) );
  OAI22X1 U1368 ( .A(n710), .B(n127), .C(n718), .D(n126), .Y(n1198) );
  OAI22X1 U1369 ( .A(n726), .B(n111), .C(n734), .D(n112), .Y(n1197) );
  AOI22X1 U1370 ( .A(n78), .B(\memory[15][0] ), .C(n74), .D(\memory[14][0] ), 
        .Y(n1195) );
  AOI22X1 U1371 ( .A(n820), .B(\memory[13][0] ), .C(n821), .D(\memory[12][0] ), 
        .Y(n1194) );
  NAND2X1 U1372 ( .A(n1200), .B(n1201), .Y(n1199) );
  NOR2X1 U1373 ( .A(n1202), .B(n1203), .Y(n1201) );
  NAND3X1 U1374 ( .A(n1204), .B(n1205), .C(n1206), .Y(n1203) );
  NOR2X1 U1375 ( .A(n1207), .B(n1208), .Y(n1206) );
  OAI22X1 U1376 ( .A(n775), .B(n121), .C(n777), .D(n120), .Y(n1208) );
  OAI22X1 U1377 ( .A(n779), .B(n102), .C(n781), .D(n104), .Y(n1207) );
  AOI22X1 U1378 ( .A(n79), .B(\opcode[23][1] ), .C(n75), .D(\opcode[22][1] ), 
        .Y(n1205) );
  AOI22X1 U1379 ( .A(n795), .B(\opcode[21][1] ), .C(n796), .D(\opcode[20][1] ), 
        .Y(n1204) );
  NAND3X1 U1380 ( .A(n1209), .B(n1210), .C(n1211), .Y(n1202) );
  NOR2X1 U1381 ( .A(n1212), .B(n1213), .Y(n1211) );
  OAI22X1 U1382 ( .A(n627), .B(n123), .C(n625), .D(n122), .Y(n1213) );
  OAI22X1 U1383 ( .A(n623), .B(n105), .C(n621), .D(n107), .Y(n1212) );
  AOI22X1 U1384 ( .A(n80), .B(\opcode[31][1] ), .C(n77), .D(\opcode[30][1] ), 
        .Y(n1210) );
  AOI22X1 U1385 ( .A(n803), .B(\opcode[29][1] ), .C(n804), .D(\opcode[28][1] ), 
        .Y(n1209) );
  NOR2X1 U1386 ( .A(n1214), .B(n1215), .Y(n1200) );
  NAND3X1 U1387 ( .A(n1216), .B(n1217), .C(n1218), .Y(n1215) );
  NOR2X1 U1388 ( .A(n1219), .B(n1220), .Y(n1218) );
  OAI22X1 U1389 ( .A(n636), .B(n108), .C(n634), .D(n110), .Y(n1220) );
  OAI22X1 U1390 ( .A(n632), .B(n125), .C(n630), .D(n124), .Y(n1219) );
  AOI22X1 U1391 ( .A(n813), .B(\opcode[4][1] ), .C(n814), .D(\opcode[5][1] ), 
        .Y(n1217) );
  AOI22X1 U1392 ( .A(n81), .B(\opcode[6][1] ), .C(n76), .D(\opcode[7][1] ), 
        .Y(n1216) );
  NAND3X1 U1393 ( .A(n1221), .B(n1222), .C(n1223), .Y(n1214) );
  NOR2X1 U1394 ( .A(n1224), .B(n1225), .Y(n1223) );
  OAI22X1 U1395 ( .A(n767), .B(n127), .C(n769), .D(n126), .Y(n1225) );
  OAI22X1 U1396 ( .A(n771), .B(n111), .C(n773), .D(n112), .Y(n1224) );
  AOI22X1 U1397 ( .A(n78), .B(\opcode[15][1] ), .C(n74), .D(\opcode[14][1] ), 
        .Y(n1222) );
  AOI22X1 U1398 ( .A(n820), .B(\opcode[13][1] ), .C(n821), .D(\opcode[12][1] ), 
        .Y(n1221) );
  NAND2X1 U1399 ( .A(n1227), .B(n1228), .Y(n1226) );
  NOR2X1 U1400 ( .A(n1229), .B(n1230), .Y(n1228) );
  NAND3X1 U1401 ( .A(n1231), .B(n1232), .C(n1233), .Y(n1230) );
  NOR2X1 U1402 ( .A(n1234), .B(n1235), .Y(n1233) );
  OAI22X1 U1403 ( .A(n776), .B(n121), .C(n778), .D(n120), .Y(n1235) );
  NAND2X1 U1404 ( .A(n1236), .B(n1237), .Y(n793) );
  OAI22X1 U1405 ( .A(n780), .B(n102), .C(n782), .D(n104), .Y(n1234) );
  AOI22X1 U1406 ( .A(n79), .B(\opcode[23][0] ), .C(n75), .D(\opcode[22][0] ), 
        .Y(n1232) );
  AOI22X1 U1407 ( .A(n795), .B(\opcode[21][0] ), .C(n796), .D(\opcode[20][0] ), 
        .Y(n1231) );
  INVX1 U1408 ( .A(n1240), .Y(n1238) );
  NAND3X1 U1409 ( .A(n57), .B(n619), .C(n53), .Y(n1240) );
  INVX1 U1410 ( .A(n1241), .Y(n1236) );
  NAND3X1 U1411 ( .A(n50), .B(n619), .C(n53), .Y(n1241) );
  NAND3X1 U1412 ( .A(n1242), .B(n1243), .C(n1244), .Y(n1229) );
  NOR2X1 U1413 ( .A(n1245), .B(n1246), .Y(n1244) );
  OAI22X1 U1414 ( .A(n628), .B(n123), .C(n626), .D(n122), .Y(n1246) );
  OAI22X1 U1415 ( .A(n624), .B(n105), .C(n622), .D(n107), .Y(n1245) );
  AOI22X1 U1416 ( .A(n80), .B(\opcode[31][0] ), .C(n77), .D(\opcode[30][0] ), 
        .Y(n1243) );
  AOI22X1 U1417 ( .A(n803), .B(\opcode[29][0] ), .C(n804), .D(\opcode[28][0] ), 
        .Y(n1242) );
  INVX1 U1418 ( .A(n1249), .Y(n1248) );
  NAND3X1 U1419 ( .A(n136), .B(n617), .C(n53), .Y(n1249) );
  INVX1 U1420 ( .A(n1250), .Y(n1247) );
  NAND3X1 U1421 ( .A(n136), .B(n50), .C(n53), .Y(n1250) );
  NOR2X1 U1422 ( .A(n1251), .B(n1252), .Y(n1227) );
  NAND3X1 U1423 ( .A(n1253), .B(n1254), .C(n1255), .Y(n1252) );
  NOR2X1 U1424 ( .A(n1256), .B(n1257), .Y(n1255) );
  OAI22X1 U1425 ( .A(n635), .B(n108), .C(n633), .D(n110), .Y(n1257) );
  OAI22X1 U1426 ( .A(n631), .B(n125), .C(n629), .D(n124), .Y(n1256) );
  AOI22X1 U1427 ( .A(n813), .B(\opcode[4][0] ), .C(n814), .D(\opcode[5][0] ), 
        .Y(n1254) );
  AOI22X1 U1428 ( .A(n81), .B(\opcode[6][0] ), .C(n76), .D(\opcode[7][0] ), 
        .Y(n1253) );
  INVX1 U1429 ( .A(n1260), .Y(n1259) );
  NAND3X1 U1430 ( .A(n619), .B(n620), .C(n50), .Y(n1260) );
  INVX1 U1431 ( .A(n1261), .Y(n1258) );
  NAND3X1 U1432 ( .A(n619), .B(n620), .C(n57), .Y(n1261) );
  NAND3X1 U1433 ( .A(n1262), .B(n1263), .C(n1264), .Y(n1251) );
  NOR2X1 U1434 ( .A(n1265), .B(n1266), .Y(n1264) );
  OAI22X1 U1435 ( .A(n768), .B(n127), .C(n770), .D(n126), .Y(n1266) );
  NOR2X1 U1436 ( .A(n49), .B(n43), .Y(n1237) );
  OAI22X1 U1437 ( .A(n772), .B(n111), .C(n774), .D(n112), .Y(n1265) );
  AOI22X1 U1438 ( .A(n78), .B(\opcode[15][0] ), .C(n74), .D(\opcode[14][0] ), 
        .Y(n1263) );
  AOI22X1 U1439 ( .A(n820), .B(\opcode[13][0] ), .C(n821), .D(\opcode[12][0] ), 
        .Y(n1262) );
  INVX1 U1440 ( .A(n1269), .Y(n1268) );
  NAND3X1 U1441 ( .A(n57), .B(n620), .C(n136), .Y(n1269) );
  NOR2X1 U1442 ( .A(n618), .B(n49), .Y(n1239) );
  INVX1 U1443 ( .A(n1270), .Y(n1267) );
  NAND3X1 U1444 ( .A(n50), .B(n620), .C(n136), .Y(n1270) );
endmodule


module memoryblock_0 ( CLK, NEXT_BYTE, RCV_DATA, RCV_OPCODE, RST, W_ENABLE, 
        EOP, EMPTY, FULL, B_READY, PRGA_IN, PRGA_OPCODE );
  input [7:0] RCV_DATA;
  input [1:0] RCV_OPCODE;
  output [7:0] PRGA_IN;
  output [1:0] PRGA_OPCODE;
  input CLK, NEXT_BYTE, RST, W_ENABLE, EOP;
  output EMPTY, FULL, B_READY;
  wire   R_ENABLE;
  wire   [4:0] BYTE_COUNT;
  wire   [7:0] DATA;
  wire   [1:0] OUT_OPCODE;

  RBUFFER_0 U_0 ( .CLK(CLK), .RST(RST), .NEXT_BYTE(NEXT_BYTE), .DATA(DATA), 
        .OPCODE(OUT_OPCODE), .BYTE_COUNT(BYTE_COUNT), .EOP(EOP), .B_READY(
        B_READY), .R_ENABLE(R_ENABLE), .PRGA_IN(PRGA_IN), .PRGA_OPCODE(
        PRGA_OPCODE) );
  RFIFO_0 U_1 ( .CLK(CLK), .RST(RST), .W_ENABLE(W_ENABLE), .R_ENABLE(R_ENABLE), 
        .RCV_DATA(RCV_DATA), .RCV_OPCODE(RCV_OPCODE), .DATA(DATA), 
        .OUT_OPCODE(OUT_OPCODE), .BYTE_COUNT(BYTE_COUNT), .EMPTY(EMPTY), 
        .FULL(FULL) );
endmodule


module rx_CRC_CALC_0 ( CLK, RST, W_ENABLE, OPCODE, RCV_DATA, RX_CRC );
  input [1:0] OPCODE;
  input [7:0] RCV_DATA;
  output [15:0] RX_CRC;
  input CLK, RST, W_ENABLE;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n100, n102, n104,
         n106, n108, n110, n112, n114, n116, n118, n120, n122, n124, n126,
         n128, n130, n131, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217;
  wire   [15:0] current_crc;
  wire   [15:0] cache_1;

  DFFPOSX1 \cache_1_reg[0]  ( .D(n186), .CLK(CLK), .Q(cache_1[0]) );
  DFFPOSX1 \cache_1_reg[8]  ( .D(n187), .CLK(CLK), .Q(cache_1[8]) );
  DFFPOSX1 \cache_1_reg[15]  ( .D(n188), .CLK(CLK), .Q(cache_1[15]) );
  DFFPOSX1 \cache_1_reg[1]  ( .D(n189), .CLK(CLK), .Q(cache_1[1]) );
  DFFPOSX1 \cache_1_reg[9]  ( .D(n190), .CLK(CLK), .Q(cache_1[9]) );
  DFFPOSX1 \cache_1_reg[2]  ( .D(n191), .CLK(CLK), .Q(cache_1[2]) );
  DFFPOSX1 \cache_1_reg[10]  ( .D(n192), .CLK(CLK), .Q(cache_1[10]) );
  DFFPOSX1 \cache_1_reg[3]  ( .D(n193), .CLK(CLK), .Q(cache_1[3]) );
  DFFPOSX1 \cache_1_reg[11]  ( .D(n194), .CLK(CLK), .Q(cache_1[11]) );
  DFFPOSX1 \cache_1_reg[4]  ( .D(n195), .CLK(CLK), .Q(cache_1[4]) );
  DFFPOSX1 \cache_1_reg[12]  ( .D(n196), .CLK(CLK), .Q(cache_1[12]) );
  DFFPOSX1 \cache_1_reg[5]  ( .D(n197), .CLK(CLK), .Q(cache_1[5]) );
  DFFPOSX1 \cache_1_reg[13]  ( .D(n198), .CLK(CLK), .Q(cache_1[13]) );
  DFFPOSX1 \cache_1_reg[6]  ( .D(n199), .CLK(CLK), .Q(cache_1[6]) );
  DFFPOSX1 \cache_1_reg[14]  ( .D(n200), .CLK(CLK), .Q(cache_1[14]) );
  DFFPOSX1 \cache_1_reg[7]  ( .D(n201), .CLK(CLK), .Q(cache_1[7]) );
  DFFPOSX1 \cache_2_reg[15]  ( .D(n202), .CLK(CLK), .Q(RX_CRC[15]) );
  DFFPOSX1 \cache_2_reg[14]  ( .D(n203), .CLK(CLK), .Q(RX_CRC[14]) );
  DFFPOSX1 \cache_2_reg[13]  ( .D(n204), .CLK(CLK), .Q(RX_CRC[13]) );
  DFFPOSX1 \cache_2_reg[12]  ( .D(n205), .CLK(CLK), .Q(RX_CRC[12]) );
  DFFPOSX1 \cache_2_reg[11]  ( .D(n206), .CLK(CLK), .Q(RX_CRC[11]) );
  DFFPOSX1 \cache_2_reg[10]  ( .D(n207), .CLK(CLK), .Q(RX_CRC[10]) );
  DFFPOSX1 \cache_2_reg[9]  ( .D(n208), .CLK(CLK), .Q(RX_CRC[9]) );
  DFFPOSX1 \cache_2_reg[8]  ( .D(n209), .CLK(CLK), .Q(RX_CRC[8]) );
  DFFPOSX1 \cache_2_reg[7]  ( .D(n210), .CLK(CLK), .Q(RX_CRC[7]) );
  DFFPOSX1 \cache_2_reg[6]  ( .D(n211), .CLK(CLK), .Q(RX_CRC[6]) );
  DFFPOSX1 \cache_2_reg[5]  ( .D(n212), .CLK(CLK), .Q(RX_CRC[5]) );
  DFFPOSX1 \cache_2_reg[4]  ( .D(n213), .CLK(CLK), .Q(RX_CRC[4]) );
  DFFPOSX1 \cache_2_reg[3]  ( .D(n214), .CLK(CLK), .Q(RX_CRC[3]) );
  DFFPOSX1 \cache_2_reg[2]  ( .D(n215), .CLK(CLK), .Q(RX_CRC[2]) );
  DFFPOSX1 \cache_2_reg[1]  ( .D(n216), .CLK(CLK), .Q(RX_CRC[1]) );
  DFFPOSX1 \cache_2_reg[0]  ( .D(n217), .CLK(CLK), .Q(RX_CRC[0]) );
  DFFSR \current_crc_reg[5]  ( .D(n175), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[5]) );
  DFFSR \current_crc_reg[3]  ( .D(n173), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[3]) );
  DFFSR \current_crc_reg[15]  ( .D(n185), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[15]) );
  DFFSR \current_crc_reg[14]  ( .D(n184), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[14]) );
  DFFSR \current_crc_reg[13]  ( .D(n183), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[13]) );
  DFFSR \current_crc_reg[10]  ( .D(n180), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[10]) );
  DFFSR \current_crc_reg[9]  ( .D(n179), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[9]) );
  DFFSR \current_crc_reg[4]  ( .D(n174), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[4]) );
  DFFSR \current_crc_reg[0]  ( .D(n170), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[0]) );
  DFFSR \current_crc_reg[12]  ( .D(n182), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[12]) );
  DFFSR \current_crc_reg[11]  ( .D(n181), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[11]) );
  DFFSR \current_crc_reg[8]  ( .D(n178), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[8]) );
  DFFSR \current_crc_reg[6]  ( .D(n176), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[6]) );
  DFFSR \current_crc_reg[2]  ( .D(n172), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[2]) );
  DFFSR \current_crc_reg[1]  ( .D(n171), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[1]) );
  DFFSR \current_crc_reg[7]  ( .D(n177), .CLK(CLK), .R(n30), .S(1'b1), .Q(
        current_crc[7]) );
  INVX2 U3 ( .A(n79), .Y(n167) );
  INVX8 U20 ( .A(n29), .Y(n26) );
  INVX4 U21 ( .A(n160), .Y(n29) );
  AND2X2 U22 ( .A(W_ENABLE), .B(OPCODE[0]), .Y(n17) );
  INVX8 U23 ( .A(n29), .Y(n27) );
  INVX1 U24 ( .A(OPCODE[1]), .Y(n51) );
  INVX2 U25 ( .A(n18), .Y(n24) );
  INVX2 U26 ( .A(n18), .Y(n25) );
  INVX2 U27 ( .A(n29), .Y(n28) );
  AND2X2 U28 ( .A(n52), .B(n79), .Y(n18) );
  INVX2 U29 ( .A(RST), .Y(n30) );
  XNOR2X1 U30 ( .A(n58), .B(n23), .Y(n59) );
  XNOR2X1 U31 ( .A(RCV_DATA[6]), .B(current_crc[14]), .Y(n156) );
  XNOR2X1 U32 ( .A(RCV_DATA[7]), .B(current_crc[15]), .Y(n124) );
  XOR2X1 U33 ( .A(RCV_DATA[0]), .B(current_crc[8]), .Y(n19) );
  XNOR2X1 U34 ( .A(RCV_DATA[5]), .B(current_crc[13]), .Y(n58) );
  XOR2X1 U35 ( .A(RCV_DATA[1]), .B(current_crc[9]), .Y(n20) );
  XOR2X1 U36 ( .A(RCV_DATA[3]), .B(current_crc[11]), .Y(n21) );
  XOR2X1 U37 ( .A(RCV_DATA[2]), .B(current_crc[10]), .Y(n22) );
  XOR2X1 U38 ( .A(RCV_DATA[4]), .B(current_crc[12]), .Y(n23) );
  INVX2 U39 ( .A(RX_CRC[0]), .Y(n33) );
  INVX2 U40 ( .A(cache_1[0]), .Y(n161) );
  NOR2X1 U41 ( .A(RST), .B(OPCODE[1]), .Y(n31) );
  NAND2X1 U42 ( .A(n31), .B(n17), .Y(n32) );
  INVX2 U43 ( .A(n32), .Y(n160) );
  MUX2X1 U44 ( .B(n33), .A(n161), .S(n26), .Y(n217) );
  INVX2 U45 ( .A(RX_CRC[1]), .Y(n34) );
  INVX2 U46 ( .A(cache_1[1]), .Y(n116) );
  MUX2X1 U47 ( .B(n34), .A(n116), .S(n26), .Y(n216) );
  INVX2 U48 ( .A(RX_CRC[2]), .Y(n35) );
  INVX2 U49 ( .A(cache_1[2]), .Y(n100) );
  MUX2X1 U50 ( .B(n35), .A(n100), .S(n26), .Y(n215) );
  INVX2 U51 ( .A(RX_CRC[3]), .Y(n36) );
  INVX2 U52 ( .A(cache_1[3]), .Y(n77) );
  MUX2X1 U53 ( .B(n36), .A(n77), .S(n26), .Y(n214) );
  INVX2 U54 ( .A(RX_CRC[4]), .Y(n37) );
  INVX2 U55 ( .A(cache_1[4]), .Y(n70) );
  MUX2X1 U56 ( .B(n37), .A(n70), .S(n26), .Y(n213) );
  INVX2 U57 ( .A(RX_CRC[5]), .Y(n38) );
  INVX2 U58 ( .A(cache_1[5]), .Y(n65) );
  MUX2X1 U59 ( .B(n38), .A(n65), .S(n26), .Y(n212) );
  INVX2 U60 ( .A(RX_CRC[6]), .Y(n39) );
  INVX2 U61 ( .A(cache_1[6]), .Y(n57) );
  MUX2X1 U62 ( .B(n39), .A(n57), .S(n26), .Y(n211) );
  INVX2 U63 ( .A(RX_CRC[7]), .Y(n40) );
  INVX2 U64 ( .A(cache_1[7]), .Y(n49) );
  MUX2X1 U65 ( .B(n40), .A(n49), .S(n26), .Y(n210) );
  INVX2 U66 ( .A(RX_CRC[8]), .Y(n41) );
  INVX2 U67 ( .A(cache_1[8]), .Y(n155) );
  MUX2X1 U68 ( .B(n41), .A(n155), .S(n26), .Y(n209) );
  INVX2 U69 ( .A(RX_CRC[9]), .Y(n42) );
  INVX2 U70 ( .A(cache_1[9]), .Y(n108) );
  MUX2X1 U71 ( .B(n42), .A(n108), .S(n26), .Y(n208) );
  INVX2 U72 ( .A(RX_CRC[10]), .Y(n43) );
  INVX2 U73 ( .A(cache_1[10]), .Y(n80) );
  MUX2X1 U74 ( .B(n43), .A(n80), .S(n26), .Y(n207) );
  INVX2 U75 ( .A(RX_CRC[11]), .Y(n44) );
  INVX2 U76 ( .A(cache_1[11]), .Y(n74) );
  MUX2X1 U77 ( .B(n44), .A(n74), .S(n26), .Y(n206) );
  INVX2 U78 ( .A(RX_CRC[12]), .Y(n45) );
  INVX2 U79 ( .A(cache_1[12]), .Y(n67) );
  MUX2X1 U80 ( .B(n45), .A(n67), .S(n26), .Y(n205) );
  INVX2 U81 ( .A(RX_CRC[13]), .Y(n46) );
  INVX2 U82 ( .A(cache_1[13]), .Y(n62) );
  MUX2X1 U83 ( .B(n46), .A(n62), .S(n27), .Y(n204) );
  INVX2 U84 ( .A(RX_CRC[14]), .Y(n47) );
  INVX2 U85 ( .A(cache_1[14]), .Y(n54) );
  MUX2X1 U86 ( .B(n47), .A(n54), .S(n27), .Y(n203) );
  INVX2 U87 ( .A(RX_CRC[15]), .Y(n48) );
  INVX2 U88 ( .A(cache_1[15]), .Y(n148) );
  MUX2X1 U89 ( .B(n48), .A(n148), .S(n27), .Y(n202) );
  INVX2 U90 ( .A(current_crc[7]), .Y(n53) );
  MUX2X1 U91 ( .B(n49), .A(n53), .S(n27), .Y(n201) );
  INVX2 U92 ( .A(n156), .Y(n50) );
  XOR2X1 U93 ( .A(n58), .B(n50), .Y(n164) );
  NAND2X1 U94 ( .A(n17), .B(n51), .Y(n79) );
  NAND2X1 U95 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n52) );
  OAI22X1 U96 ( .A(n164), .B(n79), .C(n24), .D(n53), .Y(n177) );
  INVX2 U97 ( .A(current_crc[14]), .Y(n56) );
  MUX2X1 U98 ( .B(n54), .A(n56), .S(n27), .Y(n200) );
  NAND2X1 U99 ( .A(current_crc[6]), .B(n167), .Y(n55) );
  OAI21X1 U100 ( .A(n25), .B(n56), .C(n55), .Y(n184) );
  INVX2 U101 ( .A(current_crc[6]), .Y(n61) );
  MUX2X1 U102 ( .B(n57), .A(n61), .S(n27), .Y(n199) );
  NAND2X1 U103 ( .A(n167), .B(n59), .Y(n60) );
  OAI21X1 U104 ( .A(n24), .B(n61), .C(n60), .Y(n176) );
  INVX2 U105 ( .A(current_crc[13]), .Y(n64) );
  MUX2X1 U106 ( .B(n62), .A(n64), .S(n27), .Y(n198) );
  NAND2X1 U107 ( .A(current_crc[5]), .B(n167), .Y(n63) );
  OAI21X1 U108 ( .A(n25), .B(n64), .C(n63), .Y(n183) );
  INVX2 U109 ( .A(current_crc[5]), .Y(n66) );
  MUX2X1 U110 ( .B(n65), .A(n66), .S(n27), .Y(n197) );
  XNOR2X1 U111 ( .A(n23), .B(n21), .Y(n118) );
  OAI22X1 U112 ( .A(n118), .B(n79), .C(n25), .D(n66), .Y(n175) );
  INVX2 U113 ( .A(current_crc[12]), .Y(n69) );
  MUX2X1 U114 ( .B(n67), .A(n69), .S(n27), .Y(n196) );
  NAND2X1 U115 ( .A(current_crc[4]), .B(n167), .Y(n68) );
  OAI21X1 U116 ( .A(n24), .B(n69), .C(n68), .Y(n182) );
  INVX2 U117 ( .A(current_crc[4]), .Y(n73) );
  MUX2X1 U118 ( .B(n70), .A(n73), .S(n27), .Y(n195) );
  XOR2X1 U119 ( .A(n21), .B(n22), .Y(n71) );
  NAND2X1 U120 ( .A(n167), .B(n71), .Y(n72) );
  OAI21X1 U121 ( .A(n25), .B(n73), .C(n72), .Y(n174) );
  INVX2 U122 ( .A(current_crc[11]), .Y(n76) );
  MUX2X1 U123 ( .B(n74), .A(n76), .S(n27), .Y(n194) );
  NAND2X1 U124 ( .A(current_crc[3]), .B(n167), .Y(n75) );
  OAI21X1 U125 ( .A(n24), .B(n76), .C(n75), .Y(n181) );
  INVX2 U126 ( .A(current_crc[3]), .Y(n78) );
  MUX2X1 U127 ( .B(n77), .A(n78), .S(n27), .Y(n193) );
  XNOR2X1 U128 ( .A(n22), .B(n20), .Y(n122) );
  OAI22X1 U129 ( .A(n122), .B(n79), .C(n24), .D(n78), .Y(n173) );
  INVX2 U130 ( .A(current_crc[10]), .Y(n82) );
  MUX2X1 U131 ( .B(n80), .A(n82), .S(n27), .Y(n192) );
  NAND2X1 U132 ( .A(current_crc[2]), .B(n167), .Y(n81) );
  OAI21X1 U133 ( .A(n25), .B(n82), .C(n81), .Y(n180) );
  INVX2 U134 ( .A(current_crc[2]), .Y(n106) );
  MUX2X1 U135 ( .B(n100), .A(n106), .S(n28), .Y(n191) );
  XOR2X1 U136 ( .A(n19), .B(n20), .Y(n102) );
  NAND2X1 U137 ( .A(n167), .B(n102), .Y(n104) );
  OAI21X1 U138 ( .A(n24), .B(n106), .C(n104), .Y(n172) );
  INVX2 U139 ( .A(current_crc[9]), .Y(n114) );
  MUX2X1 U140 ( .B(n108), .A(n114), .S(n28), .Y(n190) );
  INVX2 U141 ( .A(n124), .Y(n162) );
  INVX2 U142 ( .A(current_crc[1]), .Y(n131) );
  XNOR2X1 U143 ( .A(n162), .B(n131), .Y(n110) );
  NAND2X1 U144 ( .A(n167), .B(n110), .Y(n112) );
  OAI21X1 U145 ( .A(n25), .B(n114), .C(n112), .Y(n179) );
  MUX2X1 U146 ( .B(n116), .A(n131), .S(n28), .Y(n189) );
  INVX2 U147 ( .A(n118), .Y(n120) );
  XOR2X1 U148 ( .A(n122), .B(n120), .Y(n163) );
  INVX2 U149 ( .A(n163), .Y(n151) );
  XNOR2X1 U150 ( .A(n164), .B(n124), .Y(n126) );
  XNOR2X1 U151 ( .A(n151), .B(n126), .Y(n128) );
  NAND2X1 U152 ( .A(n167), .B(n128), .Y(n130) );
  OAI21X1 U153 ( .A(n24), .B(n131), .C(n130), .Y(n171) );
  INVX2 U154 ( .A(current_crc[15]), .Y(n154) );
  MUX2X1 U155 ( .B(n148), .A(n154), .S(n28), .Y(n188) );
  FAX1 U156 ( .A(current_crc[7]), .B(n19), .C(n162), .YS(n149) );
  XNOR2X1 U157 ( .A(n149), .B(n164), .Y(n150) );
  XOR2X1 U158 ( .A(n151), .B(n150), .Y(n152) );
  NAND2X1 U159 ( .A(n167), .B(n152), .Y(n153) );
  OAI21X1 U160 ( .A(n25), .B(n154), .C(n153), .Y(n185) );
  INVX2 U161 ( .A(current_crc[8]), .Y(n159) );
  MUX2X1 U162 ( .B(n155), .A(n159), .S(n28), .Y(n187) );
  INVX2 U163 ( .A(current_crc[0]), .Y(n169) );
  FAX1 U164 ( .A(n162), .B(n169), .C(n156), .YS(n157) );
  NAND2X1 U165 ( .A(n167), .B(n157), .Y(n158) );
  OAI21X1 U166 ( .A(n24), .B(n159), .C(n158), .Y(n178) );
  MUX2X1 U167 ( .B(n161), .A(n169), .S(n28), .Y(n186) );
  XOR2X1 U168 ( .A(n19), .B(n162), .Y(n165) );
  FAX1 U169 ( .A(n165), .B(n164), .C(n163), .YS(n166) );
  NAND2X1 U170 ( .A(n167), .B(n166), .Y(n168) );
  OAI21X1 U171 ( .A(n25), .B(n169), .C(n168), .Y(n170) );
endmodule


module rx_accumulator_0 ( CLK, RST, RCV_DATA, W_ENABLE, rx_CHECK_CRC );
  input [7:0] RCV_DATA;
  output [15:0] rx_CHECK_CRC;
  input CLK, RST, W_ENABLE;
  wire   n1, n2, n5, n8, n11, n14, n17, n20, n23, n56, n59, n60, n61, n63, n65,
         n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108;

  DFFSR \present_CHECK_CRC_reg[7]  ( .D(n61), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[7]) );
  DFFSR \present_CHECK_CRC_reg[15]  ( .D(n63), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[15]) );
  DFFSR \present_CHECK_CRC_reg[6]  ( .D(n65), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[6]) );
  DFFSR \present_CHECK_CRC_reg[14]  ( .D(n67), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[14]) );
  DFFSR \present_CHECK_CRC_reg[5]  ( .D(n69), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[5]) );
  DFFSR \present_CHECK_CRC_reg[13]  ( .D(n71), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[13]) );
  DFFSR \present_CHECK_CRC_reg[4]  ( .D(n73), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[4]) );
  DFFSR \present_CHECK_CRC_reg[12]  ( .D(n75), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[12]) );
  DFFSR \present_CHECK_CRC_reg[3]  ( .D(n77), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[3]) );
  DFFSR \present_CHECK_CRC_reg[11]  ( .D(n79), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[11]) );
  DFFSR \present_CHECK_CRC_reg[2]  ( .D(n81), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[2]) );
  DFFSR \present_CHECK_CRC_reg[10]  ( .D(n83), .CLK(CLK), .R(n5), .S(1'b1), 
        .Q(rx_CHECK_CRC[10]) );
  DFFSR \present_CHECK_CRC_reg[1]  ( .D(n85), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[1]) );
  DFFSR \present_CHECK_CRC_reg[9]  ( .D(n87), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[9]) );
  DFFSR \present_CHECK_CRC_reg[0]  ( .D(n89), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[0]) );
  DFFSR \present_CHECK_CRC_reg[8]  ( .D(n91), .CLK(CLK), .R(n5), .S(1'b1), .Q(
        rx_CHECK_CRC[8]) );
  OAI21X1 U2 ( .A(n8), .B(n60), .C(n108), .Y(n91) );
  NAND2X1 U3 ( .A(rx_CHECK_CRC[8]), .B(n8), .Y(n108) );
  OAI21X1 U4 ( .A(n2), .B(n60), .C(n107), .Y(n89) );
  NAND2X1 U5 ( .A(RCV_DATA[0]), .B(n2), .Y(n107) );
  OAI21X1 U7 ( .A(n8), .B(n59), .C(n106), .Y(n87) );
  NAND2X1 U8 ( .A(rx_CHECK_CRC[9]), .B(n8), .Y(n106) );
  OAI21X1 U9 ( .A(n2), .B(n59), .C(n105), .Y(n85) );
  NAND2X1 U10 ( .A(RCV_DATA[1]), .B(n2), .Y(n105) );
  OAI21X1 U12 ( .A(n8), .B(n56), .C(n104), .Y(n83) );
  NAND2X1 U13 ( .A(rx_CHECK_CRC[10]), .B(n8), .Y(n104) );
  OAI21X1 U14 ( .A(n2), .B(n56), .C(n103), .Y(n81) );
  NAND2X1 U15 ( .A(RCV_DATA[2]), .B(n2), .Y(n103) );
  OAI21X1 U17 ( .A(n8), .B(n23), .C(n102), .Y(n79) );
  NAND2X1 U18 ( .A(rx_CHECK_CRC[11]), .B(n8), .Y(n102) );
  OAI21X1 U19 ( .A(n2), .B(n23), .C(n101), .Y(n77) );
  NAND2X1 U20 ( .A(RCV_DATA[3]), .B(n2), .Y(n101) );
  OAI21X1 U22 ( .A(n8), .B(n20), .C(n100), .Y(n75) );
  NAND2X1 U23 ( .A(rx_CHECK_CRC[12]), .B(n8), .Y(n100) );
  OAI21X1 U24 ( .A(n2), .B(n20), .C(n99), .Y(n73) );
  NAND2X1 U25 ( .A(RCV_DATA[4]), .B(n2), .Y(n99) );
  OAI21X1 U27 ( .A(n8), .B(n17), .C(n98), .Y(n71) );
  NAND2X1 U28 ( .A(rx_CHECK_CRC[13]), .B(n8), .Y(n98) );
  OAI21X1 U29 ( .A(n2), .B(n17), .C(n97), .Y(n69) );
  NAND2X1 U30 ( .A(RCV_DATA[5]), .B(n2), .Y(n97) );
  OAI21X1 U32 ( .A(n8), .B(n14), .C(n96), .Y(n67) );
  NAND2X1 U33 ( .A(rx_CHECK_CRC[14]), .B(n8), .Y(n96) );
  OAI21X1 U34 ( .A(n2), .B(n14), .C(n95), .Y(n65) );
  NAND2X1 U35 ( .A(RCV_DATA[6]), .B(n2), .Y(n95) );
  OAI21X1 U37 ( .A(n8), .B(n11), .C(n94), .Y(n63) );
  NAND2X1 U38 ( .A(rx_CHECK_CRC[15]), .B(n8), .Y(n94) );
  OAI21X1 U41 ( .A(n2), .B(n11), .C(n93), .Y(n61) );
  NAND2X1 U42 ( .A(RCV_DATA[7]), .B(n2), .Y(n93) );
  INVX4 U6 ( .A(n2), .Y(n8) );
  INVX4 U11 ( .A(n1), .Y(n2) );
  INVX1 U16 ( .A(W_ENABLE), .Y(n1) );
  INVX2 U21 ( .A(RST), .Y(n5) );
  INVX2 U26 ( .A(rx_CHECK_CRC[7]), .Y(n11) );
  INVX2 U31 ( .A(rx_CHECK_CRC[6]), .Y(n14) );
  INVX2 U36 ( .A(rx_CHECK_CRC[5]), .Y(n17) );
  INVX2 U39 ( .A(rx_CHECK_CRC[4]), .Y(n20) );
  INVX2 U40 ( .A(rx_CHECK_CRC[3]), .Y(n23) );
  INVX2 U43 ( .A(rx_CHECK_CRC[2]), .Y(n56) );
  INVX2 U60 ( .A(rx_CHECK_CRC[1]), .Y(n59) );
  INVX2 U61 ( .A(rx_CHECK_CRC[0]), .Y(n60) );
endmodule


module rx_decode_0 ( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP, D_ORIG, BITSTUFF, 
        BS_ERROR );
  input CLK, RST, DP1_RX, SHIFT_ENABLE, EOP;
  output D_ORIG, BITSTUFF, BS_ERROR;
  wire   DP_hold1, DP_hold2, N29, N30, N31, N32, n6, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n18, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n48, n49, n50, n51;
  wire   [3:0] state;

  DFFSR DP_hold2_reg ( .D(n48), .CLK(CLK), .R(1'b1), .S(n9), .Q(DP_hold2) );
  DFFSR \state_reg[3]  ( .D(N32), .CLK(CLK), .R(n9), .S(1'b1), .Q(state[3]) );
  DFFSR DP_hold1_reg ( .D(n49), .CLK(CLK), .R(1'b1), .S(n9), .Q(DP_hold1) );
  NAND2X1 U20 ( .A(n51), .B(n41), .Y(n49) );
  AOI22X1 U21 ( .A(DP_hold1), .B(n42), .C(DP1_RX), .D(n50), .Y(n51) );
  XNOR2X1 U25 ( .A(DP_hold1), .B(DP_hold2), .Y(D_ORIG) );
  DFFSR \state_reg[0]  ( .D(N29), .CLK(CLK), .R(n9), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[2]  ( .D(N31), .CLK(CLK), .R(n9), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[1]  ( .D(N30), .CLK(CLK), .R(n9), .S(1'b1), .Q(state[1]) );
  INVX2 U8 ( .A(RST), .Y(n9) );
  AND2X2 U10 ( .A(state[1]), .B(state[2]), .Y(n6) );
  MUX2X1 U11 ( .B(DP_hold1), .A(DP_hold2), .S(n8), .Y(n40) );
  NAND2X1 U12 ( .A(SHIFT_ENABLE), .B(n50), .Y(n8) );
  INVX1 U13 ( .A(SHIFT_ENABLE), .Y(n31) );
  AND2X1 U14 ( .A(SHIFT_ENABLE), .B(state[0]), .Y(n22) );
  INVX2 U15 ( .A(state[0]), .Y(n15) );
  NOR2X1 U16 ( .A(state[1]), .B(state[2]), .Y(n10) );
  NAND3X1 U17 ( .A(state[3]), .B(n15), .C(n10), .Y(n11) );
  INVX2 U18 ( .A(n11), .Y(BS_ERROR) );
  NAND2X1 U19 ( .A(n6), .B(n15), .Y(n50) );
  NOR2X1 U22 ( .A(state[3]), .B(n50), .Y(BITSTUFF) );
  INVX2 U23 ( .A(n50), .Y(n42) );
  OR2X2 U24 ( .A(EOP), .B(state[3]), .Y(n37) );
  INVX2 U26 ( .A(n37), .Y(n41) );
  INVX2 U27 ( .A(DP1_RX), .Y(n12) );
  XOR2X1 U28 ( .A(n12), .B(DP_hold2), .Y(n33) );
  INVX2 U29 ( .A(n33), .Y(n24) );
  NOR2X1 U30 ( .A(state[0]), .B(n24), .Y(n13) );
  MUX2X1 U31 ( .B(n13), .A(n24), .S(n6), .Y(n14) );
  MUX2X1 U32 ( .B(n15), .A(n14), .S(SHIFT_ENABLE), .Y(n16) );
  AND2X2 U33 ( .A(n41), .B(n16), .Y(N29) );
  INVX2 U34 ( .A(state[2]), .Y(n18) );
  NAND3X1 U35 ( .A(state[1]), .B(n33), .C(n18), .Y(n35) );
  INVX2 U36 ( .A(n35), .Y(n23) );
  INVX2 U37 ( .A(state[1]), .Y(n32) );
  NAND2X1 U38 ( .A(n33), .B(n32), .Y(n20) );
  AOI21X1 U39 ( .A(SHIFT_ENABLE), .B(n20), .C(n18), .Y(n21) );
  AOI21X1 U40 ( .A(n23), .B(n22), .C(n21), .Y(n25) );
  NAND2X1 U41 ( .A(n24), .B(n42), .Y(n29) );
  AOI21X1 U42 ( .A(n25), .B(n29), .C(n37), .Y(N31) );
  NAND3X1 U43 ( .A(n33), .B(n42), .C(SHIFT_ENABLE), .Y(n28) );
  INVX2 U44 ( .A(EOP), .Y(n26) );
  NAND2X1 U45 ( .A(BS_ERROR), .B(n26), .Y(n27) );
  OAI21X1 U46 ( .A(n37), .B(n28), .C(n27), .Y(N32) );
  INVX2 U47 ( .A(n29), .Y(n30) );
  AOI21X1 U48 ( .A(state[1]), .B(n31), .C(n30), .Y(n39) );
  NAND3X1 U49 ( .A(SHIFT_ENABLE), .B(n33), .C(n32), .Y(n34) );
  MUX2X1 U50 ( .B(n35), .A(n34), .S(state[0]), .Y(n36) );
  INVX2 U51 ( .A(n36), .Y(n38) );
  AOI21X1 U52 ( .A(n39), .B(n38), .C(n37), .Y(N30) );
  NAND2X1 U53 ( .A(n41), .B(n40), .Y(n48) );
endmodule


module rx_edgedetect_0 ( CLK, RST, DP1_RX, D_EDGE );
  input CLK, RST, DP1_RX;
  output D_EDGE;
  wire   DP_hold1, DP_hold2, n2, n4;

  DFFSR DP_hold1_reg ( .D(DP1_RX), .CLK(CLK), .R(1'b1), .S(n2), .Q(DP_hold1)
         );
  DFFSR DP_hold2_reg ( .D(DP_hold1), .CLK(CLK), .R(1'b1), .S(n2), .Q(DP_hold2)
         );
  INVX2 U4 ( .A(RST), .Y(n2) );
  XNOR2X1 U6 ( .A(DP_hold2), .B(DP_hold1), .Y(n4) );
  NOR2X1 U7 ( .A(RST), .B(n4), .Y(D_EDGE) );
endmodule


module rx_eopdetect_0 ( DP1_RX, DM1_RX, EOP );
  input DP1_RX, DM1_RX;
  output EOP;


  NOR2X1 U1 ( .A(DP1_RX), .B(DM1_RX), .Y(EOP) );
endmodule


module rx_rcu_0 ( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR, 
        RX_CRC, RX_CHECK_CRC, RCV_DATA, RCVING, W_ENABLE, R_ERROR, CRC_ERROR, 
        OPCODE );
  input [15:0] RX_CRC;
  input [15:0] RX_CHECK_CRC;
  input [7:0] RCV_DATA;
  output [1:0] OPCODE;
  input CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR;
  output RCVING, W_ENABLE, R_ERROR, CRC_ERROR;
  wire   nxtR_ERROR, curR_ERROR, curCRC_ERROR, n1, n2, n3, n4, n5, n6, n7, n8,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n39, n40, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84, n85, n86, n89,
         n90, n91, n92, n93, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n152, n153, n154, n155, n160, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n234, n235, n237, n238, n239, n240,
         n241, n242, n243, n244;
  wire   [3:0] state;
  wire   [3:0] count;
  wire   [3:0] nextstate;

  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(CLK), .R(n43), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(CLK), .R(n43), .S(1'b1), .Q(
        state[0]) );
  DFFSR \count_reg[0]  ( .D(n221), .CLK(CLK), .R(n43), .S(1'b1), .Q(count[0])
         );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(CLK), .R(n43), .S(1'b1), .Q(
        state[2]) );
  DFFPOSX1 curCRC_ERROR_reg ( .D(n234), .CLK(CLK), .Q(curCRC_ERROR) );
  DFFPOSX1 curR_ERROR_reg ( .D(n235), .CLK(CLK), .Q(curR_ERROR) );
  DFFSR R_ERROR_reg ( .D(nxtR_ERROR), .CLK(CLK), .R(n43), .S(1'b1), .Q(R_ERROR) );
  DFFPOSX1 CRC_ERROR_reg ( .D(n222), .CLK(CLK), .Q(CRC_ERROR) );
  NAND2X1 U16 ( .A(n244), .B(n243), .Y(nextstate[2]) );
  OAI21X1 U19 ( .A(n5), .B(n241), .C(n35), .Y(n242) );
  NAND2X1 U20 ( .A(n188), .B(n189), .Y(n241) );
  AOI21X1 U52 ( .A(CRC_ERROR), .B(RST), .C(n238), .Y(n239) );
  OAI21X1 U56 ( .A(n43), .B(n224), .C(n237), .Y(n235) );
  NOR2X1 U79 ( .A(D_EDGE), .B(n23), .Y(n240) );
  DFFSR \count_reg[2]  ( .D(n228), .CLK(CLK), .R(n43), .S(1'b1), .Q(count[2])
         );
  DFFSR \count_reg[1]  ( .D(n229), .CLK(CLK), .R(n43), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[3]  ( .D(n227), .CLK(CLK), .R(n43), .S(1'b1), .Q(count[3])
         );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(CLK), .R(n43), .S(1'b1), .Q(
        state[1]) );
  INVX2 U3 ( .A(n117), .Y(n119) );
  AND2X2 U4 ( .A(n56), .B(n55), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n136) );
  AND2X2 U6 ( .A(n62), .B(n180), .Y(n29) );
  INVX4 U7 ( .A(n40), .Y(n58) );
  BUFX4 U8 ( .A(state[3]), .Y(n33) );
  BUFX2 U9 ( .A(n24), .Y(n2) );
  BUFX2 U10 ( .A(n24), .Y(n3) );
  BUFX2 U11 ( .A(n24), .Y(n4) );
  NAND2X1 U12 ( .A(n217), .B(n216), .Y(n5) );
  AND2X2 U13 ( .A(n40), .B(n170), .Y(n6) );
  AND2X2 U14 ( .A(n119), .B(n116), .Y(n7) );
  AND2X2 U15 ( .A(n67), .B(n39), .Y(n8) );
  INVX2 U23 ( .A(n15), .Y(n13) );
  INVX2 U24 ( .A(n153), .Y(n14) );
  INVX1 U25 ( .A(n6), .Y(n15) );
  NAND2X1 U26 ( .A(n34), .B(n4), .Y(n16) );
  NAND2X1 U27 ( .A(n6), .B(n3), .Y(n17) );
  BUFX2 U28 ( .A(n33), .Y(n18) );
  INVX1 U29 ( .A(n173), .Y(n19) );
  INVX2 U30 ( .A(n19), .Y(n20) );
  INVX2 U31 ( .A(n36), .Y(n39) );
  BUFX2 U32 ( .A(n62), .Y(n21) );
  INVX2 U33 ( .A(n36), .Y(n23) );
  BUFX2 U34 ( .A(state[1]), .Y(n35) );
  MUX2X1 U35 ( .B(n111), .A(n112), .S(n189), .Y(n227) );
  INVX1 U36 ( .A(n104), .Y(n60) );
  AND2X2 U37 ( .A(n119), .B(n110), .Y(n22) );
  NOR2X1 U38 ( .A(n22), .B(n109), .Y(n111) );
  INVX2 U39 ( .A(state[2]), .Y(n36) );
  AND2X2 U40 ( .A(state[1]), .B(n36), .Y(n24) );
  INVX1 U41 ( .A(n4), .Y(n172) );
  NAND2X1 U42 ( .A(n105), .B(n7), .Y(n114) );
  BUFX2 U43 ( .A(n104), .Y(n25) );
  BUFX2 U44 ( .A(n29), .Y(n26) );
  NAND2X1 U45 ( .A(n8), .B(n173), .Y(n62) );
  INVX1 U46 ( .A(n180), .Y(n184) );
  INVX1 U47 ( .A(n58), .Y(n27) );
  INVX1 U48 ( .A(n114), .Y(n106) );
  INVX4 U49 ( .A(n32), .Y(n170) );
  INVX1 U50 ( .A(state[1]), .Y(n67) );
  INVX2 U51 ( .A(n126), .Y(n28) );
  INVX2 U53 ( .A(RST), .Y(n43) );
  INVX1 U54 ( .A(state[1]), .Y(n178) );
  AND2X2 U55 ( .A(SHIFT_ENABLE), .B(n102), .Y(n30) );
  NOR2X1 U57 ( .A(n40), .B(n33), .Y(n31) );
  BUFX2 U58 ( .A(state[3]), .Y(n32) );
  AND2X2 U59 ( .A(n33), .B(n40), .Y(n34) );
  INVX1 U60 ( .A(n34), .Y(n153) );
  BUFX4 U61 ( .A(state[0]), .Y(n40) );
  INVX1 U62 ( .A(n108), .Y(n105) );
  INVX1 U63 ( .A(n113), .Y(n109) );
  INVX1 U64 ( .A(n182), .Y(n126) );
  NAND2X1 U65 ( .A(n39), .B(n170), .Y(n65) );
  INVX2 U66 ( .A(n65), .Y(n146) );
  NAND2X1 U67 ( .A(n35), .B(n146), .Y(n57) );
  INVX2 U68 ( .A(n57), .Y(OPCODE[0]) );
  NAND2X1 U69 ( .A(n33), .B(n39), .Y(n44) );
  NOR2X1 U70 ( .A(n40), .B(n44), .Y(n46) );
  AOI21X1 U71 ( .A(n23), .B(n58), .C(n18), .Y(n45) );
  MUX2X1 U72 ( .B(n46), .A(n45), .S(n35), .Y(n47) );
  NAND2X1 U73 ( .A(n6), .B(n4), .Y(n124) );
  NAND2X1 U74 ( .A(n34), .B(n3), .Y(n182) );
  NAND2X1 U75 ( .A(n124), .B(n182), .Y(n89) );
  OR2X2 U76 ( .A(n89), .B(n47), .Y(OPCODE[1]) );
  NAND2X1 U77 ( .A(n33), .B(n58), .Y(n85) );
  INVX2 U78 ( .A(n85), .Y(n173) );
  INVX2 U80 ( .A(RCV_DATA[1]), .Y(n49) );
  INVX2 U81 ( .A(RCV_DATA[2]), .Y(n48) );
  NAND2X1 U82 ( .A(n49), .B(n48), .Y(n52) );
  INVX2 U83 ( .A(RCV_DATA[0]), .Y(n50) );
  NAND2X1 U84 ( .A(RCV_DATA[7]), .B(n50), .Y(n51) );
  NOR2X1 U85 ( .A(n52), .B(n51), .Y(n56) );
  NOR2X1 U86 ( .A(RCV_DATA[4]), .B(RCV_DATA[3]), .Y(n54) );
  NOR2X1 U87 ( .A(RCV_DATA[6]), .B(RCV_DATA[5]), .Y(n53) );
  AND2X2 U88 ( .A(n54), .B(n53), .Y(n55) );
  NAND3X1 U89 ( .A(n1), .B(n2), .C(n31), .Y(n180) );
  NAND2X1 U90 ( .A(n29), .B(n57), .Y(W_ENABLE) );
  NAND2X1 U91 ( .A(n146), .B(n58), .Y(n166) );
  NAND3X1 U92 ( .A(n34), .B(n23), .C(n178), .Y(n181) );
  OAI21X1 U93 ( .A(n35), .B(n166), .C(n181), .Y(n122) );
  INVX2 U94 ( .A(n122), .Y(n64) );
  NAND2X1 U95 ( .A(n4), .B(n170), .Y(n61) );
  NOR2X1 U96 ( .A(n33), .B(n39), .Y(n59) );
  NAND3X1 U97 ( .A(n40), .B(n67), .C(n59), .Y(n171) );
  NAND3X1 U98 ( .A(n17), .B(n16), .C(n171), .Y(n104) );
  NAND3X1 U99 ( .A(n21), .B(n61), .C(n60), .Y(n63) );
  INVX2 U100 ( .A(n63), .Y(n91) );
  NAND3X1 U101 ( .A(n35), .B(n23), .C(n6), .Y(n130) );
  NAND3X1 U102 ( .A(n64), .B(n91), .C(n130), .Y(RCVING) );
  NAND2X1 U103 ( .A(n240), .B(n20), .Y(n75) );
  NAND2X1 U104 ( .A(n75), .B(n65), .Y(n66) );
  NAND3X1 U105 ( .A(curR_ERROR), .B(n178), .C(n66), .Y(n73) );
  NOR2X1 U106 ( .A(n27), .B(n172), .Y(n69) );
  NAND2X1 U107 ( .A(n1), .B(n170), .Y(n68) );
  NAND2X1 U108 ( .A(n69), .B(n68), .Y(n95) );
  NAND2X1 U109 ( .A(n28), .B(n171), .Y(n71) );
  INVX2 U110 ( .A(n166), .Y(n145) );
  NOR2X1 U111 ( .A(count[3]), .B(n178), .Y(n70) );
  NOR3X1 U112 ( .A(count[0]), .B(count[1]), .C(count[2]), .Y(n188) );
  NAND2X1 U113 ( .A(n70), .B(n188), .Y(n77) );
  AOI22X1 U114 ( .A(EOP), .B(n71), .C(n145), .D(n77), .Y(n72) );
  NAND3X1 U115 ( .A(n73), .B(n95), .C(n72), .Y(nxtR_ERROR) );
  INVX2 U116 ( .A(n73), .Y(n74) );
  OAI21X1 U117 ( .A(n43), .B(n74), .C(nxtR_ERROR), .Y(n237) );
  NAND2X1 U118 ( .A(curCRC_ERROR), .B(n43), .Y(n80) );
  NAND2X1 U119 ( .A(n13), .B(n23), .Y(n81) );
  NAND2X1 U120 ( .A(n81), .B(n75), .Y(n76) );
  NAND2X1 U121 ( .A(n76), .B(n178), .Y(n98) );
  INVX2 U122 ( .A(n77), .Y(n78) );
  NAND2X1 U123 ( .A(n145), .B(n78), .Y(n176) );
  INVX2 U124 ( .A(n176), .Y(n79) );
  NAND3X1 U125 ( .A(n5), .B(n43), .C(n79), .Y(n101) );
  OAI21X1 U126 ( .A(n80), .B(n98), .C(n101), .Y(n238) );
  INVX2 U127 ( .A(count[3]), .Y(n189) );
  INVX2 U128 ( .A(n81), .Y(n84) );
  INVX2 U129 ( .A(D_EDGE), .Y(n82) );
  AOI22X1 U130 ( .A(n84), .B(n82), .C(n226), .D(n145), .Y(n86) );
  MUX2X1 U131 ( .B(n86), .A(n19), .S(n35), .Y(n93) );
  NAND2X1 U132 ( .A(n188), .B(count[3]), .Y(n125) );
  INVX2 U133 ( .A(n125), .Y(n123) );
  NAND2X1 U134 ( .A(n123), .B(n89), .Y(n90) );
  OAI21X1 U135 ( .A(n225), .B(n91), .C(n90), .Y(n92) );
  NOR2X1 U136 ( .A(n93), .B(n92), .Y(n244) );
  OAI21X1 U137 ( .A(n242), .B(n166), .C(n95), .Y(n97) );
  NAND2X1 U138 ( .A(EOP), .B(n25), .Y(n116) );
  NAND2X1 U139 ( .A(n116), .B(n181), .Y(n96) );
  NOR2X1 U140 ( .A(n97), .B(n96), .Y(n243) );
  INVX2 U141 ( .A(n98), .Y(n99) );
  OAI21X1 U142 ( .A(RST), .B(n99), .C(curCRC_ERROR), .Y(n100) );
  NAND2X1 U143 ( .A(n101), .B(n100), .Y(n234) );
  AND2X2 U144 ( .A(count[1]), .B(count[0]), .Y(n103) );
  INVX2 U145 ( .A(BITSTUFF), .Y(n102) );
  NAND2X1 U146 ( .A(n103), .B(n30), .Y(n108) );
  NAND2X1 U147 ( .A(n25), .B(n125), .Y(n117) );
  NAND2X1 U148 ( .A(count[2]), .B(n106), .Y(n112) );
  INVX2 U149 ( .A(count[2]), .Y(n110) );
  INVX2 U150 ( .A(n116), .Y(n107) );
  AOI21X1 U151 ( .A(n119), .B(n108), .C(n107), .Y(n113) );
  MUX2X1 U152 ( .B(n114), .A(n113), .S(count[2]), .Y(n228) );
  NAND3X1 U153 ( .A(n30), .B(n119), .C(n116), .Y(n135) );
  INVX2 U154 ( .A(n135), .Y(n115) );
  NAND2X1 U155 ( .A(count[0]), .B(n115), .Y(n121) );
  INVX2 U156 ( .A(count[0]), .Y(n118) );
  OAI21X1 U157 ( .A(n30), .B(n117), .C(n116), .Y(n133) );
  AOI21X1 U158 ( .A(n119), .B(n118), .C(n133), .Y(n120) );
  MUX2X1 U159 ( .B(n121), .A(n120), .S(count[1]), .Y(n229) );
  NAND2X1 U161 ( .A(n122), .B(EOP), .Y(n132) );
  NAND2X1 U162 ( .A(n123), .B(n226), .Y(n141) );
  OAI21X1 U163 ( .A(n141), .B(n171), .C(n17), .Y(n129) );
  NAND3X1 U164 ( .A(n226), .B(n126), .C(n125), .Y(n127) );
  NAND2X1 U169 ( .A(n26), .B(n127), .Y(n128) );
  OAI21X1 U170 ( .A(n129), .B(n128), .C(n225), .Y(n131) );
  NAND3X1 U171 ( .A(n132), .B(n131), .C(n130), .Y(nextstate[1]) );
  INVX2 U172 ( .A(n133), .Y(n134) );
  MUX2X1 U173 ( .B(n135), .A(n134), .S(count[0]), .Y(n221) );
  NOR2X1 U174 ( .A(n226), .B(n15), .Y(n139) );
  NAND2X1 U175 ( .A(n31), .B(n136), .Y(n137) );
  OAI21X1 U176 ( .A(n153), .B(n141), .C(n137), .Y(n138) );
  OAI21X1 U177 ( .A(n139), .B(n138), .C(n225), .Y(n140) );
  NAND2X1 U178 ( .A(n3), .B(n140), .Y(n164) );
  NOR2X1 U179 ( .A(n141), .B(BS_ERROR), .Y(n142) );
  AOI22X1 U180 ( .A(n142), .B(n13), .C(n14), .D(D_EDGE), .Y(n144) );
  NAND2X1 U181 ( .A(EOP), .B(n14), .Y(n143) );
  MUX2X1 U182 ( .B(n144), .A(n143), .S(n23), .Y(n152) );
  AOI21X1 U183 ( .A(D_EDGE), .B(n146), .C(n145), .Y(n147) );
  OAI21X1 U184 ( .A(n27), .B(n223), .C(n147), .Y(n148) );
  NOR2X1 U185 ( .A(n152), .B(n148), .Y(n155) );
  AND2X2 U186 ( .A(n23), .B(n153), .Y(n154) );
  MUX2X1 U187 ( .B(n155), .A(n154), .S(n35), .Y(n160) );
  NAND2X1 U188 ( .A(n164), .B(n160), .Y(nextstate[0]) );
  NAND2X1 U189 ( .A(D_EDGE), .B(n27), .Y(n165) );
  OAI21X1 U190 ( .A(n225), .B(n170), .C(n165), .Y(n168) );
  NOR2X1 U191 ( .A(n226), .B(n166), .Y(n167) );
  AOI21X1 U192 ( .A(n23), .B(n168), .C(n167), .Y(n169) );
  OAI21X1 U193 ( .A(n223), .B(n170), .C(n169), .Y(n179) );
  OAI21X1 U194 ( .A(n20), .B(n172), .C(n171), .Y(n174) );
  NAND2X1 U195 ( .A(BS_ERROR), .B(n174), .Y(n175) );
  OAI21X1 U196 ( .A(n5), .B(n176), .C(n175), .Y(n177) );
  AOI21X1 U197 ( .A(n179), .B(n178), .C(n177), .Y(n186) );
  OAI21X1 U198 ( .A(EOP), .B(n28), .C(n181), .Y(n183) );
  NOR2X1 U199 ( .A(n184), .B(n183), .Y(n185) );
  NAND2X1 U200 ( .A(n186), .B(n185), .Y(nextstate[3]) );
  XNOR2X1 U201 ( .A(RX_CHECK_CRC[10]), .B(RX_CRC[10]), .Y(n194) );
  XNOR2X1 U202 ( .A(RX_CHECK_CRC[9]), .B(RX_CRC[9]), .Y(n193) );
  XOR2X1 U203 ( .A(RX_CHECK_CRC[7]), .B(RX_CRC[7]), .Y(n191) );
  XOR2X1 U204 ( .A(RX_CHECK_CRC[8]), .B(RX_CRC[8]), .Y(n190) );
  NOR2X1 U205 ( .A(n191), .B(n190), .Y(n192) );
  NAND3X1 U206 ( .A(n194), .B(n193), .C(n192), .Y(n201) );
  XNOR2X1 U207 ( .A(RX_CHECK_CRC[14]), .B(RX_CRC[14]), .Y(n199) );
  XNOR2X1 U208 ( .A(RX_CHECK_CRC[13]), .B(RX_CRC[13]), .Y(n198) );
  XOR2X1 U209 ( .A(RX_CHECK_CRC[11]), .B(RX_CRC[11]), .Y(n196) );
  XOR2X1 U210 ( .A(RX_CHECK_CRC[12]), .B(RX_CRC[12]), .Y(n195) );
  NOR2X1 U211 ( .A(n196), .B(n195), .Y(n197) );
  NAND3X1 U212 ( .A(n199), .B(n198), .C(n197), .Y(n200) );
  NOR2X1 U213 ( .A(n201), .B(n200), .Y(n217) );
  NOR2X1 U214 ( .A(n218), .B(RX_CHECK_CRC[0]), .Y(n202) );
  OAI22X1 U215 ( .A(RX_CRC[1]), .B(n202), .C(n202), .D(n220), .Y(n208) );
  AND2X1 U216 ( .A(RX_CHECK_CRC[0]), .B(n218), .Y(n203) );
  OAI22X1 U217 ( .A(n203), .B(n219), .C(RX_CHECK_CRC[1]), .D(n203), .Y(n207)
         );
  XOR2X1 U218 ( .A(RX_CHECK_CRC[15]), .B(RX_CRC[15]), .Y(n205) );
  XOR2X1 U219 ( .A(RX_CHECK_CRC[2]), .B(RX_CRC[2]), .Y(n204) );
  NOR2X1 U220 ( .A(n205), .B(n204), .Y(n206) );
  NAND3X1 U221 ( .A(n208), .B(n207), .C(n206), .Y(n215) );
  XNOR2X1 U222 ( .A(RX_CHECK_CRC[6]), .B(RX_CRC[6]), .Y(n213) );
  XNOR2X1 U223 ( .A(RX_CHECK_CRC[5]), .B(RX_CRC[5]), .Y(n212) );
  XOR2X1 U224 ( .A(RX_CHECK_CRC[3]), .B(RX_CRC[3]), .Y(n210) );
  XOR2X1 U225 ( .A(RX_CHECK_CRC[4]), .B(RX_CRC[4]), .Y(n209) );
  NOR2X1 U226 ( .A(n210), .B(n209), .Y(n211) );
  NAND3X1 U227 ( .A(n213), .B(n212), .C(n211), .Y(n214) );
  NOR2X1 U228 ( .A(n215), .B(n214), .Y(n216) );
  INVX2 U229 ( .A(RX_CRC[0]), .Y(n218) );
  INVX2 U230 ( .A(RX_CRC[1]), .Y(n219) );
  INVX2 U231 ( .A(RX_CHECK_CRC[1]), .Y(n220) );
  INVX2 U232 ( .A(n239), .Y(n222) );
  INVX2 U233 ( .A(n240), .Y(n223) );
  INVX2 U234 ( .A(curR_ERROR), .Y(n224) );
  INVX2 U235 ( .A(BS_ERROR), .Y(n225) );
  INVX2 U236 ( .A(EOP), .Y(n226) );
endmodule


module rx_shift_reg_0 ( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF, RCV_DATA );
  output [7:0] RCV_DATA;
  input CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF;
  wire   n1, n17, n19, n20, n22, n25, n28, n31, n34, n37, n40, n43, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  wire   [7:0] present_val;

  DFFPOSX1 \RCV_DATA_reg[7]  ( .D(n49), .CLK(CLK), .Q(RCV_DATA[7]) );
  DFFPOSX1 \RCV_DATA_reg[6]  ( .D(n51), .CLK(CLK), .Q(RCV_DATA[6]) );
  DFFPOSX1 \RCV_DATA_reg[5]  ( .D(n53), .CLK(CLK), .Q(RCV_DATA[5]) );
  DFFPOSX1 \RCV_DATA_reg[4]  ( .D(n55), .CLK(CLK), .Q(RCV_DATA[4]) );
  DFFPOSX1 \RCV_DATA_reg[3]  ( .D(n57), .CLK(CLK), .Q(RCV_DATA[3]) );
  DFFPOSX1 \RCV_DATA_reg[2]  ( .D(n59), .CLK(CLK), .Q(RCV_DATA[2]) );
  DFFPOSX1 \RCV_DATA_reg[1]  ( .D(n61), .CLK(CLK), .Q(RCV_DATA[1]) );
  DFFPOSX1 \RCV_DATA_reg[0]  ( .D(n63), .CLK(CLK), .Q(RCV_DATA[0]) );
  OAI21X1 U2 ( .A(RST), .B(n47), .C(n71), .Y(n63) );
  NAND2X1 U3 ( .A(RCV_DATA[0]), .B(RST), .Y(n71) );
  OAI21X1 U6 ( .A(RST), .B(n46), .C(n70), .Y(n61) );
  NAND2X1 U7 ( .A(RCV_DATA[1]), .B(RST), .Y(n70) );
  OAI21X1 U10 ( .A(RST), .B(n45), .C(n69), .Y(n59) );
  NAND2X1 U11 ( .A(RCV_DATA[2]), .B(RST), .Y(n69) );
  OAI21X1 U14 ( .A(RST), .B(n43), .C(n68), .Y(n57) );
  NAND2X1 U15 ( .A(RCV_DATA[3]), .B(RST), .Y(n68) );
  OAI21X1 U18 ( .A(RST), .B(n40), .C(n67), .Y(n55) );
  NAND2X1 U19 ( .A(RCV_DATA[4]), .B(RST), .Y(n67) );
  OAI21X1 U22 ( .A(RST), .B(n37), .C(n66), .Y(n53) );
  NAND2X1 U23 ( .A(RCV_DATA[5]), .B(RST), .Y(n66) );
  OAI21X1 U26 ( .A(RST), .B(n34), .C(n65), .Y(n51) );
  NAND2X1 U27 ( .A(n1), .B(RST), .Y(n65) );
  OAI21X1 U30 ( .A(RST), .B(n31), .C(n64), .Y(n49) );
  NAND2X1 U31 ( .A(n19), .B(RST), .Y(n64) );
  DFFSR \present_val_reg[0]  ( .D(n62), .CLK(CLK), .R(n22), .S(1'b1), .Q(
        present_val[0]) );
  DFFSR \present_val_reg[7]  ( .D(n48), .CLK(CLK), .R(n22), .S(1'b1), .Q(
        present_val[7]) );
  DFFSR \present_val_reg[6]  ( .D(n50), .CLK(CLK), .R(n22), .S(1'b1), .Q(
        present_val[6]) );
  DFFSR \present_val_reg[5]  ( .D(n52), .CLK(CLK), .R(n22), .S(1'b1), .Q(
        present_val[5]) );
  DFFSR \present_val_reg[4]  ( .D(n54), .CLK(CLK), .R(n22), .S(1'b1), .Q(
        present_val[4]) );
  DFFSR \present_val_reg[3]  ( .D(n56), .CLK(CLK), .R(n22), .S(1'b1), .Q(
        present_val[3]) );
  DFFSR \present_val_reg[2]  ( .D(n58), .CLK(CLK), .R(n22), .S(1'b1), .Q(
        present_val[2]) );
  DFFSR \present_val_reg[1]  ( .D(n60), .CLK(CLK), .R(n22), .S(1'b1), .Q(
        present_val[1]) );
  BUFX2 U4 ( .A(RCV_DATA[6]), .Y(n1) );
  INVX1 U21 ( .A(RCV_DATA[7]), .Y(n17) );
  INVX2 U24 ( .A(n17), .Y(n19) );
  INVX2 U25 ( .A(RST), .Y(n22) );
  AND2X2 U28 ( .A(SHIFT_ENABLE), .B(n25), .Y(n20) );
  INVX2 U29 ( .A(present_val[7]), .Y(n31) );
  INVX2 U32 ( .A(present_val[6]), .Y(n34) );
  INVX2 U33 ( .A(present_val[5]), .Y(n37) );
  INVX2 U34 ( .A(present_val[4]), .Y(n40) );
  INVX2 U35 ( .A(present_val[3]), .Y(n43) );
  INVX2 U36 ( .A(present_val[2]), .Y(n45) );
  INVX2 U37 ( .A(present_val[1]), .Y(n46) );
  INVX2 U38 ( .A(present_val[0]), .Y(n47) );
  INVX2 U39 ( .A(BITSTUFF), .Y(n25) );
  MUX2X1 U40 ( .B(n47), .A(n46), .S(n20), .Y(n62) );
  MUX2X1 U41 ( .B(n46), .A(n45), .S(n20), .Y(n60) );
  MUX2X1 U42 ( .B(n45), .A(n43), .S(n20), .Y(n58) );
  MUX2X1 U43 ( .B(n43), .A(n40), .S(n20), .Y(n56) );
  MUX2X1 U44 ( .B(n40), .A(n37), .S(n20), .Y(n54) );
  MUX2X1 U45 ( .B(n37), .A(n34), .S(n20), .Y(n52) );
  MUX2X1 U46 ( .B(n34), .A(n31), .S(n20), .Y(n50) );
  INVX2 U47 ( .A(D_ORIG), .Y(n28) );
  MUX2X1 U48 ( .B(n31), .A(n28), .S(n20), .Y(n48) );
endmodule


module rx_timer_0 ( CLK, RST, D_EDGE, RCVING, SHIFT_ENABLE );
  input CLK, RST, D_EDGE, RCVING;
  output SHIFT_ENABLE;
  wire   state, n5, n7, n9, n10, n11, n12, n13, n14, n16, n19, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36;
  wire   [3:0] count;
  wire   [3:0] nextcount;

  DFFSR state_reg ( .D(n7), .CLK(CLK), .R(n12), .S(1'b1), .Q(state) );
  DFFSR \count_reg[0]  ( .D(nextcount[0]), .CLK(CLK), .R(n12), .S(1'b1), .Q(
        count[0]) );
  DFFSR \count_reg[1]  ( .D(nextcount[1]), .CLK(CLK), .R(n12), .S(1'b1), .Q(
        count[1]) );
  DFFSR \count_reg[2]  ( .D(nextcount[2]), .CLK(CLK), .R(n12), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[3]  ( .D(nextcount[3]), .CLK(CLK), .R(n12), .S(1'b1), .Q(
        count[3]) );
  XOR2X1 U19 ( .A(n34), .B(n27), .Y(n35) );
  NOR2X1 U20 ( .A(count[3]), .B(n28), .Y(n36) );
  XOR2X1 U22 ( .A(n32), .B(count[2]), .Y(n33) );
  NAND2X1 U24 ( .A(state), .B(n30), .Y(nextcount[0]) );
  OAI21X1 U25 ( .A(D_EDGE), .B(n29), .C(n7), .Y(n30) );
  NAND2X1 U30 ( .A(count[0]), .B(count[1]), .Y(n32) );
  XNOR2X1 U32 ( .A(count[0]), .B(count[1]), .Y(n31) );
  INVX1 U7 ( .A(RCVING), .Y(n5) );
  INVX2 U9 ( .A(n5), .Y(n7) );
  NOR2X1 U10 ( .A(n24), .B(n19), .Y(SHIFT_ENABLE) );
  INVX2 U11 ( .A(n9), .Y(nextcount[2]) );
  INVX2 U12 ( .A(RST), .Y(n12) );
  OAI21X1 U13 ( .A(n10), .B(D_EDGE), .C(n7), .Y(n9) );
  NAND2X1 U14 ( .A(n33), .B(state), .Y(n10) );
  NOR2X1 U15 ( .A(D_EDGE), .B(n16), .Y(n11) );
  INVX2 U16 ( .A(count[2]), .Y(n13) );
  OAI21X1 U17 ( .A(n31), .B(n13), .C(n32), .Y(n34) );
  XOR2X1 U18 ( .A(n13), .B(n31), .Y(n27) );
  INVX2 U21 ( .A(n27), .Y(n14) );
  NAND2X1 U23 ( .A(RCVING), .B(n14), .Y(n24) );
  INVX2 U26 ( .A(state), .Y(n16) );
  INVX2 U27 ( .A(n34), .Y(n28) );
  NAND3X1 U28 ( .A(count[3]), .B(n11), .C(n28), .Y(n19) );
  AOI22X1 U29 ( .A(n36), .B(n27), .C(n35), .D(count[3]), .Y(n25) );
  NAND2X1 U31 ( .A(n7), .B(n11), .Y(n26) );
  NOR2X1 U33 ( .A(n25), .B(n26), .Y(nextcount[3]) );
  NOR2X1 U34 ( .A(n31), .B(n26), .Y(nextcount[1]) );
  INVX2 U35 ( .A(count[0]), .Y(n29) );
endmodule


module receiver_block_rewire_0 ( CLK, DM1_RX, DP1_RX, RST, BS_ERROR, CRC_ERROR, 
        EOP_external, OPCODE, RCV_DATA, R_ERROR, W_ENABLE );
  output [1:0] OPCODE;
  output [7:0] RCV_DATA;
  input CLK, DM1_RX, DP1_RX, RST;
  output BS_ERROR, CRC_ERROR, EOP_external, R_ERROR, W_ENABLE;
  wire   n8, n9, SHIFT_ENABLE, BITSTUFF, D_ORIG, D_EDGE, RCVING, n2, n3, n4,
         n5, n6;
  wire   [15:0] RX_CRC;
  wire   [15:0] rx_CHECK_CRC;

  rx_CRC_CALC_0 U_2 ( .CLK(CLK), .RST(RST), .W_ENABLE(n4), .OPCODE(OPCODE), 
        .RCV_DATA(RCV_DATA), .RX_CRC(RX_CRC) );
  rx_accumulator_0 U_3 ( .CLK(CLK), .RST(RST), .RCV_DATA(RCV_DATA), .W_ENABLE(
        n4), .rx_CHECK_CRC(rx_CHECK_CRC) );
  rx_decode_0 U_1 ( .CLK(CLK), .RST(RST), .DP1_RX(DP1_RX), .SHIFT_ENABLE(n5), 
        .EOP(EOP_external), .D_ORIG(D_ORIG), .BITSTUFF(BITSTUFF), .BS_ERROR(
        BS_ERROR) );
  rx_edgedetect_0 U_0 ( .CLK(CLK), .RST(RST), .DP1_RX(DP1_RX), .D_EDGE(D_EDGE)
         );
  rx_eopdetect_0 U_4 ( .DP1_RX(DP1_RX), .DM1_RX(DM1_RX), .EOP(EOP_external) );
  rx_rcu_0 U_5 ( .CLK(CLK), .RST(RST), .D_EDGE(D_EDGE), .EOP(EOP_external), 
        .SHIFT_ENABLE(SHIFT_ENABLE), .BITSTUFF(BITSTUFF), .BS_ERROR(BS_ERROR), 
        .RX_CRC(RX_CRC), .RX_CHECK_CRC(rx_CHECK_CRC), .RCV_DATA({n8, 
        RCV_DATA[6:0]}), .RCVING(RCVING), .W_ENABLE(n9), .R_ERROR(R_ERROR), 
        .CRC_ERROR(CRC_ERROR), .OPCODE(OPCODE) );
  rx_shift_reg_0 U_6 ( .CLK(CLK), .RST(RST), .SHIFT_ENABLE(n3), .D_ORIG(D_ORIG), .BITSTUFF(BITSTUFF), .RCV_DATA({n8, RCV_DATA[6:0]}) );
  rx_timer_0 U_7 ( .CLK(CLK), .RST(RST), .D_EDGE(D_EDGE), .RCVING(RCVING), 
        .SHIFT_ENABLE(SHIFT_ENABLE) );
  BUFX2 U1 ( .A(n8), .Y(RCV_DATA[7]) );
  INVX1 U2 ( .A(SHIFT_ENABLE), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n3) );
  INVX1 U4 ( .A(n6), .Y(n4) );
  BUFX2 U5 ( .A(SHIFT_ENABLE), .Y(n5) );
  INVX4 U6 ( .A(n6), .Y(W_ENABLE) );
  INVX2 U7 ( .A(n9), .Y(n6) );
endmodule


module tx_CRC_CALC_0 ( CLK, RST, EOP, T_STROBE, PRGA_OPCODE, PRGA_OUT, TX_CRC
 );
  input [1:0] PRGA_OPCODE;
  input [7:0] PRGA_OUT;
  output [15:0] TX_CRC;
  input CLK, RST, EOP, T_STROBE;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121;

  OAI22X1 U39 ( .A(n25), .B(n20), .C(n121), .D(n19), .Y(n96) );
  XNOR2X1 U40 ( .A(n119), .B(n79), .Y(n121) );
  OAI22X1 U41 ( .A(n37), .B(n20), .C(n19), .D(n36), .Y(n95) );
  OAI22X1 U42 ( .A(n35), .B(n20), .C(n19), .D(n34), .Y(n94) );
  OAI22X1 U43 ( .A(n33), .B(n20), .C(n19), .D(n32), .Y(n93) );
  OAI22X1 U44 ( .A(n31), .B(n20), .C(n19), .D(n30), .Y(n92) );
  OAI22X1 U45 ( .A(n29), .B(n20), .C(n19), .D(n28), .Y(n91) );
  OAI22X1 U46 ( .A(n27), .B(n20), .C(n118), .D(n19), .Y(n90) );
  XNOR2X1 U47 ( .A(TX_CRC[1]), .B(n117), .Y(n118) );
  OAI22X1 U48 ( .A(n24), .B(n20), .C(n116), .D(n19), .Y(n89) );
  XOR2X1 U49 ( .A(n115), .B(n114), .Y(n116) );
  XNOR2X1 U50 ( .A(TX_CRC[0]), .B(n117), .Y(n115) );
  OAI22X1 U51 ( .A(n79), .B(n20), .C(n113), .D(n19), .Y(n88) );
  OAI22X1 U52 ( .A(n20), .B(n36), .C(n112), .D(n19), .Y(n87) );
  XNOR2X1 U53 ( .A(n111), .B(n110), .Y(n112) );
  OAI22X1 U54 ( .A(n20), .B(n34), .C(n109), .D(n19), .Y(n86) );
  OAI22X1 U55 ( .A(n20), .B(n32), .C(n108), .D(n19), .Y(n85) );
  XNOR2X1 U56 ( .A(n107), .B(n106), .Y(n108) );
  OAI22X1 U57 ( .A(n20), .B(n30), .C(n105), .D(n19), .Y(n84) );
  OAI22X1 U58 ( .A(n20), .B(n28), .C(n104), .D(n19), .Y(n83) );
  XOR2X1 U59 ( .A(n103), .B(n102), .Y(n104) );
  OAI22X1 U60 ( .A(n20), .B(n26), .C(n101), .D(n19), .Y(n82) );
  XOR2X1 U61 ( .A(n100), .B(n99), .Y(n101) );
  XOR2X1 U62 ( .A(n117), .B(n113), .Y(n100) );
  OAI22X1 U63 ( .A(n20), .B(n23), .C(n119), .D(n19), .Y(n81) );
  XOR2X1 U64 ( .A(n98), .B(n97), .Y(n119) );
  XOR2X1 U65 ( .A(n102), .B(n117), .Y(n97) );
  XNOR2X1 U66 ( .A(n25), .B(PRGA_OUT[7]), .Y(n117) );
  XNOR2X1 U67 ( .A(n24), .B(PRGA_OUT[0]), .Y(n102) );
  XOR2X1 U68 ( .A(n113), .B(n99), .Y(n98) );
  XOR2X1 U69 ( .A(n105), .B(n109), .Y(n99) );
  XNOR2X1 U70 ( .A(n106), .B(n111), .Y(n109) );
  XOR2X1 U71 ( .A(TX_CRC[12]), .B(PRGA_OUT[4]), .Y(n111) );
  XOR2X1 U72 ( .A(TX_CRC[11]), .B(PRGA_OUT[3]), .Y(n106) );
  XOR2X1 U74 ( .A(TX_CRC[10]), .B(PRGA_OUT[2]), .Y(n107) );
  XNOR2X1 U75 ( .A(TX_CRC[9]), .B(PRGA_OUT[1]), .Y(n103) );
  XNOR2X1 U76 ( .A(n110), .B(n114), .Y(n113) );
  XNOR2X1 U77 ( .A(n37), .B(PRGA_OUT[6]), .Y(n114) );
  XOR2X1 U78 ( .A(TX_CRC[13]), .B(PRGA_OUT[5]), .Y(n110) );
  NAND3X1 U80 ( .A(PRGA_OPCODE[0]), .B(n80), .C(T_STROBE), .Y(n120) );
  DFFSR \current_crc_reg[6]  ( .D(n87), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[6]) );
  DFFSR \current_crc_reg[5]  ( .D(n86), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[5]) );
  DFFSR \current_crc_reg[4]  ( .D(n85), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[4]) );
  DFFSR \current_crc_reg[3]  ( .D(n84), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[3]) );
  DFFSR \current_crc_reg[2]  ( .D(n83), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[2]) );
  DFFSR \current_crc_reg[1]  ( .D(n82), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[1]) );
  DFFSR \current_crc_reg[0]  ( .D(n81), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[0]) );
  DFFSR \current_crc_reg[15]  ( .D(n96), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[15]) );
  DFFSR \current_crc_reg[9]  ( .D(n90), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[9]) );
  DFFSR \current_crc_reg[8]  ( .D(n89), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[8]) );
  DFFSR \current_crc_reg[14]  ( .D(n95), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[14]) );
  DFFSR \current_crc_reg[13]  ( .D(n94), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[13]) );
  DFFSR \current_crc_reg[12]  ( .D(n93), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[12]) );
  DFFSR \current_crc_reg[11]  ( .D(n92), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[11]) );
  DFFSR \current_crc_reg[10]  ( .D(n91), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[10]) );
  DFFSR \current_crc_reg[7]  ( .D(n88), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[7]) );
  INVX2 U3 ( .A(n17), .Y(n20) );
  INVX1 U20 ( .A(EOP), .Y(n22) );
  INVX2 U21 ( .A(n120), .Y(n18) );
  AND2X2 U22 ( .A(n120), .B(n22), .Y(n17) );
  INVX2 U23 ( .A(RST), .Y(n21) );
  XOR2X1 U24 ( .A(n103), .B(n107), .Y(n105) );
  INVX2 U25 ( .A(n18), .Y(n19) );
  INVX2 U26 ( .A(TX_CRC[0]), .Y(n23) );
  INVX2 U27 ( .A(TX_CRC[8]), .Y(n24) );
  INVX2 U28 ( .A(TX_CRC[15]), .Y(n25) );
  INVX2 U29 ( .A(TX_CRC[1]), .Y(n26) );
  INVX2 U30 ( .A(TX_CRC[9]), .Y(n27) );
  INVX2 U31 ( .A(TX_CRC[2]), .Y(n28) );
  INVX2 U32 ( .A(TX_CRC[10]), .Y(n29) );
  INVX2 U33 ( .A(TX_CRC[3]), .Y(n30) );
  INVX2 U34 ( .A(TX_CRC[11]), .Y(n31) );
  INVX2 U35 ( .A(TX_CRC[4]), .Y(n32) );
  INVX2 U36 ( .A(TX_CRC[12]), .Y(n33) );
  INVX2 U37 ( .A(TX_CRC[5]), .Y(n34) );
  INVX2 U38 ( .A(TX_CRC[13]), .Y(n35) );
  INVX2 U73 ( .A(TX_CRC[6]), .Y(n36) );
  INVX2 U79 ( .A(TX_CRC[14]), .Y(n37) );
  INVX2 U81 ( .A(TX_CRC[7]), .Y(n79) );
  INVX2 U82 ( .A(PRGA_OPCODE[1]), .Y(n80) );
endmodule


module tx_encode_0 ( clk, rst, SHIFT_ENABLE_E, d_encode, EOP, t_bitstuff, 
        dp_tx_out, dm_tx_out );
  input clk, rst, SHIFT_ENABLE_E, d_encode, EOP;
  output t_bitstuff, dp_tx_out, dm_tx_out;
  wire   DE_holdout, DE_holdout_BS, DE_holdout_last, DE_holdout_nxt, dm_tx_nxt,
         n3, n5, n6, n7, n8, n10, n11, n16, n17, n21, n22, n23, n24, n25, n28,
         n29, n30, n31, n33, n34, n35, n36, n38, n42, n45, n46, n47, n48, n51,
         n52, n53, n56, n57, n63, n65, n66, n67, n68, n69, n70, n71, n73, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97;
  wire   [3:0] state;
  wire   [3:0] nextstate;

  DFFSR DE_holdout_reg ( .D(DE_holdout_nxt), .CLK(clk), .R(1'b1), .S(n11), .Q(
        DE_holdout) );
  DFFPOSX1 DE_holdout_last_reg ( .D(n73), .CLK(clk), .Q(DE_holdout_last) );
  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(clk), .R(n11), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n11), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n11), .S(1'b1), .Q(
        state[1]) );
  DFFSR dp_tx_out_reg ( .D(DE_holdout_nxt), .CLK(clk), .R(1'b1), .S(n11), .Q(
        dp_tx_out) );
  DFFSR dm_tx_out_reg ( .D(dm_tx_nxt), .CLK(clk), .R(n11), .S(1'b1), .Q(
        dm_tx_out) );
  OAI21X1 U9 ( .A(n3), .B(n7), .C(n95), .Y(nextstate[1]) );
  OAI21X1 U11 ( .A(n6), .B(n8), .C(n53), .Y(n94) );
  NAND3X1 U12 ( .A(SHIFT_ENABLE_E), .B(n65), .C(n6), .Y(n97) );
  OAI21X1 U14 ( .A(n5), .B(n53), .C(n92), .Y(nextstate[0]) );
  OAI21X1 U15 ( .A(n91), .B(n90), .C(SHIFT_ENABLE_E), .Y(n92) );
  NOR2X1 U18 ( .A(n6), .B(n93), .Y(n91) );
  NAND3X1 U19 ( .A(d_encode), .B(n89), .C(n88), .Y(n93) );
  XNOR2X1 U20 ( .A(n68), .B(n67), .Y(n88) );
  NOR2X1 U22 ( .A(n63), .B(SHIFT_ENABLE_E), .Y(n96) );
  OAI22X1 U23 ( .A(n11), .B(n68), .C(rst), .D(n67), .Y(n73) );
  OAI22X1 U26 ( .A(n10), .B(n69), .C(n67), .D(n87), .Y(n71) );
  NOR2X1 U36 ( .A(EOP), .B(state[3]), .Y(n89) );
  NOR2X1 U37 ( .A(EOP), .B(n84), .Y(n86) );
  AOI22X1 U38 ( .A(n6), .B(n83), .C(n56), .D(n5), .Y(n84) );
  XNOR2X1 U40 ( .A(DE_holdout_BS), .B(n81), .Y(n83) );
  XOR2X1 U46 ( .A(DE_holdout), .B(SHIFT_ENABLE_E), .Y(n82) );
  XNOR2X1 U47 ( .A(n80), .B(n67), .Y(n85) );
  NAND2X1 U49 ( .A(SHIFT_ENABLE_E), .B(n66), .Y(n80) );
  NAND2X1 U55 ( .A(n81), .B(n69), .Y(n79) );
  NAND2X1 U57 ( .A(SHIFT_ENABLE_E), .B(d_encode), .Y(n81) );
  DFFSR DE_holdout_BS_reg ( .D(n71), .CLK(clk), .R(n11), .S(1'b1), .Q(
        DE_holdout_BS) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n11), .S(1'b1), .Q(
        state[2]) );
  INVX2 U3 ( .A(n38), .Y(n3) );
  INVX2 U4 ( .A(state[0]), .Y(n5) );
  INVX2 U5 ( .A(n5), .Y(n6) );
  INVX1 U6 ( .A(state[1]), .Y(n38) );
  BUFX4 U10 ( .A(n70), .Y(t_bitstuff) );
  INVX1 U13 ( .A(n89), .Y(n63) );
  INVX1 U16 ( .A(n52), .Y(n7) );
  INVX1 U17 ( .A(n65), .Y(n8) );
  INVX2 U21 ( .A(rst), .Y(n11) );
  NOR2X1 U24 ( .A(n48), .B(n17), .Y(n10) );
  INVX1 U25 ( .A(n10), .Y(n87) );
  NAND2X1 U27 ( .A(state[2]), .B(state[1]), .Y(n16) );
  NOR3X1 U28 ( .A(state[3]), .B(n16), .C(n5), .Y(n70) );
  INVX2 U29 ( .A(n16), .Y(n31) );
  NAND3X1 U30 ( .A(n89), .B(n5), .C(n31), .Y(n48) );
  INVX2 U31 ( .A(SHIFT_ENABLE_E), .Y(n17) );
  NAND2X1 U32 ( .A(n66), .B(n31), .Y(n21) );
  OAI21X1 U33 ( .A(n63), .B(n21), .C(n48), .Y(n90) );
  INVX2 U34 ( .A(n48), .Y(n22) );
  AOI21X1 U35 ( .A(n94), .B(n3), .C(n22), .Y(n95) );
  INVX2 U39 ( .A(state[2]), .Y(n23) );
  NAND3X1 U41 ( .A(n5), .B(n23), .C(n38), .Y(n51) );
  NAND2X1 U42 ( .A(n51), .B(state[3]), .Y(n36) );
  INVX2 U43 ( .A(n85), .Y(n24) );
  NOR2X1 U44 ( .A(n63), .B(n24), .Y(n25) );
  MUX2X1 U45 ( .B(n25), .A(n86), .S(n31), .Y(n28) );
  NAND2X1 U48 ( .A(n36), .B(n28), .Y(dm_tx_nxt) );
  OAI21X1 U50 ( .A(n69), .B(n81), .C(n79), .Y(n30) );
  AND2X2 U51 ( .A(n82), .B(n5), .Y(n29) );
  AOI21X1 U52 ( .A(n6), .B(n30), .C(n29), .Y(n33) );
  MUX2X1 U53 ( .B(n85), .A(n33), .S(n31), .Y(n34) );
  OAI21X1 U54 ( .A(state[3]), .B(n34), .C(n57), .Y(n35) );
  NAND2X1 U56 ( .A(n36), .B(n35), .Y(DE_holdout_nxt) );
  NAND2X1 U58 ( .A(n52), .B(n3), .Y(n45) );
  AOI21X1 U59 ( .A(n65), .B(n38), .C(n96), .Y(n42) );
  MUX2X1 U60 ( .B(n45), .A(n42), .S(state[2]), .Y(n46) );
  INVX2 U61 ( .A(n46), .Y(n47) );
  NAND2X1 U62 ( .A(n48), .B(n47), .Y(nextstate[2]) );
  AOI21X1 U63 ( .A(state[3]), .B(n51), .C(n57), .Y(nextstate[3]) );
  INVX2 U64 ( .A(n97), .Y(n52) );
  INVX2 U65 ( .A(n96), .Y(n53) );
  INVX2 U68 ( .A(n82), .Y(n56) );
  INVX2 U69 ( .A(EOP), .Y(n57) );
  INVX2 U74 ( .A(n93), .Y(n65) );
  INVX2 U75 ( .A(d_encode), .Y(n66) );
  INVX2 U76 ( .A(DE_holdout), .Y(n67) );
  INVX2 U77 ( .A(DE_holdout_last), .Y(n68) );
  INVX2 U78 ( .A(DE_holdout_BS), .Y(n69) );
endmodule


module tx_shiftreg_0 ( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe, 
        send_data, d_encode );
  input [7:0] send_data;
  input clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe;
  output d_encode;
  wire   n1, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79;
  wire   [7:1] present_val;
  wire   [2:0] count;

  DFFSR \count_reg[0]  ( .D(n69), .CLK(clk), .R(1'b1), .S(n17), .Q(count[0])
         );
  DFFSR \count_reg[1]  ( .D(n71), .CLK(clk), .R(1'b1), .S(n17), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n70), .CLK(clk), .R(1'b1), .S(n17), .Q(count[2])
         );
  DFFSR \present_val_reg[7]  ( .D(n78), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[7]) );
  DFFSR \present_val_reg[6]  ( .D(n77), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[6]) );
  DFFSR \present_val_reg[5]  ( .D(n76), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[5]) );
  DFFSR \present_val_reg[4]  ( .D(n75), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[4]) );
  DFFSR \present_val_reg[3]  ( .D(n74), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[3]) );
  DFFSR \present_val_reg[2]  ( .D(n73), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[2]) );
  DFFSR \present_val_reg[1]  ( .D(n72), .CLK(clk), .R(n17), .S(1'b1), .Q(
        present_val[1]) );
  DFFSR \present_val_reg[0]  ( .D(n79), .CLK(clk), .R(n17), .S(1'b1), .Q(
        d_encode) );
  AND2X2 U3 ( .A(n19), .B(count[2]), .Y(n1) );
  INVX2 U15 ( .A(n20), .Y(n13) );
  OR2X2 U16 ( .A(n13), .B(n15), .Y(n67) );
  INVX2 U17 ( .A(n15), .Y(n16) );
  INVX1 U18 ( .A(t_bitstuff), .Y(n18) );
  AND2X2 U19 ( .A(n67), .B(n16), .Y(n14) );
  INVX2 U20 ( .A(n14), .Y(n68) );
  AND2X2 U21 ( .A(n1), .B(SHIFT_ENABLE_R), .Y(n15) );
  INVX2 U22 ( .A(rst), .Y(n17) );
  INVX1 U23 ( .A(n67), .Y(n56) );
  NAND2X1 U24 ( .A(SHIFT_ENABLE_R), .B(n18), .Y(n20) );
  NAND2X1 U25 ( .A(count[1]), .B(count[0]), .Y(n64) );
  INVX2 U26 ( .A(n64), .Y(n19) );
  NAND2X1 U27 ( .A(d_encode), .B(n56), .Y(n24) );
  NAND2X1 U28 ( .A(present_val[1]), .B(n14), .Y(n23) );
  INVX2 U29 ( .A(send_data[0]), .Y(n21) );
  OR2X2 U30 ( .A(n16), .B(n21), .Y(n22) );
  NAND3X1 U31 ( .A(n24), .B(n23), .C(n22), .Y(n79) );
  NAND2X1 U32 ( .A(present_val[1]), .B(n56), .Y(n28) );
  NAND2X1 U33 ( .A(present_val[2]), .B(n14), .Y(n27) );
  INVX2 U34 ( .A(send_data[1]), .Y(n25) );
  OR2X2 U35 ( .A(n16), .B(n25), .Y(n26) );
  NAND3X1 U36 ( .A(n28), .B(n27), .C(n26), .Y(n72) );
  NAND2X1 U37 ( .A(present_val[2]), .B(n56), .Y(n32) );
  NAND2X1 U38 ( .A(present_val[3]), .B(n14), .Y(n31) );
  INVX2 U39 ( .A(send_data[2]), .Y(n29) );
  OR2X2 U40 ( .A(n16), .B(n29), .Y(n30) );
  NAND3X1 U41 ( .A(n32), .B(n31), .C(n30), .Y(n73) );
  NAND2X1 U42 ( .A(present_val[3]), .B(n56), .Y(n36) );
  NAND2X1 U43 ( .A(present_val[4]), .B(n14), .Y(n35) );
  INVX2 U44 ( .A(send_data[3]), .Y(n33) );
  OR2X2 U45 ( .A(n16), .B(n33), .Y(n34) );
  NAND3X1 U46 ( .A(n36), .B(n35), .C(n34), .Y(n74) );
  NAND2X1 U47 ( .A(present_val[4]), .B(n56), .Y(n40) );
  NAND2X1 U48 ( .A(present_val[5]), .B(n14), .Y(n39) );
  INVX2 U49 ( .A(send_data[4]), .Y(n37) );
  OR2X2 U50 ( .A(n16), .B(n37), .Y(n38) );
  NAND3X1 U51 ( .A(n40), .B(n39), .C(n38), .Y(n75) );
  NAND2X1 U52 ( .A(present_val[5]), .B(n56), .Y(n55) );
  NAND2X1 U53 ( .A(present_val[6]), .B(n14), .Y(n54) );
  INVX2 U54 ( .A(send_data[5]), .Y(n41) );
  OR2X2 U55 ( .A(n16), .B(n41), .Y(n42) );
  NAND3X1 U56 ( .A(n55), .B(n54), .C(n42), .Y(n76) );
  NAND2X1 U57 ( .A(present_val[6]), .B(n56), .Y(n60) );
  NAND2X1 U58 ( .A(present_val[7]), .B(n14), .Y(n59) );
  INVX2 U59 ( .A(send_data[6]), .Y(n57) );
  OR2X2 U60 ( .A(n16), .B(n57), .Y(n58) );
  NAND3X1 U61 ( .A(n60), .B(n59), .C(n58), .Y(n77) );
  INVX2 U62 ( .A(present_val[7]), .Y(n62) );
  INVX2 U63 ( .A(send_data[7]), .Y(n61) );
  OAI22X1 U64 ( .A(n67), .B(n62), .C(n16), .D(n61), .Y(n78) );
  NAND2X1 U65 ( .A(count[2]), .B(n16), .Y(n63) );
  OAI21X1 U66 ( .A(n64), .B(n68), .C(n63), .Y(n70) );
  NAND2X1 U67 ( .A(n14), .B(count[0]), .Y(n66) );
  AND2X2 U68 ( .A(count[0]), .B(n67), .Y(n65) );
  MUX2X1 U69 ( .B(n66), .A(n65), .S(count[1]), .Y(n71) );
  MUX2X1 U70 ( .B(n68), .A(n67), .S(count[0]), .Y(n69) );
endmodule


module tx_tcu_0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module tx_tcu_0 ( clk, rst, p_ready, t_bitstuff, PRGA_OUT, prga_opcode, t_crc, 
        sending, EOP, next_byte, send_data, t_strobe );
  input [7:0] PRGA_OUT;
  input [1:0] prga_opcode;
  input [15:0] t_crc;
  output [7:0] send_data;
  input clk, rst, p_ready, t_bitstuff;
  output sending, EOP, next_byte, t_strobe;
  wire   N59, N60, N61, N62, N63, N64, N65, N188, n1, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n175, n177, n179, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290;
  wire   [2:0] state;
  wire   [6:0] count;
  wire   [2:0] nextstate;
  wire   [7:0] flop_data;
  wire   [7:0] current_send_data;

  DFFSR \count_reg[0]  ( .D(n261), .CLK(clk), .R(n29), .S(1'b1), .Q(count[0])
         );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n29), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n29), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n29), .S(1'b1), .Q(
        state[2]) );
  DFFSR \count_reg[1]  ( .D(n267), .CLK(clk), .R(n29), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n266), .CLK(clk), .R(n29), .S(1'b1), .Q(count[2])
         );
  DFFSR \count_reg[4]  ( .D(n264), .CLK(clk), .R(n29), .S(1'b1), .Q(count[4])
         );
  DFFPOSX1 \flop_data_reg[7]  ( .D(n253), .CLK(clk), .Q(flop_data[7]) );
  DFFPOSX1 \current_send_data_reg[7]  ( .D(n275), .CLK(clk), .Q(
        current_send_data[7]) );
  DFFPOSX1 \flop_data_reg[6]  ( .D(n254), .CLK(clk), .Q(flop_data[6]) );
  DFFPOSX1 \current_send_data_reg[6]  ( .D(n276), .CLK(clk), .Q(
        current_send_data[6]) );
  DFFPOSX1 \flop_data_reg[5]  ( .D(n255), .CLK(clk), .Q(flop_data[5]) );
  DFFPOSX1 \current_send_data_reg[5]  ( .D(n277), .CLK(clk), .Q(
        current_send_data[5]) );
  DFFPOSX1 \flop_data_reg[4]  ( .D(n256), .CLK(clk), .Q(flop_data[4]) );
  DFFPOSX1 \current_send_data_reg[4]  ( .D(n278), .CLK(clk), .Q(
        current_send_data[4]) );
  DFFPOSX1 \flop_data_reg[3]  ( .D(n257), .CLK(clk), .Q(flop_data[3]) );
  DFFPOSX1 \current_send_data_reg[3]  ( .D(n279), .CLK(clk), .Q(
        current_send_data[3]) );
  DFFPOSX1 \flop_data_reg[2]  ( .D(n258), .CLK(clk), .Q(flop_data[2]) );
  DFFPOSX1 \current_send_data_reg[2]  ( .D(n280), .CLK(clk), .Q(
        current_send_data[2]) );
  DFFPOSX1 \flop_data_reg[1]  ( .D(n259), .CLK(clk), .Q(flop_data[1]) );
  DFFPOSX1 \current_send_data_reg[1]  ( .D(n281), .CLK(clk), .Q(
        current_send_data[1]) );
  DFFPOSX1 \flop_data_reg[0]  ( .D(n260), .CLK(clk), .Q(flop_data[0]) );
  DFFPOSX1 \current_send_data_reg[0]  ( .D(n282), .CLK(clk), .Q(
        current_send_data[0]) );
  DFFPOSX1 \send_data_reg[7]  ( .D(n283), .CLK(clk), .Q(send_data[7]) );
  DFFPOSX1 \send_data_reg[6]  ( .D(n284), .CLK(clk), .Q(send_data[6]) );
  DFFPOSX1 \send_data_reg[5]  ( .D(n285), .CLK(clk), .Q(send_data[5]) );
  DFFPOSX1 \send_data_reg[4]  ( .D(n286), .CLK(clk), .Q(send_data[4]) );
  DFFPOSX1 \send_data_reg[3]  ( .D(n287), .CLK(clk), .Q(send_data[3]) );
  DFFPOSX1 \send_data_reg[2]  ( .D(n288), .CLK(clk), .Q(send_data[2]) );
  DFFPOSX1 \send_data_reg[1]  ( .D(n289), .CLK(clk), .Q(send_data[1]) );
  DFFPOSX1 \send_data_reg[0]  ( .D(n290), .CLK(clk), .Q(send_data[0]) );
  tx_tcu_0_DW01_inc_0 r80 ( .A({n27, n7, n8, n9, n6, n13, count[0]}), .SUM({
        N65, N64, N63, N62, N61, N60, N59}) );
  DFFSR \count_reg[6]  ( .D(n262), .CLK(clk), .R(n29), .S(1'b1), .Q(N188) );
  DFFSR \count_reg[3]  ( .D(n265), .CLK(clk), .R(n29), .S(1'b1), .Q(count[3])
         );
  DFFSR \count_reg[5]  ( .D(n263), .CLK(clk), .R(n29), .S(1'b1), .Q(count[5])
         );
  INVX2 U3 ( .A(n11), .Y(n13) );
  INVX4 U4 ( .A(n28), .Y(n36) );
  INVX2 U5 ( .A(n187), .Y(n19) );
  INVX2 U6 ( .A(count[0]), .Y(n175) );
  NAND2X1 U7 ( .A(n14), .B(n112), .Y(n1) );
  INVX2 U11 ( .A(n125), .Y(n5) );
  INVX1 U12 ( .A(n191), .Y(n6) );
  INVX2 U13 ( .A(n154), .Y(n7) );
  BUFX4 U14 ( .A(count[4]), .Y(n8) );
  BUFX4 U15 ( .A(count[3]), .Y(n9) );
  INVX1 U16 ( .A(n147), .Y(n10) );
  INVX2 U17 ( .A(count[1]), .Y(n11) );
  INVX1 U18 ( .A(n11), .Y(n12) );
  INVX1 U19 ( .A(n20), .Y(n137) );
  AND2X2 U20 ( .A(n120), .B(n112), .Y(n15) );
  INVX2 U21 ( .A(n111), .Y(n14) );
  NAND2X1 U22 ( .A(n9), .B(count[0]), .Y(n16) );
  NAND2X1 U23 ( .A(n201), .B(n17), .Y(n192) );
  INVX2 U24 ( .A(n16), .Y(n17) );
  INVX2 U25 ( .A(count[3]), .Y(n190) );
  INVX1 U26 ( .A(n248), .Y(n62) );
  AND2X2 U27 ( .A(n132), .B(n94), .Y(n18) );
  INVX4 U28 ( .A(n18), .Y(n147) );
  INVX1 U29 ( .A(n109), .Y(n110) );
  OR2X2 U30 ( .A(n20), .B(n19), .Y(n140) );
  INVX2 U31 ( .A(n20), .Y(n186) );
  INVX1 U32 ( .A(n127), .Y(n138) );
  INVX1 U33 ( .A(n65), .Y(n34) );
  AND2X2 U34 ( .A(n6), .B(n24), .Y(n25) );
  OR2X2 U35 ( .A(n192), .B(n193), .Y(n20) );
  INVX1 U36 ( .A(n141), .Y(n90) );
  AND2X1 U37 ( .A(n13), .B(n22), .Y(n24) );
  INVX1 U38 ( .A(n93), .Y(n125) );
  INVX2 U39 ( .A(count[2]), .Y(n191) );
  INVX1 U40 ( .A(n140), .Y(n126) );
  AND2X1 U41 ( .A(n185), .B(n125), .Y(n21) );
  INVX2 U42 ( .A(rst), .Y(n29) );
  NOR2X1 U43 ( .A(t_bitstuff), .B(n175), .Y(n22) );
  BUFX4 U44 ( .A(N188), .Y(n27) );
  BUFX4 U45 ( .A(state[0]), .Y(n28) );
  AND2X2 U46 ( .A(state[2]), .B(n26), .Y(n23) );
  XOR2X1 U47 ( .A(n22), .B(n13), .Y(n116) );
  XOR2X1 U48 ( .A(n25), .B(n9), .Y(n99) );
  XOR2X1 U49 ( .A(n24), .B(n6), .Y(n105) );
  BUFX4 U50 ( .A(state[1]), .Y(n26) );
  INVX2 U51 ( .A(n27), .Y(n153) );
  INVX2 U52 ( .A(state[2]), .Y(n64) );
  INVX2 U53 ( .A(n26), .Y(n30) );
  NAND3X1 U54 ( .A(n28), .B(n64), .C(n30), .Y(n88) );
  NAND3X1 U55 ( .A(n26), .B(n64), .C(n36), .Y(n93) );
  NAND2X1 U56 ( .A(n88), .B(n93), .Y(n69) );
  NAND2X1 U57 ( .A(n69), .B(n29), .Y(n56) );
  NAND2X1 U58 ( .A(state[2]), .B(n30), .Y(n35) );
  NOR2X1 U59 ( .A(n36), .B(n35), .Y(n32) );
  INVX2 U60 ( .A(n222), .Y(n31) );
  NAND2X1 U61 ( .A(n32), .B(n31), .Y(n33) );
  OAI21X1 U62 ( .A(n189), .B(n56), .C(n33), .Y(n220) );
  NAND2X1 U63 ( .A(n23), .B(n36), .Y(n65) );
  NAND2X1 U64 ( .A(n34), .B(n29), .Y(n39) );
  INVX2 U65 ( .A(n35), .Y(n68) );
  NAND2X1 U66 ( .A(n68), .B(n36), .Y(n127) );
  NAND2X1 U67 ( .A(n138), .B(n29), .Y(n38) );
  INVX2 U68 ( .A(t_crc[15]), .Y(n37) );
  OAI22X1 U69 ( .A(n188), .B(n39), .C(n38), .D(n37), .Y(n221) );
  INVX2 U70 ( .A(n38), .Y(n53) );
  INVX2 U71 ( .A(n39), .Y(n52) );
  AOI22X1 U72 ( .A(t_crc[14]), .B(n53), .C(PRGA_OUT[6]), .D(n52), .Y(n225) );
  INVX2 U73 ( .A(flop_data[6]), .Y(n86) );
  NAND3X1 U74 ( .A(n245), .B(n28), .C(n68), .Y(n55) );
  INVX2 U75 ( .A(t_crc[6]), .Y(n40) );
  OAI22X1 U76 ( .A(n56), .B(n86), .C(n55), .D(n40), .Y(n41) );
  INVX2 U77 ( .A(n41), .Y(n226) );
  AOI22X1 U78 ( .A(t_crc[13]), .B(n53), .C(PRGA_OUT[5]), .D(n52), .Y(n228) );
  INVX2 U79 ( .A(flop_data[5]), .Y(n84) );
  INVX2 U80 ( .A(t_crc[5]), .Y(n42) );
  OAI22X1 U81 ( .A(n56), .B(n84), .C(n55), .D(n42), .Y(n43) );
  INVX2 U82 ( .A(n43), .Y(n229) );
  AOI22X1 U83 ( .A(t_crc[12]), .B(n53), .C(PRGA_OUT[4]), .D(n52), .Y(n231) );
  INVX2 U84 ( .A(flop_data[4]), .Y(n82) );
  INVX2 U85 ( .A(t_crc[4]), .Y(n44) );
  OAI22X1 U86 ( .A(n56), .B(n82), .C(n55), .D(n44), .Y(n45) );
  INVX2 U87 ( .A(n45), .Y(n232) );
  AOI22X1 U88 ( .A(t_crc[11]), .B(n53), .C(PRGA_OUT[3]), .D(n52), .Y(n234) );
  INVX2 U89 ( .A(flop_data[3]), .Y(n80) );
  INVX2 U90 ( .A(t_crc[3]), .Y(n46) );
  OAI22X1 U91 ( .A(n56), .B(n80), .C(n55), .D(n46), .Y(n47) );
  INVX2 U92 ( .A(n47), .Y(n235) );
  AOI22X1 U93 ( .A(t_crc[10]), .B(n53), .C(PRGA_OUT[2]), .D(n52), .Y(n237) );
  INVX2 U94 ( .A(flop_data[2]), .Y(n78) );
  INVX2 U95 ( .A(t_crc[2]), .Y(n48) );
  OAI22X1 U96 ( .A(n56), .B(n78), .C(n55), .D(n48), .Y(n49) );
  INVX2 U97 ( .A(n49), .Y(n238) );
  AOI22X1 U98 ( .A(t_crc[9]), .B(n53), .C(PRGA_OUT[1]), .D(n52), .Y(n240) );
  INVX2 U99 ( .A(flop_data[1]), .Y(n76) );
  INVX2 U100 ( .A(t_crc[1]), .Y(n50) );
  OAI22X1 U101 ( .A(n56), .B(n76), .C(n55), .D(n50), .Y(n51) );
  INVX2 U102 ( .A(n51), .Y(n241) );
  AOI22X1 U103 ( .A(t_crc[8]), .B(n53), .C(PRGA_OUT[0]), .D(n52), .Y(n243) );
  INVX2 U104 ( .A(flop_data[0]), .Y(n74) );
  INVX2 U105 ( .A(t_crc[0]), .Y(n54) );
  OAI22X1 U106 ( .A(n56), .B(n74), .C(n55), .D(n54), .Y(n57) );
  INVX2 U107 ( .A(n57), .Y(n244) );
  INVX2 U108 ( .A(count[4]), .Y(n155) );
  INVX2 U109 ( .A(count[5]), .Y(n154) );
  INVX2 U110 ( .A(n88), .Y(n139) );
  NAND2X1 U111 ( .A(n157), .B(n139), .Y(n58) );
  NOR2X1 U112 ( .A(n156), .B(n58), .Y(t_strobe) );
  NOR3X1 U113 ( .A(n26), .B(n28), .C(state[2]), .Y(n131) );
  INVX2 U114 ( .A(p_ready), .Y(n59) );
  NAND2X1 U115 ( .A(n131), .B(n59), .Y(n70) );
  OAI21X1 U116 ( .A(n187), .B(n5), .C(n70), .Y(n60) );
  AOI21X1 U117 ( .A(n23), .B(n28), .C(n60), .Y(n61) );
  INVX2 U118 ( .A(n61), .Y(next_byte) );
  NAND2X1 U119 ( .A(n247), .B(n27), .Y(n63) );
  NAND2X1 U120 ( .A(n68), .B(n62), .Y(n141) );
  OAI22X1 U121 ( .A(n63), .B(n141), .C(n185), .D(n93), .Y(EOP) );
  NAND2X1 U122 ( .A(n68), .B(n153), .Y(n67) );
  NAND3X1 U123 ( .A(n28), .B(n26), .C(n64), .Y(n92) );
  NAND2X1 U124 ( .A(n65), .B(n92), .Y(n142) );
  NOR2X1 U125 ( .A(n142), .B(n69), .Y(n66) );
  NAND3X1 U126 ( .A(n127), .B(n66), .C(n67), .Y(sending) );
  INVX2 U127 ( .A(PRGA_OUT[0]), .Y(n73) );
  NOR3X1 U128 ( .A(n69), .B(n23), .C(n68), .Y(n72) );
  AND2X2 U129 ( .A(n70), .B(n29), .Y(n71) );
  AND2X2 U130 ( .A(n72), .B(n71), .Y(n87) );
  MUX2X1 U131 ( .B(n74), .A(n73), .S(n87), .Y(n260) );
  INVX2 U132 ( .A(PRGA_OUT[1]), .Y(n75) );
  MUX2X1 U133 ( .B(n76), .A(n75), .S(n87), .Y(n259) );
  INVX2 U134 ( .A(PRGA_OUT[2]), .Y(n77) );
  MUX2X1 U135 ( .B(n78), .A(n77), .S(n87), .Y(n258) );
  INVX2 U136 ( .A(PRGA_OUT[3]), .Y(n79) );
  MUX2X1 U137 ( .B(n80), .A(n79), .S(n87), .Y(n257) );
  INVX2 U138 ( .A(PRGA_OUT[4]), .Y(n81) );
  MUX2X1 U139 ( .B(n82), .A(n81), .S(n87), .Y(n256) );
  INVX2 U140 ( .A(PRGA_OUT[5]), .Y(n83) );
  MUX2X1 U141 ( .B(n84), .A(n83), .S(n87), .Y(n255) );
  INVX2 U142 ( .A(PRGA_OUT[6]), .Y(n85) );
  MUX2X1 U143 ( .B(n86), .A(n85), .S(n87), .Y(n254) );
  MUX2X1 U144 ( .B(n189), .A(n188), .S(n87), .Y(n253) );
  OAI21X1 U145 ( .A(n186), .B(n127), .C(n88), .Y(n89) );
  NAND2X1 U146 ( .A(t_bitstuff), .B(n139), .Y(n100) );
  OAI21X1 U147 ( .A(n90), .B(n89), .C(n100), .Y(n91) );
  INVX2 U148 ( .A(n91), .Y(n146) );
  NAND2X1 U149 ( .A(N63), .B(n146), .Y(n98) );
  NAND2X1 U150 ( .A(n9), .B(n25), .Y(n109) );
  OR2X2 U151 ( .A(n186), .B(n92), .Y(n132) );
  NAND2X1 U152 ( .A(n125), .B(n140), .Y(n94) );
  NOR2X1 U153 ( .A(n109), .B(n10), .Y(n96) );
  NAND2X1 U154 ( .A(n109), .B(n147), .Y(n95) );
  NAND2X1 U155 ( .A(n100), .B(n95), .Y(n111) );
  MUX2X1 U156 ( .B(n96), .A(n111), .S(n8), .Y(n97) );
  NAND2X1 U157 ( .A(n98), .B(n97), .Y(n264) );
  NAND2X1 U158 ( .A(N62), .B(n146), .Y(n104) );
  NAND2X1 U159 ( .A(n99), .B(n147), .Y(n103) );
  INVX2 U160 ( .A(n100), .Y(n150) );
  INVX2 U161 ( .A(n190), .Y(n101) );
  NAND2X1 U162 ( .A(n150), .B(n101), .Y(n102) );
  NAND3X1 U163 ( .A(n104), .B(n103), .C(n102), .Y(n265) );
  NAND2X1 U164 ( .A(N61), .B(n146), .Y(n108) );
  NAND2X1 U165 ( .A(n105), .B(n147), .Y(n107) );
  NAND2X1 U166 ( .A(n150), .B(n6), .Y(n106) );
  NAND3X1 U167 ( .A(n108), .B(n107), .C(n106), .Y(n266) );
  NAND2X1 U168 ( .A(N64), .B(n146), .Y(n115) );
  NAND3X1 U169 ( .A(n110), .B(n8), .C(n147), .Y(n119) );
  INVX2 U170 ( .A(n119), .Y(n113) );
  NAND2X1 U171 ( .A(n147), .B(n155), .Y(n112) );
  MUX2X1 U172 ( .B(n113), .A(n1), .S(n7), .Y(n114) );
  NAND2X1 U173 ( .A(n115), .B(n114), .Y(n263) );
  AOI22X1 U174 ( .A(n116), .B(n147), .C(N60), .D(n146), .Y(n118) );
  NAND2X1 U175 ( .A(n150), .B(n13), .Y(n117) );
  NAND2X1 U176 ( .A(n118), .B(n117), .Y(n267) );
  NAND2X1 U177 ( .A(N65), .B(n146), .Y(n124) );
  NOR2X1 U178 ( .A(n154), .B(n119), .Y(n122) );
  NAND2X1 U179 ( .A(n147), .B(n154), .Y(n120) );
  NAND2X1 U180 ( .A(n15), .B(n14), .Y(n121) );
  MUX2X1 U181 ( .B(n122), .A(n121), .S(n27), .Y(n123) );
  NAND2X1 U182 ( .A(n124), .B(n123), .Y(n262) );
  NAND2X1 U183 ( .A(n177), .B(p_ready), .Y(n130) );
  NAND2X1 U184 ( .A(n126), .B(n21), .Y(n129) );
  AND2X2 U185 ( .A(n127), .B(n141), .Y(n128) );
  NAND3X1 U186 ( .A(n130), .B(n129), .C(n128), .Y(nextstate[2]) );
  NAND2X1 U187 ( .A(n131), .B(p_ready), .Y(n136) );
  NAND2X1 U188 ( .A(n21), .B(n140), .Y(n135) );
  INVX2 U189 ( .A(n132), .Y(n133) );
  AOI21X1 U190 ( .A(n179), .B(n139), .C(n133), .Y(n134) );
  NAND3X1 U191 ( .A(n136), .B(n135), .C(n134), .Y(nextstate[1]) );
  AOI22X1 U192 ( .A(n184), .B(n139), .C(n138), .D(n137), .Y(n145) );
  NAND3X1 U194 ( .A(n21), .B(n140), .C(p_ready), .Y(n144) );
  NOR2X1 U196 ( .A(n142), .B(n90), .Y(n143) );
  NAND3X1 U198 ( .A(n145), .B(n144), .C(n143), .Y(nextstate[0]) );
  XOR2X1 U203 ( .A(n175), .B(t_bitstuff), .Y(n148) );
  AOI22X1 U204 ( .A(n148), .B(n147), .C(N59), .D(n146), .Y(n152) );
  INVX2 U205 ( .A(n175), .Y(n149) );
  NAND2X1 U206 ( .A(n150), .B(n149), .Y(n151) );
  NAND2X1 U207 ( .A(n152), .B(n151), .Y(n261) );
  NAND2X1 U208 ( .A(n153), .B(n175), .Y(n156) );
  NOR2X1 U209 ( .A(n26), .B(n28), .Y(n177) );
  INVX1 U210 ( .A(n184), .Y(n179) );
  NAND3X1 U211 ( .A(n157), .B(n153), .C(count[0]), .Y(n184) );
  AND2X1 U212 ( .A(prga_opcode[1]), .B(prga_opcode[0]), .Y(n187) );
  NAND3X1 U213 ( .A(n8), .B(n13), .C(n7), .Y(n193) );
  NOR2X1 U214 ( .A(n27), .B(n191), .Y(n201) );
  OAI21X1 U215 ( .A(n202), .B(n203), .C(n204), .Y(n275) );
  INVX1 U216 ( .A(current_send_data[7]), .Y(n203) );
  OAI21X1 U217 ( .A(n202), .B(n205), .C(n206), .Y(n276) );
  INVX1 U218 ( .A(current_send_data[6]), .Y(n205) );
  OAI21X1 U219 ( .A(n202), .B(n207), .C(n208), .Y(n277) );
  INVX1 U220 ( .A(current_send_data[5]), .Y(n207) );
  OAI21X1 U221 ( .A(n202), .B(n209), .C(n210), .Y(n278) );
  INVX1 U222 ( .A(current_send_data[4]), .Y(n209) );
  OAI21X1 U223 ( .A(n202), .B(n211), .C(n212), .Y(n279) );
  INVX1 U224 ( .A(current_send_data[3]), .Y(n211) );
  OAI21X1 U225 ( .A(n202), .B(n213), .C(n214), .Y(n280) );
  INVX1 U226 ( .A(current_send_data[2]), .Y(n213) );
  OAI21X1 U227 ( .A(n202), .B(n215), .C(n216), .Y(n281) );
  INVX1 U228 ( .A(current_send_data[1]), .Y(n215) );
  OAI21X1 U229 ( .A(n202), .B(n217), .C(n218), .Y(n282) );
  INVX1 U230 ( .A(current_send_data[0]), .Y(n217) );
  AOI21X1 U231 ( .A(n28), .B(n26), .C(rst), .Y(n202) );
  NAND2X1 U232 ( .A(n219), .B(n204), .Y(n283) );
  NOR2X1 U233 ( .A(n220), .B(n221), .Y(n204) );
  INVX1 U234 ( .A(PRGA_OUT[7]), .Y(n188) );
  OAI21X1 U235 ( .A(n27), .B(t_crc[7]), .C(n29), .Y(n222) );
  INVX1 U236 ( .A(flop_data[7]), .Y(n189) );
  AOI22X1 U237 ( .A(n223), .B(current_send_data[7]), .C(send_data[7]), .D(rst), 
        .Y(n219) );
  NAND2X1 U238 ( .A(n224), .B(n206), .Y(n284) );
  AND2X1 U239 ( .A(n225), .B(n226), .Y(n206) );
  AOI22X1 U240 ( .A(n223), .B(current_send_data[6]), .C(send_data[6]), .D(rst), 
        .Y(n224) );
  NAND2X1 U241 ( .A(n227), .B(n208), .Y(n285) );
  AND2X1 U242 ( .A(n228), .B(n229), .Y(n208) );
  AOI22X1 U243 ( .A(n223), .B(current_send_data[5]), .C(send_data[5]), .D(rst), 
        .Y(n227) );
  NAND2X1 U244 ( .A(n230), .B(n210), .Y(n286) );
  AND2X1 U245 ( .A(n231), .B(n232), .Y(n210) );
  AOI22X1 U246 ( .A(n223), .B(current_send_data[4]), .C(send_data[4]), .D(rst), 
        .Y(n230) );
  NAND2X1 U247 ( .A(n233), .B(n212), .Y(n287) );
  AND2X1 U248 ( .A(n234), .B(n235), .Y(n212) );
  AOI22X1 U249 ( .A(n223), .B(current_send_data[3]), .C(send_data[3]), .D(rst), 
        .Y(n233) );
  NAND2X1 U250 ( .A(n236), .B(n214), .Y(n288) );
  AND2X1 U251 ( .A(n237), .B(n238), .Y(n214) );
  AOI22X1 U252 ( .A(n223), .B(current_send_data[2]), .C(send_data[2]), .D(rst), 
        .Y(n236) );
  NAND2X1 U253 ( .A(n239), .B(n216), .Y(n289) );
  AND2X1 U254 ( .A(n240), .B(n241), .Y(n216) );
  AOI22X1 U255 ( .A(n223), .B(current_send_data[1]), .C(send_data[1]), .D(rst), 
        .Y(n239) );
  NAND2X1 U256 ( .A(n242), .B(n218), .Y(n290) );
  AND2X1 U257 ( .A(n243), .B(n244), .Y(n218) );
  NOR2X1 U258 ( .A(rst), .B(n27), .Y(n245) );
  AOI22X1 U259 ( .A(n223), .B(current_send_data[0]), .C(send_data[0]), .D(rst), 
        .Y(n242) );
  INVX1 U260 ( .A(n246), .Y(n223) );
  NAND3X1 U261 ( .A(n28), .B(n29), .C(n26), .Y(n246) );
  OAI21X1 U262 ( .A(n249), .B(n250), .C(n28), .Y(n248) );
  NAND3X1 U263 ( .A(count[2]), .B(n27), .C(n9), .Y(n250) );
  NAND3X1 U264 ( .A(n155), .B(n154), .C(n251), .Y(n249) );
  NOR2X1 U265 ( .A(n12), .B(count[0]), .Y(n251) );
  NAND3X1 U266 ( .A(n157), .B(n175), .C(n27), .Y(n185) );
  NOR2X1 U267 ( .A(n247), .B(n13), .Y(n157) );
  NAND3X1 U268 ( .A(n191), .B(n190), .C(n252), .Y(n247) );
  NOR2X1 U269 ( .A(count[5]), .B(count[4]), .Y(n252) );
endmodule


module tx_timer_0 ( CLK, RST, SENDING, SHIFT_ENABLE_R, SHIFT_ENABLE_E );
  input CLK, RST, SENDING;
  output SHIFT_ENABLE_R, SHIFT_ENABLE_E;
  wire   state, nxt_SHIFT_ENABLE_E, n6, n8, n9, n10, n11, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28;
  wire   [3:0] count;
  wire   [3:0] nextcount;
  assign SHIFT_ENABLE_R = nxt_SHIFT_ENABLE_E;

  DFFSR state_reg ( .D(SENDING), .CLK(CLK), .R(n6), .S(1'b1), .Q(state) );
  DFFSR \count_reg[0]  ( .D(nextcount[0]), .CLK(CLK), .R(n6), .S(1'b1), .Q(
        count[0]) );
  DFFSR \count_reg[2]  ( .D(nextcount[2]), .CLK(CLK), .R(n6), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[1]  ( .D(nextcount[1]), .CLK(CLK), .R(n6), .S(1'b1), .Q(
        count[1]) );
  DFFSR \count_reg[3]  ( .D(nextcount[3]), .CLK(CLK), .R(n6), .S(1'b1), .Q(
        count[3]) );
  DFFSR SHIFT_ENABLE_E_reg ( .D(nxt_SHIFT_ENABLE_E), .CLK(CLK), .R(n6), .S(
        1'b1), .Q(SHIFT_ENABLE_E) );
  NOR2X1 U14 ( .A(n28), .B(n27), .Y(nextcount[3]) );
  XNOR2X1 U15 ( .A(count[3]), .B(n26), .Y(n28) );
  NOR2X1 U16 ( .A(n25), .B(n20), .Y(n26) );
  AOI21X1 U17 ( .A(n24), .B(state), .C(n21), .Y(nextcount[2]) );
  XNOR2X1 U18 ( .A(n25), .B(n20), .Y(n24) );
  NAND2X1 U19 ( .A(count[1]), .B(count[0]), .Y(n25) );
  NOR2X1 U20 ( .A(n23), .B(n27), .Y(nextcount[1]) );
  NAND3X1 U21 ( .A(SENDING), .B(n22), .C(state), .Y(n27) );
  XNOR2X1 U22 ( .A(count[0]), .B(count[1]), .Y(n23) );
  OAI21X1 U23 ( .A(count[0]), .B(n21), .C(state), .Y(nextcount[0]) );
  INVX1 U8 ( .A(SENDING), .Y(n21) );
  INVX2 U10 ( .A(RST), .Y(n6) );
  NOR2X1 U11 ( .A(count[0]), .B(count[2]), .Y(n9) );
  INVX2 U12 ( .A(count[1]), .Y(n8) );
  NAND2X1 U13 ( .A(n9), .B(n8), .Y(n22) );
  INVX2 U24 ( .A(n22), .Y(n11) );
  AND2X2 U25 ( .A(count[3]), .B(state), .Y(n10) );
  NAND3X1 U26 ( .A(SENDING), .B(n11), .C(n10), .Y(n19) );
  INVX2 U27 ( .A(n19), .Y(nxt_SHIFT_ENABLE_E) );
  INVX2 U28 ( .A(count[2]), .Y(n20) );
endmodule


module transmitter_block_0 ( PRGA_OUT, clk, p_ready, prga_opcode, rst, SENDING, 
        dm_tx_out, dp_tx_out, NEXT_BYTE );
  input [7:0] PRGA_OUT;
  input [1:0] prga_opcode;
  input clk, p_ready, rst;
  output SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE;
  wire   t_strobe, EOP, SHIFT_ENABLE_E, d_encode, t_bitstuff, SHIFT_ENABLE_R;
  wire   [15:0] TX_CRC;
  wire   [7:0] send_data;

  tx_CRC_CALC_0 U_1 ( .CLK(clk), .RST(rst), .EOP(EOP), .T_STROBE(t_strobe), 
        .PRGA_OPCODE(prga_opcode), .PRGA_OUT(PRGA_OUT), .TX_CRC(TX_CRC) );
  tx_encode_0 U_0 ( .clk(clk), .rst(rst), .SHIFT_ENABLE_E(SHIFT_ENABLE_E), 
        .d_encode(d_encode), .EOP(EOP), .t_bitstuff(t_bitstuff), .dp_tx_out(
        dp_tx_out), .dm_tx_out(dm_tx_out) );
  tx_shiftreg_0 U_2 ( .clk(clk), .rst(rst), .SHIFT_ENABLE_R(SHIFT_ENABLE_R), 
        .t_bitstuff(t_bitstuff), .t_strobe(t_strobe), .send_data(send_data), 
        .d_encode(d_encode) );
  tx_tcu_0 U_3 ( .clk(clk), .rst(rst), .p_ready(p_ready), .t_bitstuff(
        t_bitstuff), .PRGA_OUT(PRGA_OUT), .prga_opcode(prga_opcode), .t_crc(
        TX_CRC), .sending(SENDING), .EOP(EOP), .next_byte(NEXT_BYTE), 
        .send_data(send_data), .t_strobe(t_strobe) );
  tx_timer_0 U_4 ( .CLK(clk), .RST(rst), .SENDING(SENDING), .SHIFT_ENABLE_R(
        SHIFT_ENABLE_R), .SHIFT_ENABLE_E(SHIFT_ENABLE_E) );
endmodule


module RMEDT_REWIRE_0 ( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN, DATA_IN, BS_ERROR, 
        CRC_ERROR, EMPTY, FULL, KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, 
        R_ERROR, SENDING, dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE, DATA, 
        ADDR );
  input [7:0] DATA_IN;
  output [7:0] DATA;
  output [7:0] ADDR;
  input CLK, DM1_RX, DP1_RX, RST, SERIAL_IN;
  output BS_ERROR, CRC_ERROR, EMPTY, FULL, KEY_ERROR, PROG_ERROR, PARITY_ERROR,
         RBUF_FULL, R_ERROR, SENDING, dm_tx_out, dp_tx_out, W_ENABLE_R,
         R_ENABLE;
  wire   B_READY, PDATA_READY, EOP_external, NEXT_BYTE, W_ENABLE;
  wire   [7:0] PRGA_IN;
  wire   [1:0] PRGA_OPCODE;
  wire   [7:0] PROCESSED_DATA;
  wire   [7:0] RCV_DATA;
  wire   [1:0] OPCODE;

  EDBlock_0 U_0 ( .BYTE(PRGA_IN), .BYTE_READY(B_READY), .CLK(CLK), .OPCODE(
        PRGA_OPCODE), .RST(RST), .SERIAL_IN(SERIAL_IN), .DATA_IN(DATA_IN), 
        .KEY_ERROR(KEY_ERROR), .PARITY_ERROR(PARITY_ERROR), .PDATA_READY(
        PDATA_READY), .PROCESSED_DATA(PROCESSED_DATA), .PROG_ERROR(PROG_ERROR), 
        .RBUF_FULL(RBUF_FULL), .W_ENABLE(W_ENABLE_R), .R_ENABLE(R_ENABLE), 
        .DATA(DATA), .ADDR(ADDR) );
  memoryblock_0 U_1 ( .CLK(CLK), .NEXT_BYTE(NEXT_BYTE), .RCV_DATA(RCV_DATA), 
        .RCV_OPCODE(OPCODE), .RST(RST), .W_ENABLE(W_ENABLE), .EOP(EOP_external), .EMPTY(EMPTY), .FULL(FULL), .B_READY(B_READY), .PRGA_IN(PRGA_IN), 
        .PRGA_OPCODE(PRGA_OPCODE) );
  receiver_block_rewire_0 U_2 ( .CLK(CLK), .DM1_RX(DM1_RX), .DP1_RX(DP1_RX), 
        .RST(RST), .BS_ERROR(BS_ERROR), .CRC_ERROR(CRC_ERROR), .EOP_external(
        EOP_external), .OPCODE(OPCODE), .RCV_DATA(RCV_DATA), .R_ERROR(R_ERROR), 
        .W_ENABLE(W_ENABLE) );
  transmitter_block_0 U_3 ( .PRGA_OUT(PROCESSED_DATA), .clk(CLK), .p_ready(
        PDATA_READY), .prga_opcode(PRGA_OPCODE), .rst(RST), .SENDING(SENDING), 
        .dm_tx_out(dm_tx_out), .dp_tx_out(dp_tx_out), .NEXT_BYTE(NEXT_BYTE) );
endmodule


module rmedt_square_t ( CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN, DATA_IN_H, 
        DATA_IN_S, BSE_H, BSE_S, CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, 
        EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, 
        c_parity_error, c_prog_error, host_is_sending, slave_is_sending, 
        W_ENABLE_H, W_ENABLE_S, R_ENABLE_H, R_ENABLE_S, DATA_H, DATA_S, ADDR_H, 
        ADDR_S );
  input [7:0] DATA_IN_H;
  input [7:0] DATA_IN_S;
  output [7:0] DATA_H;
  output [7:0] DATA_S;
  output [7:0] ADDR_H;
  output [7:0] ADDR_S;
  input CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN;
  output BSE_H, BSE_S, CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, EMPTY_H,
         EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, c_parity_error,
         c_prog_error, host_is_sending, slave_is_sending, W_ENABLE_H,
         W_ENABLE_S, R_ENABLE_H, R_ENABLE_S;
  wire   KEY_ERROR, KEY_ERROR1, PARITY_ERROR, PARITY_ERROR1, PROG_ERROR,
         PROG_ERROR1;

  OR2X2 U1 ( .A(PROG_ERROR), .B(PROG_ERROR1), .Y(c_prog_error) );
  OR2X2 U2 ( .A(PARITY_ERROR), .B(PARITY_ERROR1), .Y(c_parity_error) );
  OR2X2 U3 ( .A(KEY_ERROR), .B(KEY_ERROR1), .Y(c_key_error) );
  RMEDT_REWIRE_1 U_0 ( .CLK(CLK), .DM1_RX(DMRH), .DP1_RX(DPRH), .RST(RST), 
        .SERIAL_IN(SERIAL_IN), .DATA_IN(DATA_IN_H), .BS_ERROR(BSE_H), 
        .CRC_ERROR(CRCE_H), .EMPTY(EMPTY_H), .FULL(FULL_H), .KEY_ERROR(
        KEY_ERROR), .PROG_ERROR(PROG_ERROR), .PARITY_ERROR(PARITY_ERROR), 
        .R_ERROR(RE_H), .SENDING(host_is_sending), .dm_tx_out(DMTS), 
        .dp_tx_out(DPTS), .W_ENABLE_R(W_ENABLE_H), .R_ENABLE(R_ENABLE_H), 
        .DATA(DATA_H), .ADDR(ADDR_H) );
  RMEDT_REWIRE_0 U_1 ( .CLK(CLK), .DM1_RX(DMRS), .DP1_RX(DPRS), .RST(RST), 
        .SERIAL_IN(SERIAL_IN), .DATA_IN(DATA_IN_S), .BS_ERROR(BSE_S), 
        .CRC_ERROR(CRCE_S), .EMPTY(EMPTY_S), .FULL(FULL_S), .KEY_ERROR(
        KEY_ERROR1), .PROG_ERROR(PROG_ERROR1), .PARITY_ERROR(PARITY_ERROR1), 
        .R_ERROR(RE_S), .SENDING(slave_is_sending), .dm_tx_out(DMTH), 
        .dp_tx_out(DPTH), .W_ENABLE_R(W_ENABLE_S), .R_ENABLE(R_ENABLE_S), 
        .DATA(DATA_S), .ADDR(ADDR_S) );
endmodule

module  rmedt_square ( CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN, BSE_H, BSE_S, 
	CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, DPHS, DMHS, DPSS, DMSS, EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, 
	RE_S, c_key_error, c_parity_error, c_prog_error, host_is_sending, slave_is_sending );

input   CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN;
output  BSE_H, BSE_S, CRCE_H, CRCE_S, EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, c_parity_error, c_prog_error, DMTH, DMTS, DPTH, DPTS, slave_is_sending, host_is_sending;
inout   DPHS, DMHS, DPSS, DMSS;
wire	nCLK, nDMRH, nDMRS, nDPRH, nDPRS, nRST, nSERIAL_IN, nBSE_H, nBSE_S, nCRCE_H, nCRCE_S, nDMTH, nDMTS, nDPTH, nDPTS, nEMPTY_H, nEMPTY_S, nFULL_H, nFULL_S, nRE_H, nRE_S, nc_key_error, nc_parity_error, nc_prog_error, nhost_is_sending, nslave_is_sending;

        rmedt_square_t I0 ( .CLK(nCLK), .DMRH(nDMRH), .DMRS(nDMRS), .DPRH(nDPRH), 
	.DPRS(nDPRS), .RST(nRST), .SERIAL_IN(nSERIAL_IN), .BSE_H(nBSE_H), .BSE_S(nBSE_S), 
	.CRCE_H(nCRCE_H), .CRCE_S(nCRCE_S), .DMTH(nDMTH), .DMTS(nDMTS), 
	.DPTH(nDPTH), .DPTS(nDPTS), .EMPTY_H(nEMPTY_H), .EMPTY_S(nSERIAL_IN), 
	.FULL_H(nFULL_H), .FULL_S(nFULL_S), .RE_H(nRE_H), .RE_S(nRE_S), 
	.c_key_error(nc_key_error), .c_parity_error(nc_parity_error), .c_prog_error(nc_prog_error), .host_is_sending(nhost_is_sending), 
	.slave_is_sending(nslave_is_sending));

PADVDD UVDD (  );
PADGND UGND (  );
PADINC UCLK ( .DI(nCLK), .YPAD(CLK) );
PADINC URST ( .DI(nRST), .YPAD(RST) );
PADINC U_SERIAL_IN ( .DI(nSERIAL_IN), .YPAD(SERIAL_IN) );
PADINOUT U_HOST_PLUS ( .DI(nDPRH), .DO(nDPTH), .OEN(nslave_is_sending), .YPAD(DPHS));
PADINOUT U_HOST_MINUS( .DI(nDMRH), .DO(nDMTH), .OEN(nslave_is_sending), .YPAD(DMHS));
PADINOUT U_SLAVE_PLUS ( .DI(nDPRS), .DO(nDPTS), .OEN(nhost_is_sending), .YPAD(DPSS));
PADINOUT U_SLAVE_MINUS ( .DI(nDMRS), .DO(nDMTS), .OEN(nhost_is_sending), .YPAD(DMSS));
//PADOUT U_BSE_H ( .DO(BSE_H), .YPAD(nBSE_H) );
//PADOUT U_BSE_S ( .DO(BSE_S), .YPAD(nBSE_S) );
PADOUT U_CRCE_H ( .DO(CRCE_H), .YPAD(nCRCE_H) );
PADOUT U_CRCE_S ( .DO(CRCE_S), .YPAD(nCRCE_S) );
PADOUT U_EMPTY_H ( .DO(EMPTY_H), .YPAD(nEMPTY_H) );
PADOUT U_EMPTY_S ( .DO(EMPTY_S), .YPAD(nEMPTY_S) );
PADOUT U_FULL_H ( .DO(FULL_H), .YPAD(nFULL_H) );
PADOUT U_FULL_S ( .DO(FULL_S), .YPAD(nFULL_S) );
PADOUT U_RE_H ( .DO(RE_H), .YPAD(nRE_H) );
PADOUT U_RE_S ( .DO(RE_S), .YPAD(nRE_S) );
PADOUT U_KEY ( .DO(c_key_error), .YPAD(nc_key_error) );
PADOUT U_PARITY ( .DO(c_parity_error), .YPAD(nc_parity_error) );
PADOUT U_PROG ( .DO(c_prog_error), .YPAD(nc_prog_error) );

endmodule
