
module rmedt_square_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module rmedt_square_DW01_add_2 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_add_3 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module rmedt_square_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module rmedt_square_DW01_inc_5 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module rmedt_square_DW01_add_6 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_add_7 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_inc_6 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module rmedt_square_DW01_inc_7 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module rmedt_square_DW01_inc_8 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module rmedt_square_DW01_add_9 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_inc_10 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module rmedt_square_DW01_inc_11 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module rmedt_square_DW01_add_11 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_inc_13 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module rmedt_square_DW01_add_15 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_add_14 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_add_13 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_DW01_add_12 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module rmedt_square_t ( CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN, DATA_IN_H, 
        DATA_IN_S, BSE_H, BSE_S, CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, 
        EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, 
        c_parity_error, c_prog_error, host_is_sending, slave_is_sending, 
        W_ENABLE_H, W_ENABLE_S, R_ENABLE_H, R_ENABLE_S, DATA_H, DATA_S, ADDR_H, 
        ADDR_S );
  input [7:0] DATA_IN_H;
  input [7:0] DATA_IN_S;
  output [7:0] DATA_H;
  output [7:0] DATA_S;
  output [7:0] ADDR_H;
  output [7:0] ADDR_S;
  input CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN;
  output BSE_H, BSE_S, CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, EMPTY_H,
         EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, c_parity_error,
         c_prog_error, host_is_sending, slave_is_sending, W_ENABLE_H,
         W_ENABLE_S, R_ENABLE_H, R_ENABLE_S;
  wire   PARITY_ERROR, PARITY_ERROR1, \U_0/PDATA_READY , \U_0/PRGA_OPCODE[0] ,
         \U_0/PRGA_OPCODE[1] , \U_0/B_READY , \U_0/RBUF_FULL ,
         \U_0/U_0/U_0/N527 , \U_0/U_0/U_0/N526 , \U_0/U_0/U_0/N525 ,
         \U_0/U_0/U_0/N524 , \U_0/U_0/U_0/N523 , \U_0/U_0/U_0/N522 ,
         \U_0/U_0/U_0/N521 , \U_0/U_0/U_0/N520 , \U_0/U_0/U_0/N519 ,
         \U_0/U_0/U_0/N518 , \U_0/U_0/U_0/N517 , \U_0/U_0/U_0/N516 ,
         \U_0/U_0/U_0/N515 , \U_0/U_0/U_0/N514 , \U_0/U_0/U_0/N513 ,
         \U_0/U_0/U_0/N512 , \U_0/U_0/U_0/N503 , \U_0/U_0/U_0/N502 ,
         \U_0/U_0/U_0/N501 , \U_0/U_0/U_0/N500 , \U_0/U_0/U_0/N499 ,
         \U_0/U_0/U_0/N498 , \U_0/U_0/U_0/N497 , \U_0/U_0/U_0/N496 ,
         \U_0/U_0/U_0/N487 , \U_0/U_0/U_0/N486 , \U_0/U_0/U_0/N485 ,
         \U_0/U_0/U_0/N484 , \U_0/U_0/U_0/N483 , \U_0/U_0/U_0/N482 ,
         \U_0/U_0/U_0/N481 , \U_0/U_0/U_0/N480 , \U_0/U_0/U_0/N479 ,
         \U_0/U_0/U_0/N478 , \U_0/U_0/U_0/N477 , \U_0/U_0/U_0/N476 ,
         \U_0/U_0/U_0/N475 , \U_0/U_0/U_0/N474 , \U_0/U_0/U_0/N473 ,
         \U_0/U_0/U_0/N472 , \U_0/U_0/U_0/N448 , \U_0/U_0/U_0/N447 ,
         \U_0/U_0/U_0/N446 , \U_0/U_0/U_0/N445 , \U_0/U_0/U_0/N444 ,
         \U_0/U_0/U_0/N443 , \U_0/U_0/U_0/N442 , \U_0/U_0/U_0/N431 ,
         \U_0/U_0/U_0/N430 , \U_0/U_0/U_0/N429 , \U_0/U_0/U_0/N428 ,
         \U_0/U_0/U_0/N427 , \U_0/U_0/U_0/N426 , \U_0/U_0/U_0/N425 ,
         \U_0/U_0/U_0/N424 , \U_0/U_0/U_0/N414 , \U_0/U_0/U_0/N413 ,
         \U_0/U_0/U_0/N412 , \U_0/U_0/U_0/N411 , \U_0/U_0/U_0/N410 ,
         \U_0/U_0/U_0/N409 , \U_0/U_0/U_0/N408 , \U_0/U_0/U_0/N407 ,
         \U_0/U_0/U_0/fr_enable , \U_0/U_0/U_0/fw_enable ,
         \U_0/U_0/U_0/prefillCounter[0] , \U_0/U_0/U_0/prefillCounter[1] ,
         \U_0/U_0/U_0/prefillCounter[2] , \U_0/U_0/U_0/prefillCounter[3] ,
         \U_0/U_0/U_0/prefillCounter[4] , \U_0/U_0/U_0/prefillCounter[5] ,
         \U_0/U_0/U_0/prefillCounter[6] , \U_0/U_0/U_0/prefillCounter[7] ,
         \U_0/U_0/U_0/keyTable[0][7] , \U_0/U_0/U_0/keyTable[0][6] ,
         \U_0/U_0/U_0/keyTable[0][5] , \U_0/U_0/U_0/keyTable[0][4] ,
         \U_0/U_0/U_0/keyTable[0][3] , \U_0/U_0/U_0/keyTable[0][2] ,
         \U_0/U_0/U_0/keyTable[0][1] , \U_0/U_0/U_0/keyTable[0][0] ,
         \U_0/U_0/U_0/keyTable[1][7] , \U_0/U_0/U_0/keyTable[1][6] ,
         \U_0/U_0/U_0/keyTable[1][5] , \U_0/U_0/U_0/keyTable[1][4] ,
         \U_0/U_0/U_0/keyTable[1][3] , \U_0/U_0/U_0/keyTable[1][2] ,
         \U_0/U_0/U_0/keyTable[1][1] , \U_0/U_0/U_0/keyTable[1][0] ,
         \U_0/U_0/U_0/keyTable[2][7] , \U_0/U_0/U_0/keyTable[2][6] ,
         \U_0/U_0/U_0/keyTable[2][5] , \U_0/U_0/U_0/keyTable[2][4] ,
         \U_0/U_0/U_0/keyTable[2][3] , \U_0/U_0/U_0/keyTable[2][2] ,
         \U_0/U_0/U_0/keyTable[2][1] , \U_0/U_0/U_0/keyTable[2][0] ,
         \U_0/U_0/U_0/keyTable[3][7] , \U_0/U_0/U_0/keyTable[3][6] ,
         \U_0/U_0/U_0/keyTable[3][5] , \U_0/U_0/U_0/keyTable[3][4] ,
         \U_0/U_0/U_0/keyTable[3][3] , \U_0/U_0/U_0/keyTable[3][2] ,
         \U_0/U_0/U_0/keyTable[3][1] , \U_0/U_0/U_0/keyTable[3][0] ,
         \U_0/U_0/U_0/keyTable[4][7] , \U_0/U_0/U_0/keyTable[4][6] ,
         \U_0/U_0/U_0/keyTable[4][5] , \U_0/U_0/U_0/keyTable[4][4] ,
         \U_0/U_0/U_0/keyTable[4][3] , \U_0/U_0/U_0/keyTable[4][2] ,
         \U_0/U_0/U_0/keyTable[4][1] , \U_0/U_0/U_0/keyTable[4][0] ,
         \U_0/U_0/U_0/keyTable[5][7] , \U_0/U_0/U_0/keyTable[5][6] ,
         \U_0/U_0/U_0/keyTable[5][5] , \U_0/U_0/U_0/keyTable[5][4] ,
         \U_0/U_0/U_0/keyTable[5][3] , \U_0/U_0/U_0/keyTable[5][2] ,
         \U_0/U_0/U_0/keyTable[5][1] , \U_0/U_0/U_0/keyTable[5][0] ,
         \U_0/U_0/U_0/keyTable[6][7] , \U_0/U_0/U_0/keyTable[6][6] ,
         \U_0/U_0/U_0/keyTable[6][5] , \U_0/U_0/U_0/keyTable[6][4] ,
         \U_0/U_0/U_0/keyTable[6][3] , \U_0/U_0/U_0/keyTable[6][2] ,
         \U_0/U_0/U_0/keyTable[6][1] , \U_0/U_0/U_0/keyTable[6][0] ,
         \U_0/U_0/U_0/keyTable[7][7] , \U_0/U_0/U_0/keyTable[7][6] ,
         \U_0/U_0/U_0/keyTable[7][5] , \U_0/U_0/U_0/keyTable[7][4] ,
         \U_0/U_0/U_0/keyTable[7][3] , \U_0/U_0/U_0/keyTable[7][2] ,
         \U_0/U_0/U_0/keyTable[7][1] , \U_0/U_0/U_0/keyTable[7][0] ,
         \U_0/U_0/U_0/nextProcessedData[0] ,
         \U_0/U_0/U_0/nextProcessedData[1] ,
         \U_0/U_0/U_0/nextProcessedData[2] ,
         \U_0/U_0/U_0/nextProcessedData[3] ,
         \U_0/U_0/U_0/nextProcessedData[4] ,
         \U_0/U_0/U_0/nextProcessedData[5] ,
         \U_0/U_0/U_0/nextProcessedData[6] ,
         \U_0/U_0/U_0/nextProcessedData[7] , \U_0/U_0/U_0/extratemp[0] ,
         \U_0/U_0/U_0/extratemp[1] , \U_0/U_0/U_0/extratemp[2] ,
         \U_0/U_0/U_0/extratemp[3] , \U_0/U_0/U_0/extratemp[4] ,
         \U_0/U_0/U_0/extratemp[5] , \U_0/U_0/U_0/extratemp[6] ,
         \U_0/U_0/U_0/extratemp[7] , \U_0/U_0/U_0/temp[0] ,
         \U_0/U_0/U_0/temp[1] , \U_0/U_0/U_0/temp[2] , \U_0/U_0/U_0/temp[3] ,
         \U_0/U_0/U_0/temp[4] , \U_0/U_0/U_0/temp[5] , \U_0/U_0/U_0/temp[6] ,
         \U_0/U_0/U_0/temp[7] , \U_0/U_0/U_0/permuteComplete ,
         \U_0/U_0/U_0/keyi[0] , \U_0/U_0/U_0/keyi[1] , \U_0/U_0/U_0/keyi[2] ,
         \U_0/U_0/U_0/intj[0] , \U_0/U_0/U_0/intj[1] , \U_0/U_0/U_0/intj[2] ,
         \U_0/U_0/U_0/intj[3] , \U_0/U_0/U_0/intj[4] , \U_0/U_0/U_0/intj[5] ,
         \U_0/U_0/U_0/intj[6] , \U_0/U_0/U_0/intj[7] , \U_0/U_0/U_0/inti[0] ,
         \U_0/U_0/U_0/inti[1] , \U_0/U_0/U_0/inti[2] , \U_0/U_0/U_0/inti[3] ,
         \U_0/U_0/U_0/inti[4] , \U_0/U_0/U_0/inti[5] , \U_0/U_0/U_0/inti[6] ,
         \U_0/U_0/U_0/inti[7] , \U_0/U_0/U_0/sj[0] , \U_0/U_0/U_0/sj[1] ,
         \U_0/U_0/U_0/sj[2] , \U_0/U_0/U_0/sj[3] , \U_0/U_0/U_0/sj[4] ,
         \U_0/U_0/U_0/sj[5] , \U_0/U_0/U_0/sj[6] , \U_0/U_0/U_0/sj[7] ,
         \U_0/U_0/U_0/si[0] , \U_0/U_0/U_0/si[1] , \U_0/U_0/U_0/si[2] ,
         \U_0/U_0/U_0/si[3] , \U_0/U_0/U_0/si[4] , \U_0/U_0/U_0/si[5] ,
         \U_0/U_0/U_0/si[6] , \U_0/U_0/U_0/si[7] , \U_0/U_0/U_0/state[0] ,
         \U_0/U_0/U_0/state[1] , \U_0/U_0/U_0/state[2] ,
         \U_0/U_0/U_0/state[3] , \U_0/U_0/U_0/state[4] , \U_0/U_0/U_1/SBE ,
         \U_0/U_0/U_1/TIMER_TRIG , \U_0/U_0/U_1/SET_RBUF_FULL ,
         \U_0/U_0/U_1/SBC_EN , \U_0/U_0/U_1/SBC_CLR , \U_0/U_0/U_1/RBUF_LOAD ,
         \U_0/U_0/U_1/SB_DETECT , \U_0/U_0/U_1/OE , \U_0/U_0/U_1/CHK_ERROR ,
         \U_0/U_0/U_1/U_0/Q_int2 , \U_0/U_0/U_1/U_0/Q_int ,
         \U_0/U_0/U_1/U_1/OE_prime , \U_0/U_0/U_1/U_2/N99 ,
         \U_0/U_0/U_1/U_2/N38 , \U_0/U_0/U_1/U_2/N37 , \U_0/U_0/U_1/U_2/N36 ,
         \U_0/U_0/U_1/U_2/N35 , \U_0/U_0/U_1/U_2/N34 , \U_0/U_0/U_1/U_2/N33 ,
         \U_0/U_0/U_1/U_2/N32 , \U_0/U_0/U_1/U_2/N31 , \U_0/U_0/U_1/U_2/N30 ,
         \U_0/U_0/U_1/U_2/N29 , \U_0/U_0/U_1/U_2/N28 , \U_0/U_0/U_1/U_2/N27 ,
         \U_0/U_0/U_1/U_2/N26 , \U_0/U_0/U_1/U_2/N25 , \U_0/U_0/U_1/U_2/N24 ,
         \U_0/U_0/U_1/U_2/N23 , \U_0/U_0/U_1/U_2/nextState[0] ,
         \U_0/U_0/U_1/U_2/nextState[1] , \U_0/U_0/U_1/U_2/nextState[2] ,
         \U_0/U_0/U_1/U_2/count[1] , \U_0/U_0/U_1/U_2/count[2] ,
         \U_0/U_0/U_1/U_2/count[3] , \U_0/U_0/U_1/U_2/count[4] ,
         \U_0/U_0/U_1/U_2/count[5] , \U_0/U_0/U_1/U_2/count[6] ,
         \U_0/U_0/U_1/U_2/count[7] , \U_0/U_0/U_1/U_2/timerRunning ,
         \U_0/U_0/U_1/U_2/state[0] , \U_0/U_0/U_1/U_2/state[1] ,
         \U_0/U_0/U_1/U_2/state[2] , \U_0/U_0/U_1/U_5/sb_detect_flag ,
         \U_0/U_0/U_1/U_5/SBE_prime , \U_0/U_0/U_1/U_8/N1799 ,
         \U_0/U_0/U_1/U_8/N1798 , \U_0/U_0/U_1/U_8/N1797 ,
         \U_0/U_0/U_1/U_8/N1796 , \U_0/U_0/U_1/U_8/N1795 ,
         \U_0/U_0/U_1/U_8/N1794 , \U_0/U_0/U_1/U_8/N1793 ,
         \U_0/U_0/U_1/U_8/N1792 , \U_0/U_0/U_1/U_8/nextParityError ,
         \U_0/U_0/U_1/U_8/parityAccumulator[0] ,
         \U_0/U_0/U_1/U_8/parityAccumulator[1] ,
         \U_0/U_0/U_1/U_8/parityAccumulator[2] ,
         \U_0/U_0/U_1/U_8/parityAccumulator[3] ,
         \U_0/U_0/U_1/U_8/parityAccumulator[4] ,
         \U_0/U_0/U_1/U_8/parityAccumulator[5] ,
         \U_0/U_0/U_1/U_8/parityAccumulator[6] ,
         \U_0/U_0/U_1/U_8/parityAccumulator[7] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[0] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[1] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[2] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[3] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[4] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[5] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[6] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[7] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[8] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[9] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[10] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[11] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[12] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[13] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[14] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[15] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[16] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[17] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[18] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[19] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[20] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[21] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[22] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[23] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[24] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[25] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[26] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[27] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[28] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[29] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[30] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[31] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[32] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[33] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[34] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[35] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[36] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[37] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[38] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[39] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[40] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[41] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[42] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[43] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[44] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[45] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[46] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[47] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[48] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[49] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[50] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[51] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[52] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[53] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[54] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[55] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[56] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[57] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[58] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[59] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[60] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[61] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[62] ,
         \U_0/U_0/U_1/U_8/currentPlainKey[63] , \U_0/U_0/U_1/U_8/address[0] ,
         \U_0/U_0/U_1/U_8/address[1] , \U_0/U_0/U_1/U_8/address[2] ,
         \U_0/U_0/U_1/U_8/address[3] , \U_0/U_0/U_1/U_8/address[4] ,
         \U_0/U_0/U_1/U_8/address[5] , \U_0/U_0/U_1/U_8/address[6] ,
         \U_0/U_0/U_1/U_8/address[7] , \U_0/U_0/U_1/U_8/keyCount[0] ,
         \U_0/U_0/U_1/U_8/keyCount[1] , \U_0/U_0/U_1/U_8/keyCount[2] ,
         \U_0/U_0/U_1/U_8/keyCount[3] , \U_0/U_0/U_1/U_8/parityError ,
         \U_0/U_0/U_1/U_8/state[0] , \U_0/U_0/U_1/U_8/state[1] ,
         \U_0/U_0/U_1/U_8/state[2] , \U_0/U_0/U_1/U_8/state[3] ,
         \U_0/U_0/U_1/U_7/N33 , \U_0/U_0/U_1/U_7/N32 , \U_0/U_0/U_1/U_7/N31 ,
         \U_0/U_0/U_1/U_7/N30 , \U_0/U_0/U_1/U_7/N29 , \U_0/U_0/U_1/U_7/N28 ,
         \U_0/U_0/U_1/U_7/N27 , \U_0/U_0/U_1/U_7/N26 ,
         \U_0/U_0/U_1/U_7/nextState[0] , \U_0/U_0/U_1/U_7/nextState[1] ,
         \U_0/U_0/U_1/U_7/nextState[2] , \U_0/U_0/U_1/U_7/nextState[3] ,
         \U_0/U_0/U_1/U_7/nextState[4] , \U_0/U_0/U_1/U_7/nextState[5] ,
         \U_0/U_0/U_1/U_7/nextState[6] , \U_0/U_0/U_1/U_7/nextState[7] ,
         \U_0/U_0/U_1/U_7/state[0] , \U_0/U_0/U_1/U_7/state[1] ,
         \U_0/U_0/U_1/U_7/state[2] , \U_0/U_0/U_1/U_7/state[3] ,
         \U_0/U_0/U_1/U_7/state[4] , \U_0/U_0/U_1/U_7/state[5] ,
         \U_0/U_0/U_1/U_7/state[6] , \U_0/U_0/U_1/U_7/state[7] ,
         \U_0/U_1/R_ENABLE , \U_0/U_1/U_0/N40 , \U_0/U_1/U_0/N39 ,
         \U_0/U_1/U_0/state[0] , \U_0/U_1/U_0/state[1] ,
         \U_0/U_1/U_0/state[2] , \U_0/U_1/U_1/N355 , \U_0/U_1/U_1/N349 ,
         \U_0/U_1/U_1/N347 , \U_0/U_1/U_1/N346 , \U_0/U_1/U_1/N345 ,
         \U_0/U_1/U_1/N344 , \U_0/U_1/U_1/N343 , \U_0/U_1/U_1/N342 ,
         \U_0/U_1/U_1/N341 , \U_0/U_1/U_1/N340 , \U_0/U_1/U_1/N339 ,
         \U_0/U_1/U_1/N338 , \U_0/U_1/U_1/N337 , \U_0/U_1/U_1/N336 ,
         \U_0/U_1/U_1/N335 , \U_0/U_1/U_1/N334 , \U_0/U_1/U_1/N333 ,
         \U_0/U_1/U_1/N195 , \U_0/U_1/U_1/N194 , \U_0/U_1/U_1/N193 ,
         \U_0/U_1/U_1/N192 , \U_0/U_1/U_1/N191 , \U_0/U_1/U_1/N190 ,
         \U_0/U_1/U_1/N189 , \U_0/U_1/U_1/N51 , \U_0/U_1/U_1/N50 ,
         \U_0/U_1/U_1/N49 , \U_0/U_1/U_1/N48 , \U_0/U_1/U_1/memory[0][7] ,
         \U_0/U_1/U_1/memory[0][6] , \U_0/U_1/U_1/memory[0][5] ,
         \U_0/U_1/U_1/memory[0][4] , \U_0/U_1/U_1/memory[0][3] ,
         \U_0/U_1/U_1/memory[0][2] , \U_0/U_1/U_1/memory[0][1] ,
         \U_0/U_1/U_1/memory[0][0] , \U_0/U_1/U_1/memory[1][7] ,
         \U_0/U_1/U_1/memory[1][6] , \U_0/U_1/U_1/memory[1][5] ,
         \U_0/U_1/U_1/memory[1][4] , \U_0/U_1/U_1/memory[1][3] ,
         \U_0/U_1/U_1/memory[1][2] , \U_0/U_1/U_1/memory[1][1] ,
         \U_0/U_1/U_1/memory[1][0] , \U_0/U_1/U_1/memory[2][7] ,
         \U_0/U_1/U_1/memory[2][6] , \U_0/U_1/U_1/memory[2][5] ,
         \U_0/U_1/U_1/memory[2][4] , \U_0/U_1/U_1/memory[2][3] ,
         \U_0/U_1/U_1/memory[2][2] , \U_0/U_1/U_1/memory[2][1] ,
         \U_0/U_1/U_1/memory[2][0] , \U_0/U_1/U_1/memory[3][7] ,
         \U_0/U_1/U_1/memory[3][6] , \U_0/U_1/U_1/memory[3][5] ,
         \U_0/U_1/U_1/memory[3][4] , \U_0/U_1/U_1/memory[3][3] ,
         \U_0/U_1/U_1/memory[3][2] , \U_0/U_1/U_1/memory[3][1] ,
         \U_0/U_1/U_1/memory[3][0] , \U_0/U_1/U_1/memory[4][7] ,
         \U_0/U_1/U_1/memory[4][6] , \U_0/U_1/U_1/memory[4][5] ,
         \U_0/U_1/U_1/memory[4][4] , \U_0/U_1/U_1/memory[4][3] ,
         \U_0/U_1/U_1/memory[4][2] , \U_0/U_1/U_1/memory[4][1] ,
         \U_0/U_1/U_1/memory[4][0] , \U_0/U_1/U_1/memory[5][7] ,
         \U_0/U_1/U_1/memory[5][6] , \U_0/U_1/U_1/memory[5][5] ,
         \U_0/U_1/U_1/memory[5][4] , \U_0/U_1/U_1/memory[5][3] ,
         \U_0/U_1/U_1/memory[5][2] , \U_0/U_1/U_1/memory[5][1] ,
         \U_0/U_1/U_1/memory[5][0] , \U_0/U_1/U_1/memory[6][7] ,
         \U_0/U_1/U_1/memory[6][6] , \U_0/U_1/U_1/memory[6][5] ,
         \U_0/U_1/U_1/memory[6][4] , \U_0/U_1/U_1/memory[6][3] ,
         \U_0/U_1/U_1/memory[6][2] , \U_0/U_1/U_1/memory[6][1] ,
         \U_0/U_1/U_1/memory[6][0] , \U_0/U_1/U_1/memory[7][7] ,
         \U_0/U_1/U_1/memory[7][6] , \U_0/U_1/U_1/memory[7][5] ,
         \U_0/U_1/U_1/memory[7][4] , \U_0/U_1/U_1/memory[7][3] ,
         \U_0/U_1/U_1/memory[7][2] , \U_0/U_1/U_1/memory[7][1] ,
         \U_0/U_1/U_1/memory[7][0] , \U_0/U_1/U_1/memory[8][7] ,
         \U_0/U_1/U_1/memory[8][6] , \U_0/U_1/U_1/memory[8][5] ,
         \U_0/U_1/U_1/memory[8][4] , \U_0/U_1/U_1/memory[8][3] ,
         \U_0/U_1/U_1/memory[8][2] , \U_0/U_1/U_1/memory[8][1] ,
         \U_0/U_1/U_1/memory[8][0] , \U_0/U_1/U_1/memory[9][7] ,
         \U_0/U_1/U_1/memory[9][6] , \U_0/U_1/U_1/memory[9][5] ,
         \U_0/U_1/U_1/memory[9][4] , \U_0/U_1/U_1/memory[9][3] ,
         \U_0/U_1/U_1/memory[9][2] , \U_0/U_1/U_1/memory[9][1] ,
         \U_0/U_1/U_1/memory[9][0] , \U_0/U_1/U_1/memory[10][7] ,
         \U_0/U_1/U_1/memory[10][6] , \U_0/U_1/U_1/memory[10][5] ,
         \U_0/U_1/U_1/memory[10][4] , \U_0/U_1/U_1/memory[10][3] ,
         \U_0/U_1/U_1/memory[10][2] , \U_0/U_1/U_1/memory[10][1] ,
         \U_0/U_1/U_1/memory[10][0] , \U_0/U_1/U_1/memory[11][7] ,
         \U_0/U_1/U_1/memory[11][6] , \U_0/U_1/U_1/memory[11][5] ,
         \U_0/U_1/U_1/memory[11][4] , \U_0/U_1/U_1/memory[11][3] ,
         \U_0/U_1/U_1/memory[11][2] , \U_0/U_1/U_1/memory[11][1] ,
         \U_0/U_1/U_1/memory[11][0] , \U_0/U_1/U_1/memory[12][7] ,
         \U_0/U_1/U_1/memory[12][6] , \U_0/U_1/U_1/memory[12][5] ,
         \U_0/U_1/U_1/memory[12][4] , \U_0/U_1/U_1/memory[12][3] ,
         \U_0/U_1/U_1/memory[12][2] , \U_0/U_1/U_1/memory[12][1] ,
         \U_0/U_1/U_1/memory[12][0] , \U_0/U_1/U_1/memory[13][7] ,
         \U_0/U_1/U_1/memory[13][6] , \U_0/U_1/U_1/memory[13][5] ,
         \U_0/U_1/U_1/memory[13][4] , \U_0/U_1/U_1/memory[13][3] ,
         \U_0/U_1/U_1/memory[13][2] , \U_0/U_1/U_1/memory[13][1] ,
         \U_0/U_1/U_1/memory[13][0] , \U_0/U_1/U_1/memory[14][7] ,
         \U_0/U_1/U_1/memory[14][6] , \U_0/U_1/U_1/memory[14][5] ,
         \U_0/U_1/U_1/memory[14][4] , \U_0/U_1/U_1/memory[14][3] ,
         \U_0/U_1/U_1/memory[14][2] , \U_0/U_1/U_1/memory[14][1] ,
         \U_0/U_1/U_1/memory[14][0] , \U_0/U_1/U_1/memory[15][7] ,
         \U_0/U_1/U_1/memory[15][6] , \U_0/U_1/U_1/memory[15][5] ,
         \U_0/U_1/U_1/memory[15][4] , \U_0/U_1/U_1/memory[15][3] ,
         \U_0/U_1/U_1/memory[15][2] , \U_0/U_1/U_1/memory[15][1] ,
         \U_0/U_1/U_1/memory[15][0] , \U_0/U_1/U_1/memory[16][7] ,
         \U_0/U_1/U_1/memory[16][6] , \U_0/U_1/U_1/memory[16][5] ,
         \U_0/U_1/U_1/memory[16][4] , \U_0/U_1/U_1/memory[16][3] ,
         \U_0/U_1/U_1/memory[16][2] , \U_0/U_1/U_1/memory[16][1] ,
         \U_0/U_1/U_1/memory[16][0] , \U_0/U_1/U_1/memory[17][7] ,
         \U_0/U_1/U_1/memory[17][6] , \U_0/U_1/U_1/memory[17][5] ,
         \U_0/U_1/U_1/memory[17][4] , \U_0/U_1/U_1/memory[17][3] ,
         \U_0/U_1/U_1/memory[17][2] , \U_0/U_1/U_1/memory[17][1] ,
         \U_0/U_1/U_1/memory[17][0] , \U_0/U_1/U_1/memory[18][7] ,
         \U_0/U_1/U_1/memory[18][6] , \U_0/U_1/U_1/memory[18][5] ,
         \U_0/U_1/U_1/memory[18][4] , \U_0/U_1/U_1/memory[18][3] ,
         \U_0/U_1/U_1/memory[18][2] , \U_0/U_1/U_1/memory[18][1] ,
         \U_0/U_1/U_1/memory[18][0] , \U_0/U_1/U_1/memory[19][7] ,
         \U_0/U_1/U_1/memory[19][6] , \U_0/U_1/U_1/memory[19][5] ,
         \U_0/U_1/U_1/memory[19][4] , \U_0/U_1/U_1/memory[19][3] ,
         \U_0/U_1/U_1/memory[19][2] , \U_0/U_1/U_1/memory[19][1] ,
         \U_0/U_1/U_1/memory[19][0] , \U_0/U_1/U_1/memory[20][7] ,
         \U_0/U_1/U_1/memory[20][6] , \U_0/U_1/U_1/memory[20][5] ,
         \U_0/U_1/U_1/memory[20][4] , \U_0/U_1/U_1/memory[20][3] ,
         \U_0/U_1/U_1/memory[20][2] , \U_0/U_1/U_1/memory[20][1] ,
         \U_0/U_1/U_1/memory[20][0] , \U_0/U_1/U_1/memory[21][7] ,
         \U_0/U_1/U_1/memory[21][6] , \U_0/U_1/U_1/memory[21][5] ,
         \U_0/U_1/U_1/memory[21][4] , \U_0/U_1/U_1/memory[21][3] ,
         \U_0/U_1/U_1/memory[21][2] , \U_0/U_1/U_1/memory[21][1] ,
         \U_0/U_1/U_1/memory[21][0] , \U_0/U_1/U_1/memory[22][7] ,
         \U_0/U_1/U_1/memory[22][6] , \U_0/U_1/U_1/memory[22][5] ,
         \U_0/U_1/U_1/memory[22][4] , \U_0/U_1/U_1/memory[22][3] ,
         \U_0/U_1/U_1/memory[22][2] , \U_0/U_1/U_1/memory[22][1] ,
         \U_0/U_1/U_1/memory[22][0] , \U_0/U_1/U_1/memory[23][7] ,
         \U_0/U_1/U_1/memory[23][6] , \U_0/U_1/U_1/memory[23][5] ,
         \U_0/U_1/U_1/memory[23][4] , \U_0/U_1/U_1/memory[23][3] ,
         \U_0/U_1/U_1/memory[23][2] , \U_0/U_1/U_1/memory[23][1] ,
         \U_0/U_1/U_1/memory[23][0] , \U_0/U_1/U_1/memory[24][7] ,
         \U_0/U_1/U_1/memory[24][6] , \U_0/U_1/U_1/memory[24][5] ,
         \U_0/U_1/U_1/memory[24][4] , \U_0/U_1/U_1/memory[24][3] ,
         \U_0/U_1/U_1/memory[24][2] , \U_0/U_1/U_1/memory[24][1] ,
         \U_0/U_1/U_1/memory[24][0] , \U_0/U_1/U_1/memory[25][7] ,
         \U_0/U_1/U_1/memory[25][6] , \U_0/U_1/U_1/memory[25][5] ,
         \U_0/U_1/U_1/memory[25][4] , \U_0/U_1/U_1/memory[25][3] ,
         \U_0/U_1/U_1/memory[25][2] , \U_0/U_1/U_1/memory[25][1] ,
         \U_0/U_1/U_1/memory[25][0] , \U_0/U_1/U_1/memory[26][7] ,
         \U_0/U_1/U_1/memory[26][6] , \U_0/U_1/U_1/memory[26][5] ,
         \U_0/U_1/U_1/memory[26][4] , \U_0/U_1/U_1/memory[26][3] ,
         \U_0/U_1/U_1/memory[26][2] , \U_0/U_1/U_1/memory[26][1] ,
         \U_0/U_1/U_1/memory[26][0] , \U_0/U_1/U_1/memory[27][7] ,
         \U_0/U_1/U_1/memory[27][6] , \U_0/U_1/U_1/memory[27][5] ,
         \U_0/U_1/U_1/memory[27][4] , \U_0/U_1/U_1/memory[27][3] ,
         \U_0/U_1/U_1/memory[27][2] , \U_0/U_1/U_1/memory[27][1] ,
         \U_0/U_1/U_1/memory[27][0] , \U_0/U_1/U_1/memory[28][7] ,
         \U_0/U_1/U_1/memory[28][6] , \U_0/U_1/U_1/memory[28][5] ,
         \U_0/U_1/U_1/memory[28][4] , \U_0/U_1/U_1/memory[28][3] ,
         \U_0/U_1/U_1/memory[28][2] , \U_0/U_1/U_1/memory[28][1] ,
         \U_0/U_1/U_1/memory[28][0] , \U_0/U_1/U_1/memory[29][7] ,
         \U_0/U_1/U_1/memory[29][6] , \U_0/U_1/U_1/memory[29][5] ,
         \U_0/U_1/U_1/memory[29][4] , \U_0/U_1/U_1/memory[29][3] ,
         \U_0/U_1/U_1/memory[29][2] , \U_0/U_1/U_1/memory[29][1] ,
         \U_0/U_1/U_1/memory[29][0] , \U_0/U_1/U_1/memory[30][7] ,
         \U_0/U_1/U_1/memory[30][6] , \U_0/U_1/U_1/memory[30][5] ,
         \U_0/U_1/U_1/memory[30][4] , \U_0/U_1/U_1/memory[30][3] ,
         \U_0/U_1/U_1/memory[30][2] , \U_0/U_1/U_1/memory[30][1] ,
         \U_0/U_1/U_1/memory[30][0] , \U_0/U_1/U_1/memory[31][7] ,
         \U_0/U_1/U_1/memory[31][6] , \U_0/U_1/U_1/memory[31][5] ,
         \U_0/U_1/U_1/memory[31][4] , \U_0/U_1/U_1/memory[31][3] ,
         \U_0/U_1/U_1/memory[31][2] , \U_0/U_1/U_1/memory[31][1] ,
         \U_0/U_1/U_1/memory[31][0] , \U_0/U_1/U_1/opcode[0][1] ,
         \U_0/U_1/U_1/opcode[0][0] , \U_0/U_1/U_1/opcode[1][1] ,
         \U_0/U_1/U_1/opcode[1][0] , \U_0/U_1/U_1/opcode[2][1] ,
         \U_0/U_1/U_1/opcode[2][0] , \U_0/U_1/U_1/opcode[3][1] ,
         \U_0/U_1/U_1/opcode[3][0] , \U_0/U_1/U_1/opcode[4][1] ,
         \U_0/U_1/U_1/opcode[4][0] , \U_0/U_1/U_1/opcode[5][1] ,
         \U_0/U_1/U_1/opcode[5][0] , \U_0/U_1/U_1/opcode[6][1] ,
         \U_0/U_1/U_1/opcode[6][0] , \U_0/U_1/U_1/opcode[7][1] ,
         \U_0/U_1/U_1/opcode[7][0] , \U_0/U_1/U_1/opcode[8][1] ,
         \U_0/U_1/U_1/opcode[8][0] , \U_0/U_1/U_1/opcode[9][1] ,
         \U_0/U_1/U_1/opcode[9][0] , \U_0/U_1/U_1/opcode[10][1] ,
         \U_0/U_1/U_1/opcode[10][0] , \U_0/U_1/U_1/opcode[11][1] ,
         \U_0/U_1/U_1/opcode[11][0] , \U_0/U_1/U_1/opcode[12][1] ,
         \U_0/U_1/U_1/opcode[12][0] , \U_0/U_1/U_1/opcode[13][1] ,
         \U_0/U_1/U_1/opcode[13][0] , \U_0/U_1/U_1/opcode[14][1] ,
         \U_0/U_1/U_1/opcode[14][0] , \U_0/U_1/U_1/opcode[15][1] ,
         \U_0/U_1/U_1/opcode[15][0] , \U_0/U_1/U_1/opcode[16][1] ,
         \U_0/U_1/U_1/opcode[16][0] , \U_0/U_1/U_1/opcode[17][1] ,
         \U_0/U_1/U_1/opcode[17][0] , \U_0/U_1/U_1/opcode[18][1] ,
         \U_0/U_1/U_1/opcode[18][0] , \U_0/U_1/U_1/opcode[19][1] ,
         \U_0/U_1/U_1/opcode[19][0] , \U_0/U_1/U_1/opcode[20][1] ,
         \U_0/U_1/U_1/opcode[20][0] , \U_0/U_1/U_1/opcode[21][1] ,
         \U_0/U_1/U_1/opcode[21][0] , \U_0/U_1/U_1/opcode[22][1] ,
         \U_0/U_1/U_1/opcode[22][0] , \U_0/U_1/U_1/opcode[23][1] ,
         \U_0/U_1/U_1/opcode[23][0] , \U_0/U_1/U_1/opcode[24][1] ,
         \U_0/U_1/U_1/opcode[24][0] , \U_0/U_1/U_1/opcode[25][1] ,
         \U_0/U_1/U_1/opcode[25][0] , \U_0/U_1/U_1/opcode[26][1] ,
         \U_0/U_1/U_1/opcode[26][0] , \U_0/U_1/U_1/opcode[27][1] ,
         \U_0/U_1/U_1/opcode[27][0] , \U_0/U_1/U_1/opcode[28][1] ,
         \U_0/U_1/U_1/opcode[28][0] , \U_0/U_1/U_1/opcode[29][1] ,
         \U_0/U_1/U_1/opcode[29][0] , \U_0/U_1/U_1/opcode[30][1] ,
         \U_0/U_1/U_1/opcode[30][0] , \U_0/U_1/U_1/opcode[31][1] ,
         \U_0/U_1/U_1/opcode[31][0] , \U_0/U_1/U_1/N46 , \U_0/U_1/U_1/N45 ,
         \U_0/U_1/U_1/N44 , \U_0/U_1/U_1/N43 , \U_0/U_1/U_1/N36 ,
         \U_0/U_1/U_1/N35 , \U_0/U_1/U_1/N34 , \U_0/U_1/U_1/N33 ,
         \U_0/U_1/U_1/N32 , \U_0/U_1/U_1/state , \U_0/U_1/U_1/writeptr[0] ,
         \U_0/U_1/U_1/writeptr[1] , \U_0/U_1/U_1/writeptr[2] ,
         \U_0/U_1/U_1/writeptr[3] , \U_0/U_1/U_1/writeptr[4] ,
         \U_0/U_1/U_1/readptr[0] , \U_0/U_1/U_1/readptr[1] ,
         \U_0/U_1/U_1/readptr[2] , \U_0/U_1/U_1/readptr[3] ,
         \U_0/U_1/U_1/readptr[4] , \U_0/U_2/U_2/current_crc[0] ,
         \U_0/U_2/U_2/current_crc[1] , \U_0/U_2/U_2/current_crc[2] ,
         \U_0/U_2/U_2/current_crc[3] , \U_0/U_2/U_2/current_crc[4] ,
         \U_0/U_2/U_2/current_crc[5] , \U_0/U_2/U_2/current_crc[6] ,
         \U_0/U_2/U_2/current_crc[7] , \U_0/U_2/U_2/current_crc[8] ,
         \U_0/U_2/U_2/current_crc[9] , \U_0/U_2/U_2/current_crc[10] ,
         \U_0/U_2/U_2/current_crc[11] , \U_0/U_2/U_2/current_crc[12] ,
         \U_0/U_2/U_2/current_crc[13] , \U_0/U_2/U_2/current_crc[14] ,
         \U_0/U_2/U_2/current_crc[15] , \U_0/U_2/U_1/N32 , \U_0/U_2/U_1/N31 ,
         \U_0/U_2/U_1/N29 , \U_0/U_2/U_1/state[0] , \U_0/U_2/U_1/state[1] ,
         \U_0/U_2/U_1/state[2] , \U_0/U_2/U_1/state[3] ,
         \U_0/U_2/U_1/DP_hold2 , \U_0/U_2/U_1/DP_hold1 ,
         \U_0/U_2/U_0/DP_hold2 , \U_0/U_2/U_0/DP_hold1 , \U_0/U_2/U_5/N170 ,
         \U_0/U_2/U_5/curCRC_ERROR , \U_0/U_2/U_5/curR_ERROR ,
         \U_0/U_2/U_5/count[0] , \U_0/U_2/U_5/count[1] ,
         \U_0/U_2/U_5/count[2] , \U_0/U_2/U_5/count[3] ,
         \U_0/U_2/U_5/state[0] , \U_0/U_2/U_5/state[1] ,
         \U_0/U_2/U_5/state[2] , \U_0/U_2/U_5/state[3] , \U_0/U_2/U_7/state ,
         \U_0/U_2/U_7/count[0] , \U_0/U_2/U_7/count[1] ,
         \U_0/U_2/U_7/count[2] , \U_0/U_2/U_7/count[3] , \U_0/U_3/d_encode ,
         \U_0/U_3/SHIFT_ENABLE_E , \U_0/U_3/U_0/N59 , \U_0/U_3/U_0/dm_tx_nxt ,
         \U_0/U_3/U_0/DE_holdout_nxt , \U_0/U_3/U_0/DE_holdout_last ,
         \U_0/U_3/U_0/state[0] , \U_0/U_3/U_0/state[1] ,
         \U_0/U_3/U_0/state[2] , \U_0/U_3/U_0/state[3] ,
         \U_0/U_3/U_0/DE_holdout_BS , \U_0/U_3/U_0/DE_holdout ,
         \U_0/U_3/U_2/count[0] , \U_0/U_3/U_2/count[1] ,
         \U_0/U_3/U_2/count[2] , \U_0/U_3/U_3/N188 , \U_0/U_3/U_3/N187 ,
         \U_0/U_3/U_3/N90 , \U_0/U_3/U_3/N89 , \U_0/U_3/U_3/N88 ,
         \U_0/U_3/U_3/N87 , \U_0/U_3/U_3/N86 , \U_0/U_3/U_3/N85 ,
         \U_0/U_3/U_3/N84 , \U_0/U_3/U_3/N65 , \U_0/U_3/U_3/N64 ,
         \U_0/U_3/U_3/N63 , \U_0/U_3/U_3/N62 , \U_0/U_3/U_3/N61 ,
         \U_0/U_3/U_3/N60 , \U_0/U_3/U_3/N59 , \U_0/U_3/U_3/count[0] ,
         \U_0/U_3/U_3/count[1] , \U_0/U_3/U_3/count[2] ,
         \U_0/U_3/U_3/count[3] , \U_0/U_3/U_3/count[4] ,
         \U_0/U_3/U_3/count[5] , \U_0/U_3/U_3/state[0] ,
         \U_0/U_3/U_3/state[1] , \U_0/U_3/U_3/state[2] , \U_0/U_3/U_4/state ,
         \U_0/U_3/U_4/count[0] , \U_0/U_3/U_4/count[1] ,
         \U_0/U_3/U_4/count[2] , \U_0/U_3/U_4/count[3] , \U_1/PDATA_READY ,
         \U_1/PRGA_OPCODE[0] , \U_1/PRGA_OPCODE[1] , \U_1/B_READY ,
         \U_1/RBUF_FULL , \U_1/U_0/U_0/N527 , \U_1/U_0/U_0/N526 ,
         \U_1/U_0/U_0/N525 , \U_1/U_0/U_0/N524 , \U_1/U_0/U_0/N523 ,
         \U_1/U_0/U_0/N522 , \U_1/U_0/U_0/N521 , \U_1/U_0/U_0/N520 ,
         \U_1/U_0/U_0/N519 , \U_1/U_0/U_0/N518 , \U_1/U_0/U_0/N517 ,
         \U_1/U_0/U_0/N516 , \U_1/U_0/U_0/N515 , \U_1/U_0/U_0/N514 ,
         \U_1/U_0/U_0/N513 , \U_1/U_0/U_0/N512 , \U_1/U_0/U_0/N503 ,
         \U_1/U_0/U_0/N502 , \U_1/U_0/U_0/N501 , \U_1/U_0/U_0/N500 ,
         \U_1/U_0/U_0/N499 , \U_1/U_0/U_0/N498 , \U_1/U_0/U_0/N497 ,
         \U_1/U_0/U_0/N496 , \U_1/U_0/U_0/N487 , \U_1/U_0/U_0/N486 ,
         \U_1/U_0/U_0/N485 , \U_1/U_0/U_0/N484 , \U_1/U_0/U_0/N483 ,
         \U_1/U_0/U_0/N482 , \U_1/U_0/U_0/N481 , \U_1/U_0/U_0/N480 ,
         \U_1/U_0/U_0/N479 , \U_1/U_0/U_0/N478 , \U_1/U_0/U_0/N477 ,
         \U_1/U_0/U_0/N476 , \U_1/U_0/U_0/N475 , \U_1/U_0/U_0/N474 ,
         \U_1/U_0/U_0/N473 , \U_1/U_0/U_0/N472 , \U_1/U_0/U_0/N448 ,
         \U_1/U_0/U_0/N447 , \U_1/U_0/U_0/N446 , \U_1/U_0/U_0/N445 ,
         \U_1/U_0/U_0/N444 , \U_1/U_0/U_0/N443 , \U_1/U_0/U_0/N442 ,
         \U_1/U_0/U_0/N431 , \U_1/U_0/U_0/N430 , \U_1/U_0/U_0/N429 ,
         \U_1/U_0/U_0/N428 , \U_1/U_0/U_0/N427 , \U_1/U_0/U_0/N426 ,
         \U_1/U_0/U_0/N425 , \U_1/U_0/U_0/N424 , \U_1/U_0/U_0/N414 ,
         \U_1/U_0/U_0/N413 , \U_1/U_0/U_0/N412 , \U_1/U_0/U_0/N411 ,
         \U_1/U_0/U_0/N410 , \U_1/U_0/U_0/N409 , \U_1/U_0/U_0/N408 ,
         \U_1/U_0/U_0/N407 , \U_1/U_0/U_0/fr_enable , \U_1/U_0/U_0/fw_enable ,
         \U_1/U_0/U_0/prefillCounter[0] , \U_1/U_0/U_0/prefillCounter[1] ,
         \U_1/U_0/U_0/prefillCounter[2] , \U_1/U_0/U_0/prefillCounter[3] ,
         \U_1/U_0/U_0/prefillCounter[4] , \U_1/U_0/U_0/prefillCounter[5] ,
         \U_1/U_0/U_0/prefillCounter[6] , \U_1/U_0/U_0/prefillCounter[7] ,
         \U_1/U_0/U_0/keyTable[0][7] , \U_1/U_0/U_0/keyTable[0][6] ,
         \U_1/U_0/U_0/keyTable[0][5] , \U_1/U_0/U_0/keyTable[0][4] ,
         \U_1/U_0/U_0/keyTable[0][3] , \U_1/U_0/U_0/keyTable[0][2] ,
         \U_1/U_0/U_0/keyTable[0][1] , \U_1/U_0/U_0/keyTable[0][0] ,
         \U_1/U_0/U_0/keyTable[1][7] , \U_1/U_0/U_0/keyTable[1][6] ,
         \U_1/U_0/U_0/keyTable[1][5] , \U_1/U_0/U_0/keyTable[1][4] ,
         \U_1/U_0/U_0/keyTable[1][3] , \U_1/U_0/U_0/keyTable[1][2] ,
         \U_1/U_0/U_0/keyTable[1][1] , \U_1/U_0/U_0/keyTable[1][0] ,
         \U_1/U_0/U_0/keyTable[2][7] , \U_1/U_0/U_0/keyTable[2][6] ,
         \U_1/U_0/U_0/keyTable[2][5] , \U_1/U_0/U_0/keyTable[2][4] ,
         \U_1/U_0/U_0/keyTable[2][3] , \U_1/U_0/U_0/keyTable[2][2] ,
         \U_1/U_0/U_0/keyTable[2][1] , \U_1/U_0/U_0/keyTable[2][0] ,
         \U_1/U_0/U_0/keyTable[3][7] , \U_1/U_0/U_0/keyTable[3][6] ,
         \U_1/U_0/U_0/keyTable[3][5] , \U_1/U_0/U_0/keyTable[3][4] ,
         \U_1/U_0/U_0/keyTable[3][3] , \U_1/U_0/U_0/keyTable[3][2] ,
         \U_1/U_0/U_0/keyTable[3][1] , \U_1/U_0/U_0/keyTable[3][0] ,
         \U_1/U_0/U_0/keyTable[4][7] , \U_1/U_0/U_0/keyTable[4][6] ,
         \U_1/U_0/U_0/keyTable[4][5] , \U_1/U_0/U_0/keyTable[4][4] ,
         \U_1/U_0/U_0/keyTable[4][3] , \U_1/U_0/U_0/keyTable[4][2] ,
         \U_1/U_0/U_0/keyTable[4][1] , \U_1/U_0/U_0/keyTable[4][0] ,
         \U_1/U_0/U_0/keyTable[5][7] , \U_1/U_0/U_0/keyTable[5][6] ,
         \U_1/U_0/U_0/keyTable[5][5] , \U_1/U_0/U_0/keyTable[5][4] ,
         \U_1/U_0/U_0/keyTable[5][3] , \U_1/U_0/U_0/keyTable[5][2] ,
         \U_1/U_0/U_0/keyTable[5][1] , \U_1/U_0/U_0/keyTable[5][0] ,
         \U_1/U_0/U_0/keyTable[6][7] , \U_1/U_0/U_0/keyTable[6][6] ,
         \U_1/U_0/U_0/keyTable[6][5] , \U_1/U_0/U_0/keyTable[6][4] ,
         \U_1/U_0/U_0/keyTable[6][3] , \U_1/U_0/U_0/keyTable[6][2] ,
         \U_1/U_0/U_0/keyTable[6][1] , \U_1/U_0/U_0/keyTable[6][0] ,
         \U_1/U_0/U_0/keyTable[7][7] , \U_1/U_0/U_0/keyTable[7][6] ,
         \U_1/U_0/U_0/keyTable[7][5] , \U_1/U_0/U_0/keyTable[7][4] ,
         \U_1/U_0/U_0/keyTable[7][3] , \U_1/U_0/U_0/keyTable[7][2] ,
         \U_1/U_0/U_0/keyTable[7][1] , \U_1/U_0/U_0/keyTable[7][0] ,
         \U_1/U_0/U_0/nextProcessedData[0] ,
         \U_1/U_0/U_0/nextProcessedData[1] ,
         \U_1/U_0/U_0/nextProcessedData[2] ,
         \U_1/U_0/U_0/nextProcessedData[3] ,
         \U_1/U_0/U_0/nextProcessedData[4] ,
         \U_1/U_0/U_0/nextProcessedData[5] ,
         \U_1/U_0/U_0/nextProcessedData[6] ,
         \U_1/U_0/U_0/nextProcessedData[7] , \U_1/U_0/U_0/extratemp[0] ,
         \U_1/U_0/U_0/extratemp[1] , \U_1/U_0/U_0/extratemp[2] ,
         \U_1/U_0/U_0/extratemp[3] , \U_1/U_0/U_0/extratemp[4] ,
         \U_1/U_0/U_0/extratemp[5] , \U_1/U_0/U_0/extratemp[6] ,
         \U_1/U_0/U_0/extratemp[7] , \U_1/U_0/U_0/temp[0] ,
         \U_1/U_0/U_0/temp[1] , \U_1/U_0/U_0/temp[2] , \U_1/U_0/U_0/temp[3] ,
         \U_1/U_0/U_0/temp[4] , \U_1/U_0/U_0/temp[5] , \U_1/U_0/U_0/temp[6] ,
         \U_1/U_0/U_0/temp[7] , \U_1/U_0/U_0/permuteComplete ,
         \U_1/U_0/U_0/keyi[0] , \U_1/U_0/U_0/keyi[1] , \U_1/U_0/U_0/keyi[2] ,
         \U_1/U_0/U_0/intj[0] , \U_1/U_0/U_0/intj[1] , \U_1/U_0/U_0/intj[2] ,
         \U_1/U_0/U_0/intj[3] , \U_1/U_0/U_0/intj[4] , \U_1/U_0/U_0/intj[5] ,
         \U_1/U_0/U_0/intj[6] , \U_1/U_0/U_0/intj[7] , \U_1/U_0/U_0/inti[0] ,
         \U_1/U_0/U_0/inti[1] , \U_1/U_0/U_0/inti[2] , \U_1/U_0/U_0/inti[3] ,
         \U_1/U_0/U_0/inti[4] , \U_1/U_0/U_0/inti[5] , \U_1/U_0/U_0/inti[6] ,
         \U_1/U_0/U_0/inti[7] , \U_1/U_0/U_0/sj[0] , \U_1/U_0/U_0/sj[1] ,
         \U_1/U_0/U_0/sj[2] , \U_1/U_0/U_0/sj[3] , \U_1/U_0/U_0/sj[4] ,
         \U_1/U_0/U_0/sj[5] , \U_1/U_0/U_0/sj[6] , \U_1/U_0/U_0/sj[7] ,
         \U_1/U_0/U_0/si[0] , \U_1/U_0/U_0/si[1] , \U_1/U_0/U_0/si[2] ,
         \U_1/U_0/U_0/si[3] , \U_1/U_0/U_0/si[4] , \U_1/U_0/U_0/si[5] ,
         \U_1/U_0/U_0/si[6] , \U_1/U_0/U_0/si[7] , \U_1/U_0/U_0/state[0] ,
         \U_1/U_0/U_0/state[1] , \U_1/U_0/U_0/state[2] ,
         \U_1/U_0/U_0/state[3] , \U_1/U_0/U_0/state[4] , \U_1/U_0/U_1/SBE ,
         \U_1/U_0/U_1/TIMER_TRIG , \U_1/U_0/U_1/SET_RBUF_FULL ,
         \U_1/U_0/U_1/SBC_EN , \U_1/U_0/U_1/SBC_CLR , \U_1/U_0/U_1/RBUF_LOAD ,
         \U_1/U_0/U_1/SB_DETECT , \U_1/U_0/U_1/OE , \U_1/U_0/U_1/CHK_ERROR ,
         \U_1/U_0/U_1/U_0/Q_int2 , \U_1/U_0/U_1/U_0/Q_int ,
         \U_1/U_0/U_1/U_1/OE_prime , \U_1/U_0/U_1/U_2/N99 ,
         \U_1/U_0/U_1/U_2/N38 , \U_1/U_0/U_1/U_2/N37 , \U_1/U_0/U_1/U_2/N36 ,
         \U_1/U_0/U_1/U_2/N35 , \U_1/U_0/U_1/U_2/N34 , \U_1/U_0/U_1/U_2/N33 ,
         \U_1/U_0/U_1/U_2/N32 , \U_1/U_0/U_1/U_2/N31 , \U_1/U_0/U_1/U_2/N30 ,
         \U_1/U_0/U_1/U_2/N29 , \U_1/U_0/U_1/U_2/N28 , \U_1/U_0/U_1/U_2/N27 ,
         \U_1/U_0/U_1/U_2/N26 , \U_1/U_0/U_1/U_2/N25 , \U_1/U_0/U_1/U_2/N24 ,
         \U_1/U_0/U_1/U_2/N23 , \U_1/U_0/U_1/U_2/nextState[0] ,
         \U_1/U_0/U_1/U_2/nextState[1] , \U_1/U_0/U_1/U_2/nextState[2] ,
         \U_1/U_0/U_1/U_2/count[1] , \U_1/U_0/U_1/U_2/count[2] ,
         \U_1/U_0/U_1/U_2/count[3] , \U_1/U_0/U_1/U_2/count[4] ,
         \U_1/U_0/U_1/U_2/count[5] , \U_1/U_0/U_1/U_2/count[6] ,
         \U_1/U_0/U_1/U_2/count[7] , \U_1/U_0/U_1/U_2/timerRunning ,
         \U_1/U_0/U_1/U_2/state[0] , \U_1/U_0/U_1/U_2/state[1] ,
         \U_1/U_0/U_1/U_2/state[2] , \U_1/U_0/U_1/U_5/sb_detect_flag ,
         \U_1/U_0/U_1/U_5/SBE_prime , \U_1/U_0/U_1/U_8/N1799 ,
         \U_1/U_0/U_1/U_8/N1798 , \U_1/U_0/U_1/U_8/N1797 ,
         \U_1/U_0/U_1/U_8/N1796 , \U_1/U_0/U_1/U_8/N1795 ,
         \U_1/U_0/U_1/U_8/N1794 , \U_1/U_0/U_1/U_8/N1793 ,
         \U_1/U_0/U_1/U_8/N1792 , \U_1/U_0/U_1/U_8/nextParityError ,
         \U_1/U_0/U_1/U_8/parityAccumulator[0] ,
         \U_1/U_0/U_1/U_8/parityAccumulator[1] ,
         \U_1/U_0/U_1/U_8/parityAccumulator[2] ,
         \U_1/U_0/U_1/U_8/parityAccumulator[3] ,
         \U_1/U_0/U_1/U_8/parityAccumulator[4] ,
         \U_1/U_0/U_1/U_8/parityAccumulator[5] ,
         \U_1/U_0/U_1/U_8/parityAccumulator[6] ,
         \U_1/U_0/U_1/U_8/parityAccumulator[7] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[0] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[1] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[2] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[3] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[4] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[5] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[6] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[7] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[8] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[9] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[10] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[11] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[12] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[13] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[14] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[15] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[16] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[17] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[18] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[19] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[20] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[21] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[22] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[23] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[24] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[25] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[26] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[27] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[28] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[29] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[30] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[31] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[32] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[33] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[34] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[35] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[36] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[37] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[38] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[39] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[40] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[41] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[42] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[43] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[44] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[45] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[46] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[47] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[48] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[49] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[50] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[51] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[52] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[53] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[54] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[55] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[56] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[57] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[58] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[59] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[60] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[61] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[62] ,
         \U_1/U_0/U_1/U_8/currentPlainKey[63] , \U_1/U_0/U_1/U_8/address[0] ,
         \U_1/U_0/U_1/U_8/address[1] , \U_1/U_0/U_1/U_8/address[2] ,
         \U_1/U_0/U_1/U_8/address[3] , \U_1/U_0/U_1/U_8/address[4] ,
         \U_1/U_0/U_1/U_8/address[5] , \U_1/U_0/U_1/U_8/address[6] ,
         \U_1/U_0/U_1/U_8/address[7] , \U_1/U_0/U_1/U_8/keyCount[0] ,
         \U_1/U_0/U_1/U_8/keyCount[1] , \U_1/U_0/U_1/U_8/keyCount[2] ,
         \U_1/U_0/U_1/U_8/keyCount[3] , \U_1/U_0/U_1/U_8/parityError ,
         \U_1/U_0/U_1/U_8/state[0] , \U_1/U_0/U_1/U_8/state[1] ,
         \U_1/U_0/U_1/U_8/state[2] , \U_1/U_0/U_1/U_8/state[3] ,
         \U_1/U_0/U_1/U_7/N33 , \U_1/U_0/U_1/U_7/N32 , \U_1/U_0/U_1/U_7/N31 ,
         \U_1/U_0/U_1/U_7/N30 , \U_1/U_0/U_1/U_7/N29 , \U_1/U_0/U_1/U_7/N28 ,
         \U_1/U_0/U_1/U_7/N27 , \U_1/U_0/U_1/U_7/N26 ,
         \U_1/U_0/U_1/U_7/nextState[0] , \U_1/U_0/U_1/U_7/nextState[1] ,
         \U_1/U_0/U_1/U_7/nextState[2] , \U_1/U_0/U_1/U_7/nextState[3] ,
         \U_1/U_0/U_1/U_7/nextState[4] , \U_1/U_0/U_1/U_7/nextState[5] ,
         \U_1/U_0/U_1/U_7/nextState[6] , \U_1/U_0/U_1/U_7/nextState[7] ,
         \U_1/U_0/U_1/U_7/state[0] , \U_1/U_0/U_1/U_7/state[1] ,
         \U_1/U_0/U_1/U_7/state[2] , \U_1/U_0/U_1/U_7/state[3] ,
         \U_1/U_0/U_1/U_7/state[4] , \U_1/U_0/U_1/U_7/state[5] ,
         \U_1/U_0/U_1/U_7/state[6] , \U_1/U_0/U_1/U_7/state[7] ,
         \U_1/U_1/R_ENABLE , \U_1/U_1/U_0/N40 , \U_1/U_1/U_0/N39 ,
         \U_1/U_1/U_0/state[0] , \U_1/U_1/U_0/state[1] ,
         \U_1/U_1/U_0/state[2] , \U_1/U_1/U_1/N355 , \U_1/U_1/U_1/N349 ,
         \U_1/U_1/U_1/N347 , \U_1/U_1/U_1/N346 , \U_1/U_1/U_1/N345 ,
         \U_1/U_1/U_1/N344 , \U_1/U_1/U_1/N343 , \U_1/U_1/U_1/N342 ,
         \U_1/U_1/U_1/N341 , \U_1/U_1/U_1/N340 , \U_1/U_1/U_1/N339 ,
         \U_1/U_1/U_1/N338 , \U_1/U_1/U_1/N337 , \U_1/U_1/U_1/N336 ,
         \U_1/U_1/U_1/N335 , \U_1/U_1/U_1/N334 , \U_1/U_1/U_1/N333 ,
         \U_1/U_1/U_1/N195 , \U_1/U_1/U_1/N194 , \U_1/U_1/U_1/N193 ,
         \U_1/U_1/U_1/N192 , \U_1/U_1/U_1/N191 , \U_1/U_1/U_1/N190 ,
         \U_1/U_1/U_1/N189 , \U_1/U_1/U_1/N51 , \U_1/U_1/U_1/N50 ,
         \U_1/U_1/U_1/N49 , \U_1/U_1/U_1/N48 , \U_1/U_1/U_1/memory[0][7] ,
         \U_1/U_1/U_1/memory[0][6] , \U_1/U_1/U_1/memory[0][5] ,
         \U_1/U_1/U_1/memory[0][4] , \U_1/U_1/U_1/memory[0][3] ,
         \U_1/U_1/U_1/memory[0][2] , \U_1/U_1/U_1/memory[0][1] ,
         \U_1/U_1/U_1/memory[0][0] , \U_1/U_1/U_1/memory[1][7] ,
         \U_1/U_1/U_1/memory[1][6] , \U_1/U_1/U_1/memory[1][5] ,
         \U_1/U_1/U_1/memory[1][4] , \U_1/U_1/U_1/memory[1][3] ,
         \U_1/U_1/U_1/memory[1][2] , \U_1/U_1/U_1/memory[1][1] ,
         \U_1/U_1/U_1/memory[1][0] , \U_1/U_1/U_1/memory[2][7] ,
         \U_1/U_1/U_1/memory[2][6] , \U_1/U_1/U_1/memory[2][5] ,
         \U_1/U_1/U_1/memory[2][4] , \U_1/U_1/U_1/memory[2][3] ,
         \U_1/U_1/U_1/memory[2][2] , \U_1/U_1/U_1/memory[2][1] ,
         \U_1/U_1/U_1/memory[2][0] , \U_1/U_1/U_1/memory[3][7] ,
         \U_1/U_1/U_1/memory[3][6] , \U_1/U_1/U_1/memory[3][5] ,
         \U_1/U_1/U_1/memory[3][4] , \U_1/U_1/U_1/memory[3][3] ,
         \U_1/U_1/U_1/memory[3][2] , \U_1/U_1/U_1/memory[3][1] ,
         \U_1/U_1/U_1/memory[3][0] , \U_1/U_1/U_1/memory[4][7] ,
         \U_1/U_1/U_1/memory[4][6] , \U_1/U_1/U_1/memory[4][5] ,
         \U_1/U_1/U_1/memory[4][4] , \U_1/U_1/U_1/memory[4][3] ,
         \U_1/U_1/U_1/memory[4][2] , \U_1/U_1/U_1/memory[4][1] ,
         \U_1/U_1/U_1/memory[4][0] , \U_1/U_1/U_1/memory[5][7] ,
         \U_1/U_1/U_1/memory[5][6] , \U_1/U_1/U_1/memory[5][5] ,
         \U_1/U_1/U_1/memory[5][4] , \U_1/U_1/U_1/memory[5][3] ,
         \U_1/U_1/U_1/memory[5][2] , \U_1/U_1/U_1/memory[5][1] ,
         \U_1/U_1/U_1/memory[5][0] , \U_1/U_1/U_1/memory[6][7] ,
         \U_1/U_1/U_1/memory[6][6] , \U_1/U_1/U_1/memory[6][5] ,
         \U_1/U_1/U_1/memory[6][4] , \U_1/U_1/U_1/memory[6][3] ,
         \U_1/U_1/U_1/memory[6][2] , \U_1/U_1/U_1/memory[6][1] ,
         \U_1/U_1/U_1/memory[6][0] , \U_1/U_1/U_1/memory[7][7] ,
         \U_1/U_1/U_1/memory[7][6] , \U_1/U_1/U_1/memory[7][5] ,
         \U_1/U_1/U_1/memory[7][4] , \U_1/U_1/U_1/memory[7][3] ,
         \U_1/U_1/U_1/memory[7][2] , \U_1/U_1/U_1/memory[7][1] ,
         \U_1/U_1/U_1/memory[7][0] , \U_1/U_1/U_1/memory[8][7] ,
         \U_1/U_1/U_1/memory[8][6] , \U_1/U_1/U_1/memory[8][5] ,
         \U_1/U_1/U_1/memory[8][4] , \U_1/U_1/U_1/memory[8][3] ,
         \U_1/U_1/U_1/memory[8][2] , \U_1/U_1/U_1/memory[8][1] ,
         \U_1/U_1/U_1/memory[8][0] , \U_1/U_1/U_1/memory[9][7] ,
         \U_1/U_1/U_1/memory[9][6] , \U_1/U_1/U_1/memory[9][5] ,
         \U_1/U_1/U_1/memory[9][4] , \U_1/U_1/U_1/memory[9][3] ,
         \U_1/U_1/U_1/memory[9][2] , \U_1/U_1/U_1/memory[9][1] ,
         \U_1/U_1/U_1/memory[9][0] , \U_1/U_1/U_1/memory[10][7] ,
         \U_1/U_1/U_1/memory[10][6] , \U_1/U_1/U_1/memory[10][5] ,
         \U_1/U_1/U_1/memory[10][4] , \U_1/U_1/U_1/memory[10][3] ,
         \U_1/U_1/U_1/memory[10][2] , \U_1/U_1/U_1/memory[10][1] ,
         \U_1/U_1/U_1/memory[10][0] , \U_1/U_1/U_1/memory[11][7] ,
         \U_1/U_1/U_1/memory[11][6] , \U_1/U_1/U_1/memory[11][5] ,
         \U_1/U_1/U_1/memory[11][4] , \U_1/U_1/U_1/memory[11][3] ,
         \U_1/U_1/U_1/memory[11][2] , \U_1/U_1/U_1/memory[11][1] ,
         \U_1/U_1/U_1/memory[11][0] , \U_1/U_1/U_1/memory[12][7] ,
         \U_1/U_1/U_1/memory[12][6] , \U_1/U_1/U_1/memory[12][5] ,
         \U_1/U_1/U_1/memory[12][4] , \U_1/U_1/U_1/memory[12][3] ,
         \U_1/U_1/U_1/memory[12][2] , \U_1/U_1/U_1/memory[12][1] ,
         \U_1/U_1/U_1/memory[12][0] , \U_1/U_1/U_1/memory[13][7] ,
         \U_1/U_1/U_1/memory[13][6] , \U_1/U_1/U_1/memory[13][5] ,
         \U_1/U_1/U_1/memory[13][4] , \U_1/U_1/U_1/memory[13][3] ,
         \U_1/U_1/U_1/memory[13][2] , \U_1/U_1/U_1/memory[13][1] ,
         \U_1/U_1/U_1/memory[13][0] , \U_1/U_1/U_1/memory[14][7] ,
         \U_1/U_1/U_1/memory[14][6] , \U_1/U_1/U_1/memory[14][5] ,
         \U_1/U_1/U_1/memory[14][4] , \U_1/U_1/U_1/memory[14][3] ,
         \U_1/U_1/U_1/memory[14][2] , \U_1/U_1/U_1/memory[14][1] ,
         \U_1/U_1/U_1/memory[14][0] , \U_1/U_1/U_1/memory[15][7] ,
         \U_1/U_1/U_1/memory[15][6] , \U_1/U_1/U_1/memory[15][5] ,
         \U_1/U_1/U_1/memory[15][4] , \U_1/U_1/U_1/memory[15][3] ,
         \U_1/U_1/U_1/memory[15][2] , \U_1/U_1/U_1/memory[15][1] ,
         \U_1/U_1/U_1/memory[15][0] , \U_1/U_1/U_1/memory[16][7] ,
         \U_1/U_1/U_1/memory[16][6] , \U_1/U_1/U_1/memory[16][5] ,
         \U_1/U_1/U_1/memory[16][4] , \U_1/U_1/U_1/memory[16][3] ,
         \U_1/U_1/U_1/memory[16][2] , \U_1/U_1/U_1/memory[16][1] ,
         \U_1/U_1/U_1/memory[16][0] , \U_1/U_1/U_1/memory[17][7] ,
         \U_1/U_1/U_1/memory[17][6] , \U_1/U_1/U_1/memory[17][5] ,
         \U_1/U_1/U_1/memory[17][4] , \U_1/U_1/U_1/memory[17][3] ,
         \U_1/U_1/U_1/memory[17][2] , \U_1/U_1/U_1/memory[17][1] ,
         \U_1/U_1/U_1/memory[17][0] , \U_1/U_1/U_1/memory[18][7] ,
         \U_1/U_1/U_1/memory[18][6] , \U_1/U_1/U_1/memory[18][5] ,
         \U_1/U_1/U_1/memory[18][4] , \U_1/U_1/U_1/memory[18][3] ,
         \U_1/U_1/U_1/memory[18][2] , \U_1/U_1/U_1/memory[18][1] ,
         \U_1/U_1/U_1/memory[18][0] , \U_1/U_1/U_1/memory[19][7] ,
         \U_1/U_1/U_1/memory[19][6] , \U_1/U_1/U_1/memory[19][5] ,
         \U_1/U_1/U_1/memory[19][4] , \U_1/U_1/U_1/memory[19][3] ,
         \U_1/U_1/U_1/memory[19][2] , \U_1/U_1/U_1/memory[19][1] ,
         \U_1/U_1/U_1/memory[19][0] , \U_1/U_1/U_1/memory[20][7] ,
         \U_1/U_1/U_1/memory[20][6] , \U_1/U_1/U_1/memory[20][5] ,
         \U_1/U_1/U_1/memory[20][4] , \U_1/U_1/U_1/memory[20][3] ,
         \U_1/U_1/U_1/memory[20][2] , \U_1/U_1/U_1/memory[20][1] ,
         \U_1/U_1/U_1/memory[20][0] , \U_1/U_1/U_1/memory[21][7] ,
         \U_1/U_1/U_1/memory[21][6] , \U_1/U_1/U_1/memory[21][5] ,
         \U_1/U_1/U_1/memory[21][4] , \U_1/U_1/U_1/memory[21][3] ,
         \U_1/U_1/U_1/memory[21][2] , \U_1/U_1/U_1/memory[21][1] ,
         \U_1/U_1/U_1/memory[21][0] , \U_1/U_1/U_1/memory[22][7] ,
         \U_1/U_1/U_1/memory[22][6] , \U_1/U_1/U_1/memory[22][5] ,
         \U_1/U_1/U_1/memory[22][4] , \U_1/U_1/U_1/memory[22][3] ,
         \U_1/U_1/U_1/memory[22][2] , \U_1/U_1/U_1/memory[22][1] ,
         \U_1/U_1/U_1/memory[22][0] , \U_1/U_1/U_1/memory[23][7] ,
         \U_1/U_1/U_1/memory[23][6] , \U_1/U_1/U_1/memory[23][5] ,
         \U_1/U_1/U_1/memory[23][4] , \U_1/U_1/U_1/memory[23][3] ,
         \U_1/U_1/U_1/memory[23][2] , \U_1/U_1/U_1/memory[23][1] ,
         \U_1/U_1/U_1/memory[23][0] , \U_1/U_1/U_1/memory[24][7] ,
         \U_1/U_1/U_1/memory[24][6] , \U_1/U_1/U_1/memory[24][5] ,
         \U_1/U_1/U_1/memory[24][4] , \U_1/U_1/U_1/memory[24][3] ,
         \U_1/U_1/U_1/memory[24][2] , \U_1/U_1/U_1/memory[24][1] ,
         \U_1/U_1/U_1/memory[24][0] , \U_1/U_1/U_1/memory[25][7] ,
         \U_1/U_1/U_1/memory[25][6] , \U_1/U_1/U_1/memory[25][5] ,
         \U_1/U_1/U_1/memory[25][4] , \U_1/U_1/U_1/memory[25][3] ,
         \U_1/U_1/U_1/memory[25][2] , \U_1/U_1/U_1/memory[25][1] ,
         \U_1/U_1/U_1/memory[25][0] , \U_1/U_1/U_1/memory[26][7] ,
         \U_1/U_1/U_1/memory[26][6] , \U_1/U_1/U_1/memory[26][5] ,
         \U_1/U_1/U_1/memory[26][4] , \U_1/U_1/U_1/memory[26][3] ,
         \U_1/U_1/U_1/memory[26][2] , \U_1/U_1/U_1/memory[26][1] ,
         \U_1/U_1/U_1/memory[26][0] , \U_1/U_1/U_1/memory[27][7] ,
         \U_1/U_1/U_1/memory[27][6] , \U_1/U_1/U_1/memory[27][5] ,
         \U_1/U_1/U_1/memory[27][4] , \U_1/U_1/U_1/memory[27][3] ,
         \U_1/U_1/U_1/memory[27][2] , \U_1/U_1/U_1/memory[27][1] ,
         \U_1/U_1/U_1/memory[27][0] , \U_1/U_1/U_1/memory[28][7] ,
         \U_1/U_1/U_1/memory[28][6] , \U_1/U_1/U_1/memory[28][5] ,
         \U_1/U_1/U_1/memory[28][4] , \U_1/U_1/U_1/memory[28][3] ,
         \U_1/U_1/U_1/memory[28][2] , \U_1/U_1/U_1/memory[28][1] ,
         \U_1/U_1/U_1/memory[28][0] , \U_1/U_1/U_1/memory[29][7] ,
         \U_1/U_1/U_1/memory[29][6] , \U_1/U_1/U_1/memory[29][5] ,
         \U_1/U_1/U_1/memory[29][4] , \U_1/U_1/U_1/memory[29][3] ,
         \U_1/U_1/U_1/memory[29][2] , \U_1/U_1/U_1/memory[29][1] ,
         \U_1/U_1/U_1/memory[29][0] , \U_1/U_1/U_1/memory[30][7] ,
         \U_1/U_1/U_1/memory[30][6] , \U_1/U_1/U_1/memory[30][5] ,
         \U_1/U_1/U_1/memory[30][4] , \U_1/U_1/U_1/memory[30][3] ,
         \U_1/U_1/U_1/memory[30][2] , \U_1/U_1/U_1/memory[30][1] ,
         \U_1/U_1/U_1/memory[30][0] , \U_1/U_1/U_1/memory[31][7] ,
         \U_1/U_1/U_1/memory[31][6] , \U_1/U_1/U_1/memory[31][5] ,
         \U_1/U_1/U_1/memory[31][4] , \U_1/U_1/U_1/memory[31][3] ,
         \U_1/U_1/U_1/memory[31][2] , \U_1/U_1/U_1/memory[31][1] ,
         \U_1/U_1/U_1/memory[31][0] , \U_1/U_1/U_1/opcode[0][1] ,
         \U_1/U_1/U_1/opcode[0][0] , \U_1/U_1/U_1/opcode[1][1] ,
         \U_1/U_1/U_1/opcode[1][0] , \U_1/U_1/U_1/opcode[2][1] ,
         \U_1/U_1/U_1/opcode[2][0] , \U_1/U_1/U_1/opcode[3][1] ,
         \U_1/U_1/U_1/opcode[3][0] , \U_1/U_1/U_1/opcode[4][1] ,
         \U_1/U_1/U_1/opcode[4][0] , \U_1/U_1/U_1/opcode[5][1] ,
         \U_1/U_1/U_1/opcode[5][0] , \U_1/U_1/U_1/opcode[6][1] ,
         \U_1/U_1/U_1/opcode[6][0] , \U_1/U_1/U_1/opcode[7][1] ,
         \U_1/U_1/U_1/opcode[7][0] , \U_1/U_1/U_1/opcode[8][1] ,
         \U_1/U_1/U_1/opcode[8][0] , \U_1/U_1/U_1/opcode[9][1] ,
         \U_1/U_1/U_1/opcode[9][0] , \U_1/U_1/U_1/opcode[10][1] ,
         \U_1/U_1/U_1/opcode[10][0] , \U_1/U_1/U_1/opcode[11][1] ,
         \U_1/U_1/U_1/opcode[11][0] , \U_1/U_1/U_1/opcode[12][1] ,
         \U_1/U_1/U_1/opcode[12][0] , \U_1/U_1/U_1/opcode[13][1] ,
         \U_1/U_1/U_1/opcode[13][0] , \U_1/U_1/U_1/opcode[14][1] ,
         \U_1/U_1/U_1/opcode[14][0] , \U_1/U_1/U_1/opcode[15][1] ,
         \U_1/U_1/U_1/opcode[15][0] , \U_1/U_1/U_1/opcode[16][1] ,
         \U_1/U_1/U_1/opcode[16][0] , \U_1/U_1/U_1/opcode[17][1] ,
         \U_1/U_1/U_1/opcode[17][0] , \U_1/U_1/U_1/opcode[18][1] ,
         \U_1/U_1/U_1/opcode[18][0] , \U_1/U_1/U_1/opcode[19][1] ,
         \U_1/U_1/U_1/opcode[19][0] , \U_1/U_1/U_1/opcode[20][1] ,
         \U_1/U_1/U_1/opcode[20][0] , \U_1/U_1/U_1/opcode[21][1] ,
         \U_1/U_1/U_1/opcode[21][0] , \U_1/U_1/U_1/opcode[22][1] ,
         \U_1/U_1/U_1/opcode[22][0] , \U_1/U_1/U_1/opcode[23][1] ,
         \U_1/U_1/U_1/opcode[23][0] , \U_1/U_1/U_1/opcode[24][1] ,
         \U_1/U_1/U_1/opcode[24][0] , \U_1/U_1/U_1/opcode[25][1] ,
         \U_1/U_1/U_1/opcode[25][0] , \U_1/U_1/U_1/opcode[26][1] ,
         \U_1/U_1/U_1/opcode[26][0] , \U_1/U_1/U_1/opcode[27][1] ,
         \U_1/U_1/U_1/opcode[27][0] , \U_1/U_1/U_1/opcode[28][1] ,
         \U_1/U_1/U_1/opcode[28][0] , \U_1/U_1/U_1/opcode[29][1] ,
         \U_1/U_1/U_1/opcode[29][0] , \U_1/U_1/U_1/opcode[30][1] ,
         \U_1/U_1/U_1/opcode[30][0] , \U_1/U_1/U_1/opcode[31][1] ,
         \U_1/U_1/U_1/opcode[31][0] , \U_1/U_1/U_1/N46 , \U_1/U_1/U_1/N45 ,
         \U_1/U_1/U_1/N44 , \U_1/U_1/U_1/N43 , \U_1/U_1/U_1/N36 ,
         \U_1/U_1/U_1/N35 , \U_1/U_1/U_1/N34 , \U_1/U_1/U_1/N33 ,
         \U_1/U_1/U_1/N32 , \U_1/U_1/U_1/state , \U_1/U_1/U_1/writeptr[0] ,
         \U_1/U_1/U_1/writeptr[1] , \U_1/U_1/U_1/writeptr[2] ,
         \U_1/U_1/U_1/writeptr[3] , \U_1/U_1/U_1/writeptr[4] ,
         \U_1/U_1/U_1/readptr[0] , \U_1/U_1/U_1/readptr[1] ,
         \U_1/U_1/U_1/readptr[2] , \U_1/U_1/U_1/readptr[3] ,
         \U_1/U_1/U_1/readptr[4] , \U_1/U_2/U_2/current_crc[0] ,
         \U_1/U_2/U_2/current_crc[1] , \U_1/U_2/U_2/current_crc[2] ,
         \U_1/U_2/U_2/current_crc[3] , \U_1/U_2/U_2/current_crc[4] ,
         \U_1/U_2/U_2/current_crc[5] , \U_1/U_2/U_2/current_crc[6] ,
         \U_1/U_2/U_2/current_crc[7] , \U_1/U_2/U_2/current_crc[8] ,
         \U_1/U_2/U_2/current_crc[9] , \U_1/U_2/U_2/current_crc[10] ,
         \U_1/U_2/U_2/current_crc[11] , \U_1/U_2/U_2/current_crc[12] ,
         \U_1/U_2/U_2/current_crc[13] , \U_1/U_2/U_2/current_crc[14] ,
         \U_1/U_2/U_2/current_crc[15] , \U_1/U_2/U_1/N32 , \U_1/U_2/U_1/N31 ,
         \U_1/U_2/U_1/N29 , \U_1/U_2/U_1/state[0] , \U_1/U_2/U_1/state[1] ,
         \U_1/U_2/U_1/state[2] , \U_1/U_2/U_1/state[3] ,
         \U_1/U_2/U_1/DP_hold2 , \U_1/U_2/U_1/DP_hold1 ,
         \U_1/U_2/U_0/DP_hold2 , \U_1/U_2/U_0/DP_hold1 , \U_1/U_2/U_5/N170 ,
         \U_1/U_2/U_5/curCRC_ERROR , \U_1/U_2/U_5/curR_ERROR ,
         \U_1/U_2/U_5/count[0] , \U_1/U_2/U_5/count[1] ,
         \U_1/U_2/U_5/count[2] , \U_1/U_2/U_5/count[3] ,
         \U_1/U_2/U_5/state[0] , \U_1/U_2/U_5/state[1] ,
         \U_1/U_2/U_5/state[2] , \U_1/U_2/U_5/state[3] , \U_1/U_2/U_7/state ,
         \U_1/U_2/U_7/count[0] , \U_1/U_2/U_7/count[1] ,
         \U_1/U_2/U_7/count[2] , \U_1/U_2/U_7/count[3] , \U_1/U_3/d_encode ,
         \U_1/U_3/SHIFT_ENABLE_E , \U_1/U_3/U_0/N59 , \U_1/U_3/U_0/dm_tx_nxt ,
         \U_1/U_3/U_0/DE_holdout_nxt , \U_1/U_3/U_0/DE_holdout_last ,
         \U_1/U_3/U_0/state[0] , \U_1/U_3/U_0/state[1] ,
         \U_1/U_3/U_0/state[2] , \U_1/U_3/U_0/state[3] ,
         \U_1/U_3/U_0/DE_holdout_BS , \U_1/U_3/U_0/DE_holdout ,
         \U_1/U_3/U_2/count[0] , \U_1/U_3/U_2/count[1] ,
         \U_1/U_3/U_2/count[2] , \U_1/U_3/U_3/N188 , \U_1/U_3/U_3/N187 ,
         \U_1/U_3/U_3/N90 , \U_1/U_3/U_3/N89 , \U_1/U_3/U_3/N88 ,
         \U_1/U_3/U_3/N87 , \U_1/U_3/U_3/N86 , \U_1/U_3/U_3/N85 ,
         \U_1/U_3/U_3/N84 , \U_1/U_3/U_3/N65 , \U_1/U_3/U_3/N64 ,
         \U_1/U_3/U_3/N63 , \U_1/U_3/U_3/N62 , \U_1/U_3/U_3/N61 ,
         \U_1/U_3/U_3/N60 , \U_1/U_3/U_3/N59 , \U_1/U_3/U_3/count[0] ,
         \U_1/U_3/U_3/count[1] , \U_1/U_3/U_3/count[2] ,
         \U_1/U_3/U_3/count[3] , \U_1/U_3/U_3/count[4] ,
         \U_1/U_3/U_3/count[5] , \U_1/U_3/U_3/state[0] ,
         \U_1/U_3/U_3/state[1] , \U_1/U_3/U_3/state[2] , \U_1/U_3/U_4/state ,
         \U_1/U_3/U_4/count[0] , \U_1/U_3/U_4/count[1] ,
         \U_1/U_3/U_4/count[2] , \U_1/U_3/U_4/count[3] , n177, n178, n179,
         n180, n182, n184, n185, n186, n187, n189, n190, n191, n193, n194,
         n196, n197, n198, n200, n201, n202, n204, n205, n206, n207, n209,
         n210, n211, n212, n214, n215, n216, n217, n219, n220, n221, n222,
         n224, n225, n226, n227, n228, n230, n231, n232, n236, n237, n238,
         n240, n243, n244, n245, n247, n248, n250, n251, n252, n254, n255,
         n257, n258, n259, n261, n262, n264, n265, n266, n268, n269, n271,
         n272, n273, n275, n276, n278, n279, n280, n282, n283, n285, n286,
         n287, n289, n290, n292, n293, n294, n296, n297, n298, n299, n300,
         n301, n303, n304, n306, n307, n308, n309, n310, n311, n312, n314,
         n315, n316, n317, n318, n320, n321, n322, n325, n326, n329, n333,
         n337, n341, n345, n349, n353, n357, n362, n364, n369, n371, n372,
         n374, n375, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n460, n463, n464, n465, n466,
         n468, n470, n471, n472, n473, n475, n477, n479, n480, n482, n483,
         n484, n485, n486, n487, n488, n490, n491, n492, n493, n495, n496,
         n497, n498, n500, n501, n502, n503, n505, n506, n507, n508, n510,
         n511, n512, n513, n514, n516, n517, n518, n519, n522, n523, n525,
         n528, n530, n532, n533, n535, n536, n538, n539, n541, n542, n544,
         n545, n547, n548, n550, n551, n553, n554, n555, n556, n557, n559,
         n560, n561, n562, n566, n567, n568, n569, n571, n574, n577, n580,
         n583, n586, n589, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n604, n607, n609, n610, n613, n617, n621,
         n625, n629, n633, n637, n641, n646, n648, n653, n655, n656, n658,
         n659, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n744, n747, n748, n749, n750, n753,
         n754, n756, n757, n758, n760, n761, n762, n763, n764, n767, n768,
         n770, n771, n772, n774, n776, n777, n781, n783, n784, n785, n786,
         n788, n790, n791, n792, n794, n796, n798, n800, n802, n804, n806,
         n808, n809, n812, n813, n814, n815, n818, n819, n820, n833, n834,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n852, n853, n854, n856, n857, n862, n864,
         n865, n867, n868, n869, n870, n871, n872, n873, n874, n875, n877,
         n879, n880, n881, n882, n884, n886, n888, n890, n892, n893, n895,
         n896, n898, n900, n902, n904, n906, n908, n910, n912, n913, n914,
         n916, n917, n918, n919, n921, n926, n931, n934, n935, n937, n939,
         n941, n943, n944, n945, n946, n947, n948, n949, n950, n951, n954,
         n956, n959, n962, n964, n966, n968, n970, n972, n974, n975, n977,
         n979, n980, n981, n984, n986, n988, n990, n992, n994, n996, n998,
         n1000, n1001, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1013, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1032, n1033, n1034, n1036,
         n1052, n1054, n1055, n1056, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1067, n1068, n1070, n1072, n1074, n1076, n1078, n1080,
         n1082, n1084, n1085, n1087, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1101, n1102, n1105, n1106, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1185,
         n1187, n1189, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1202, n1204, n1206, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1221, n1223, n1225,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1238, n1240, n1242, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1262, n1263, n1264,
         n1265, n1266, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1282,
         n1283, n1284, n1285, n1286, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1305, n1306, n1307, n1308, n1309, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1325, n1326, n1327, n1328,
         n1329, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1348, n1349, n1350, n1351, n1352, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1368, n1369, n1370, n1371, n1372, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1391, n1392,
         n1393, n1394, n1395, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1411, n1412, n1413, n1414, n1415, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1434, n1435, n1436, n1437, n1438,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1454, n1455, n1456,
         n1457, n1458, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1477, n1478, n1479, n1480, n1481, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1497, n1498, n1499, n1500, n1501, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1520,
         n1521, n1522, n1523, n1524, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1540, n1541, n1542, n1543, n1544, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1563, n1564, n1565, n1566,
         n1567, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1583, n1584,
         n1585, n1586, n1587, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1605, n1609, n1610, n1611, n1612, n1613, n1615,
         n1616, n1617, n1618, n1619, n1626, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1642, n1644, n1645, n1646, n1647, n1648, n1649,
         n1657, n1658, n1659, n1660, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1710, n1712, n1714, n1716, n1718, n1720, n1722, n1724, n1725, n1726,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1768, n1770, n1772, n1774,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1856, n1858, n1860, n1862, n1863, n1866, n1868, n1869,
         n1870, n1871, n1872, n1873, n1875, n1876, n1877, n1878, n1880, n1881,
         n1882, n1883, n1885, n1886, n1888, n1889, n1891, n1893, n1894, n1896,
         n1897, n1899, n1902, n1904, n1906, n1908, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1918, n1919, n1920, n1922, n1923, n1924, n1925,
         n1927, n1928, n1929, n1930, n1932, n1934, n1935, n1937, n1939, n1941,
         n1942, n1943, n1945, n1946, n1947, n1949, n1950, n1951, n1953, n1954,
         n1955, n1956, n1958, n1959, n1960, n1962, n1963, n1964, n1965, n1967,
         n1968, n1969, n1971, n1974, n1975, n1977, n1979, n1982, n1984, n1986,
         n1987, n1988, n1990, n1991, n1992, n1993, n1994, n1996, n1997, n1999,
         n2000, n2004, n2005, n2010, n2012, n2014, n2016, n2019, n2021, n2023,
         n2025, n2027, n2029, n2031, n2033, n2034, n2037, n2044, n2048, n2052,
         n2056, n2060, n2062, n2063, n2065, n2067, n2068, n2069, n2071, n2073,
         n2075, n2076, n2077, n2078, n2080, n2081, n2083, n2084, n2085, n2086,
         n2088, n2089, n2091, n2092, n2093, n2094, n2096, n2098, n2099, n2100,
         n2102, n2104, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2119, n2122, n2123, n2125, n2126, n2127, n2128, n2130,
         n2133, n2135, n2136, n2138, n2139, n2140, n2142, n2144, n2146, n2147,
         n2150, n2152, n2153, n2155, n2156, n2157, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2167, n2168, n2169, n2170, n2172, n2173, n2175,
         n2176, n2177, n2179, n2180, n2181, n2183, n2185, n2186, n2187, n2189,
         n2191, n2192, n2193, n2194, n2196, n2197, n2199, n2200, n2202, n2203,
         n2204, n2205, n2206, n2207, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2232, n2234, n2235, n2236, n2237,
         n2239, n2240, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2252, n2253, n2254, n2255, n2256, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2266, n2267, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2283, n2284, n2286, n2287,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2319, n2320,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2335, n2336, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2351, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2366, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2381, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2396, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2411, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2426, n2429, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2443, n2444, n2445,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2459, n2460, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2474, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2488, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2502, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2516, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2530, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2544, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2558, n2559, n2560, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2574, n2575, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2589, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2603, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2617, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2631,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2645, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2659, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2673, n2675, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2689, n2690,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2704, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2718, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2732, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2746, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2760,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2774, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2788, n2789, n2790, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2804, n2805, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2819, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2833, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2847, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2861, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2875, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2889, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2903, n2905, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2919, n2920, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2934, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2948, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2962, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2976, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2990, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3004, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3018, n3019, n3020, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3034, n3035, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3049, n3051, n3052,
         n3053, n3054, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3064,
         n3065, n3066, n3067, n3068, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3078, n3079, n3080, n3081, n3083, n3084, n3085, n3086, n3088,
         n3089, n3090, n3091, n3092, n3094, n3095, n3096, n3097, n3098, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3109, n3110, n3111,
         n3112, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3122, n3123,
         n3124, n3125, n3130, n3131, n3132, n3133, n3135, n3136, n3137, n3138,
         n3140, n3141, n3142, n3144, n3146, n3147, n3149, n3151, n3153, n3155,
         n3157, n3159, n3161, n3162, n3164, n3167, n3168, n3171, n3174, n3176,
         n3179, n3180, n3181, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3193, n3195, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3207, n3208, n3209, n3215, n3216, n3217, n3218, n3220, n3222,
         n3223, n3224, n3225, n3227, n3229, n3230, n3231, n3232, n3234, n3235,
         n3236, n3237, n3239, n3242, n3243, n3244, n3247, n3248, n3250, n3251,
         n3255, n3256, n3257, n3259, n3260, n3261, n3262, n3263, n3266, n3268,
         n3269, n3270, n3271, n3273, n3274, n3275, n3276, n3277, n3279, n3280,
         n3281, n3283, n3285, n3287, n3289, n3291, n3293, n3295, n3296, n3297,
         n3298, n3299, n3300, n3303, n3305, n3306, n3307, n3308, n3310, n3312,
         n3313, n3314, n3316, n3318, n3320, n3322, n3324, n3326, n3328, n3330,
         n3331, n3334, n3335, n3336, n3337, n3340, n3341, n3342, n3355, n3356,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3374, n3375, n3376, n3378, n3379,
         n3384, n3386, n3387, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3400, n3402, n3403, n3404, n3405, n3407, n3409,
         n3411, n3413, n3415, n3418, n3419, n3421, n3423, n3425, n3427, n3429,
         n3431, n3433, n3434, n3436, n3437, n3438, n3440, n3441, n3442, n3443,
         n3444, n3447, n3448, n3450, n3452, n3454, n3456, n3460, n3461, n3464,
         n3468, n3469, n3470, n3471, n3472, n3473, n3475, n3476, n3477, n3480,
         n3481, n3483, n3485, n3487, n3489, n3491, n3493, n3495, n3496, n3497,
         n3498, n3500, n3501, n3502, n3503, n3504, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3518, n3522, n3523, n3525,
         n3527, n3529, n3531, n3533, n3535, n3537, n3538, n3541, n3542, n3543,
         n3545, n3547, n3549, n3551, n3553, n3555, n3557, n3558, n3559, n3561,
         n3562, n3563, n3565, n3566, n3569, n3570, n3571, n3572, n3573, n3574,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3589, n3590, n3591, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3654, n3655, n3656, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3688, n3690, n3692, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3705, n3707, n3709, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3724, n3726, n3728, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3741, n3743, n3745, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3765, n3766, n3767, n3768, n3769, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3785, n3786, n3787, n3788, n3789, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3808, n3809,
         n3810, n3811, n3812, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3828, n3829, n3830, n3831, n3832, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3851, n3852, n3853, n3854, n3855,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3871, n3872, n3873,
         n3874, n3875, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3894, n3895, n3896, n3897, n3898, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3914, n3915, n3916, n3917, n3918, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3937,
         n3938, n3939, n3940, n3941, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3957, n3958, n3959, n3960, n3961, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3980, n3981, n3982, n3983,
         n3984, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n4000, n4001,
         n4002, n4003, n4004, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4023, n4024, n4025, n4026, n4027, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4043, n4044, n4045, n4046, n4047,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4066, n4067, n4068, n4069, n4070, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4086, n4087, n4088, n4089, n4090, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4108, n4112, n4113,
         n4114, n4115, n4116, n4118, n4119, n4120, n4121, n4122, n4129, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4145, n4147, n4148,
         n4149, n4150, n4151, n4152, n4160, n4161, n4162, n4163, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4213, n4215, n4217, n4219, n4221, n4223,
         n4225, n4227, n4228, n4229, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4271, n4273, n4275, n4277, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4359, n4361, n4363, n4365,
         n4366, n4369, n4371, n4372, n4373, n4374, n4375, n4376, n4378, n4379,
         n4380, n4381, n4383, n4384, n4385, n4386, n4388, n4389, n4391, n4392,
         n4394, n4396, n4397, n4399, n4400, n4402, n4405, n4407, n4409, n4411,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4421, n4422, n4423,
         n4425, n4426, n4427, n4428, n4430, n4431, n4432, n4433, n4435, n4437,
         n4438, n4440, n4442, n4444, n4445, n4446, n4448, n4449, n4450, n4452,
         n4453, n4454, n4456, n4457, n4458, n4459, n4461, n4462, n4463, n4465,
         n4466, n4467, n4468, n4470, n4471, n4472, n4474, n4477, n4478, n4480,
         n4482, n4485, n4487, n4489, n4490, n4491, n4493, n4494, n4495, n4496,
         n4497, n4499, n4500, n4501, n4502, n4505, n4511, n4513, n4515, n4517,
         n4520, n4522, n4524, n4526, n4528, n4530, n4532, n4534, n4535, n4538,
         n4545, n4549, n4553, n4557, n4561, n4563, n4564, n4566, n4568, n4569,
         n4570, n4572, n4574, n4576, n4577, n4578, n4579, n4581, n4582, n4584,
         n4585, n4586, n4587, n4589, n4590, n4592, n4593, n4594, n4595, n4597,
         n4599, n4600, n4601, n4603, n4605, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4620, n4623, n4624, n4626, n4627,
         n4628, n4629, n4631, n4634, n4636, n4637, n4639, n4640, n4641, n4643,
         n4645, n4647, n4648, n4651, n4653, n4654, n4656, n4657, n4658, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4668, n4669, n4670, n4671,
         n4673, n4674, n4676, n4677, n4678, n4680, n4681, n4682, n4684, n4686,
         n4687, n4688, n4690, n4692, n4693, n4694, n4695, n4697, n4698, n4700,
         n4701, n4703, n4704, n4705, n4706, n4707, n4708, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4733, n4735,
         n4736, n4737, n4738, n4740, n4741, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4753, n4754, n4755, n4756, n4757, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4767, n4768, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4784,
         n4785, n4787, n4788, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4820, n4821, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4836, n4837, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4852, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4867,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4882, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4897, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4912, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4927, n4930, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4944, n4945, n4946, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4960, n4961, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4975, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4989,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5003, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5017, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5031, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5045, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5059,
         n5060, n5061, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5075, n5076, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5090, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5104, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5118, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5132, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5146, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5160, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5174, n5176,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5190, n5191, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5205, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5219, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5233, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5247, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5261, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5275, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5289, n5290, n5291, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5305, n5306, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5320, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5334, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5348, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5362,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5376, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5390, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5404, n5406, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5420, n5421,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5435, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5449, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5463, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5477, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5491,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5505, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5519, n5520, n5521, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5535, n5536, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5550, n5552, n5553, n5554, n5555, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5565, n5566, n5567, n5568, n5569, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5579, n5580, n5581, n5582, n5584, n5585,
         n5586, n5587, n5589, n5590, n5591, n5592, n5593, n5595, n5596, n5597,
         n5598, n5599, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5610, n5611, n5612, n5613, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5623, n5624, n5625, n5626, n5631, n5632, n5633, n5634, n5636,
         n5637, n5638, n5639, n5641, n5642, n5643, n5645, n5647, n5648, n5650,
         n5652, n5654, n5656, n5658, n5660, n5662, n5663, n5665, n5668, n5669,
         n5672, n5675, n5677, n5680, n5681, n5682, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5694, n5696, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5708, n5709, n5710, n5716, n5717, n5718,
         n5719, n5721, n5723, n5724, n5725, n5726, n5728, n5730, n5731, n5732,
         n5733, n5735, n5736, n5737, n5738, n5740, n5743, n5744, n5745, n5748,
         n5749, n5751, n5752, n5755, n5756, n5757, n5759, n5760, n5761, n5762,
         n5763, n5766, n5768, n5769, n5770, n5771, n5773, n5774, n5775, n5776,
         n5777, n5779, n5780, n5781, n5783, n5785, n5787, n5789, n5791, n5793,
         n5795, n5796, n5797, n5798, n5799, n5800, n5803, n5804, n5805, n5806,
         n5808, n5810, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5825, n5827, n5828, n5829, n5831, n5832, n5834,
         n5835, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5849, n5850, n5851, n5852, n5854, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5876, n5877, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5888, n5889, n5890, n5892, n5893, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5911, n5912, n5913, n5914, n5915, n5916, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5927, n5928, n5929, n5930, n5931, n5932, n5934,
         n5935, n5937, n5938, n5941, n5942, n5943, n5944, n5945, n5947, n5948,
         n5949, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5963, n5964, n5965, n5966, n5968, n5969, n5970, n5972, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5982, n5983, n5984, n5985,
         n5986, n5989, n5991, n5992, n5994, n5995, n5996, n5997, n6000, n6001,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6014, n6016,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6027, n6028,
         n6029, n6031, n6032, n6033, n6034, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6049, n6050, n6051, n6052, n6054,
         n6055, n6056, n6058, n6059, n6060, n6061, n6063, n6065, n6066, n6067,
         n6069, n6070, n6071, n6073, n6074, n6075, n6077, n6078, n6079, n6081,
         n6082, n6083, n6085, n6086, n6087, n6089, n6090, n6091, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6152, n6153, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6165, n6166, n6167, n6168, n6170,
         n6171, n6172, n6173, n6174, n6175, n6177, n6178, n6180, n6181, n6182,
         n6183, n6184, n6185, n6187, n6188, n6189, n6191, n6192, n6193, n6194,
         n6196, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6215, n6216, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6229, n6230,
         n6231, n6232, n6234, n6236, n6237, n6238, n6240, n6241, n6242, n6243,
         n6247, n6248, n6250, n6251, n6253, n6254, n6256, n6257, n6259, n6260,
         n6262, n6263, n6265, n6266, n6268, n6269, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6280, n6282, n6283, n6284, n6287, n6288,
         n6289, n6290, n6291, n6293, n6294, n6296, n6298, n6303, n6304, n6305,
         n6306, n6307, n6311, n6312, n6313, n6314, n6315, n6319, n6320, n6321,
         n6322, n6323, n6327, n6328, n6329, n6330, n6331, n6336, n6337, n6338,
         n6339, n6340, n6345, n6346, n6347, n6348, n6349, n6354, n6355, n6356,
         n6357, n6358, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6372, n6374, n6377, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6389, n6391, n6392, n6393, n6395, n6396, n6398, n6399,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6413,
         n6414, n6415, n6416, n6418, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6440, n6441, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6452,
         n6453, n6454, n6456, n6457, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6475,
         n6476, n6477, n6478, n6479, n6480, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6491, n6492, n6493, n6494, n6495, n6496, n6498, n6499,
         n6501, n6502, n6505, n6506, n6507, n6508, n6509, n6511, n6512, n6513,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6527, n6528, n6529, n6530, n6532, n6533, n6534, n6536, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6546, n6547, n6548, n6549, n6550,
         n6553, n6555, n6556, n6558, n6559, n6560, n6561, n6564, n6565, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6578, n6580, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6591, n6592, n6593,
         n6595, n6596, n6597, n6598, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6613, n6614, n6615, n6616, n6618, n6619,
         n6620, n6622, n6623, n6624, n6625, n6626, n6627, n6630, n6631, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6658, n6660, n6661, n6662, n6663, n6664, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6717, n6718,
         n6719, n6721, n6722, n6723, n6724, n6725, n6727, n6728, n6729, n6731,
         n6732, n6735, n6736, n6737, n6739, n6740, n6741, n6742, n6743, n6745,
         n6746, n6747, n6748, n6749, n6751, n6753, n6754, n6756, n6757, n6758,
         n6759, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6774, n6775, n6776, n6777, n6778, n6779, n6781,
         n6782, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6793, n6794,
         n6795, n6797, n6799, n6800, n6801, n6803, n6804, n6806, n6807, n6808,
         n6810, n6811, n6813, n6814, n6816, n6817, n6819, n6820, n6822, n6823,
         n6825, n6826, n6828, n6829, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6839, n6840, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6850, n6851, n6853, n6855, n6860, n6861, n6862, n6863, n6864, n6868,
         n6869, n6870, n6871, n6872, n6876, n6877, n6878, n6879, n6880, n6884,
         n6885, n6886, n6887, n6888, n6893, n6894, n6895, n6896, n6897, n6902,
         n6903, n6904, n6905, n6906, n6911, n6912, n6913, n6914, n6915, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6998, n7017, n7020, n7023, n7026, n7029,
         n7032, n7035, n7038, n7041, n7044, n7047, n7050, n7053, n7056, n7074,
         n7075, n7076, n7077, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7130, n7140, n7207, n7267, n7268, n7269, n7270,
         n7274, n7277, n7280, n7283, n7286, n7289, n7295, n7299, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7390, n7392, n7394,
         n7396, n7398, n7400, n7402, n7404, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7461, n7462, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7522, n7532, n7599, n7659, n7660, n7661, n7662,
         n7666, n7669, n7672, n7675, n7678, n7681, n7687, n7691, n7748, n7749,
         n7750, n7751, n7754, n7756, n7757, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7869, n7870,
         n7871, n7872, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8564, n8565,
         n8566, n8567, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, \U_0/U_0/U_0/N456 , \U_0/U_0/U_0/N455 ,
         \U_0/U_0/U_0/N454 , \U_0/U_0/U_0/N453 , \U_0/U_0/U_0/N452 ,
         \U_0/U_0/U_0/N451 , \U_0/U_0/U_0/N450 , \U_0/U_0/U_0/N449 ,
         \U_1/U_0/U_0/N456 , \U_1/U_0/U_0/N455 , \U_1/U_0/U_0/N454 ,
         \U_1/U_0/U_0/N453 , \U_1/U_0/U_0/N452 , \U_1/U_0/U_0/N451 ,
         \U_1/U_0/U_0/N450 , \U_1/U_0/U_0/N449 ,
         \U_1/U_1/U_1/add_76_aco/carry[4] , \U_1/U_1/U_1/add_76_aco/carry[3] ,
         \U_1/U_1/U_1/add_76_aco/carry[2] , \U_1/U_1/U_1/add_76_aco/carry[1] ,
         \U_1/U_1/U_1/sub_72/carry[4] , \U_1/U_1/U_1/sub_72/carry[3] ,
         \U_1/U_1/U_1/sub_72/carry[2] , \U_1/U_1/U_1/sub_72/carry[1] ,
         \U_1/U_1/U_1/add_67/carry[4] , \U_1/U_1/U_1/add_67/carry[3] ,
         \U_1/U_1/U_1/add_67/carry[2] , \U_1/U_0/U_1/U_2/add_46/carry[7] ,
         \U_1/U_0/U_1/U_2/add_46/carry[6] , \U_1/U_0/U_1/U_2/add_46/carry[5] ,
         \U_1/U_0/U_1/U_2/add_46/carry[4] , \U_1/U_0/U_1/U_2/add_46/carry[3] ,
         \U_0/U_1/U_1/add_76_aco/carry[4] , \U_0/U_1/U_1/add_76_aco/carry[3] ,
         \U_0/U_1/U_1/add_76_aco/carry[2] , \U_0/U_1/U_1/add_76_aco/carry[1] ,
         \U_0/U_1/U_1/sub_72/carry[4] , \U_0/U_1/U_1/sub_72/carry[3] ,
         \U_0/U_1/U_1/sub_72/carry[2] , \U_0/U_1/U_1/sub_72/carry[1] ,
         \U_0/U_1/U_1/add_67/carry[4] , \U_0/U_1/U_1/add_67/carry[3] ,
         \U_0/U_1/U_1/add_67/carry[2] , \U_0/U_0/U_1/U_2/add_46/carry[7] ,
         \U_0/U_0/U_1/U_2/add_46/carry[6] , \U_0/U_0/U_1/U_2/add_46/carry[5] ,
         \U_0/U_0/U_1/U_2/add_46/carry[4] , \U_0/U_0/U_1/U_2/add_46/carry[3] ,
         \r2042/carry[6] , \r2042/carry[5] , \r2042/carry[4] ,
         \r2042/carry[3] , \r2042/carry[2] , \r2042/carry[1] ,
         \r2028/carry[4] , \r2028/carry[3] , \r2028/carry[2] ,
         \r2008/carry[6] , \r2008/carry[5] , \r2008/carry[4] ,
         \r2008/carry[3] , \r2008/carry[2] , \r2008/carry[1] ,
         \r1994/carry[4] , \r1994/carry[3] , \r1994/carry[2] , n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9560, n9561, n9562, n9563, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077;
  wire   [7:0] \U_0/RCV_DATA ;
  wire   [7:0] \U_0/PROCESSED_DATA ;
  wire   [7:0] \U_0/PRGA_IN ;
  wire   [63:0] \U_0/U_0/PLAINKEY ;
  wire   [7:0] \U_0/U_0/U_0/fdata ;
  wire   [7:0] \U_0/U_0/U_0/faddr ;
  wire   [7:0] \U_0/U_0/U_0/delaydata ;
  wire   [4:0] \U_0/U_0/U_0/nextState ;
  wire   [7:0] \U_0/U_0/U_0/currentProcessedData ;
  wire   [1:0] \U_0/U_0/U_1/STOP_DATA ;
  wire   [7:0] \U_0/U_0/U_1/RCV_DATA ;
  wire   [7:0] \U_0/U_0/U_1/LOAD_DATA ;
  wire   [7:0] \U_0/U_0/U_1/U_2/nextCount ;
  wire   [1:0] \U_0/U_1/OUT_OPCODE ;
  wire   [7:0] \U_0/U_1/DATA ;
  wire   [4:0] \U_0/U_1/BYTE_COUNT ;
  wire   [1:0] \U_0/U_1/U_0/tempOpcode ;
  wire   [7:0] \U_0/U_1/U_0/tempData ;
  wire   [2:0] \U_0/U_1/U_0/nextState ;
  wire   [15:0] \U_0/U_2/rx_CHECK_CRC ;
  wire   [15:0] \U_0/U_2/RX_CRC ;
  wire   [15:0] \U_0/U_2/U_2/cache_1 ;
  wire   [3:0] \U_0/U_2/U_5/nextstate ;
  wire   [3:0] \U_0/U_2/U_7/nextcount ;
  wire   [7:0] \U_0/U_3/send_data ;
  wire   [15:0] \U_0/U_3/TX_CRC ;
  wire   [3:0] \U_0/U_3/U_0/nextstate ;
  wire   [7:1] \U_0/U_3/U_2/present_val ;
  wire   [7:0] \U_0/U_3/U_3/current_send_data ;
  wire   [7:0] \U_0/U_3/U_3/flop_data ;
  wire   [2:0] \U_0/U_3/U_3/nextstate ;
  wire   [3:0] \U_0/U_3/U_4/nextcount ;
  wire   [7:0] \U_1/RCV_DATA ;
  wire   [7:0] \U_1/PROCESSED_DATA ;
  wire   [7:0] \U_1/PRGA_IN ;
  wire   [63:0] \U_1/U_0/PLAINKEY ;
  wire   [7:0] \U_1/U_0/U_0/fdata ;
  wire   [7:0] \U_1/U_0/U_0/faddr ;
  wire   [7:0] \U_1/U_0/U_0/delaydata ;
  wire   [4:0] \U_1/U_0/U_0/nextState ;
  wire   [7:0] \U_1/U_0/U_0/currentProcessedData ;
  wire   [1:0] \U_1/U_0/U_1/STOP_DATA ;
  wire   [7:0] \U_1/U_0/U_1/RCV_DATA ;
  wire   [7:0] \U_1/U_0/U_1/LOAD_DATA ;
  wire   [7:0] \U_1/U_0/U_1/U_2/nextCount ;
  wire   [1:0] \U_1/U_1/OUT_OPCODE ;
  wire   [7:0] \U_1/U_1/DATA ;
  wire   [4:0] \U_1/U_1/BYTE_COUNT ;
  wire   [1:0] \U_1/U_1/U_0/tempOpcode ;
  wire   [7:0] \U_1/U_1/U_0/tempData ;
  wire   [2:0] \U_1/U_1/U_0/nextState ;
  wire   [15:0] \U_1/U_2/rx_CHECK_CRC ;
  wire   [15:0] \U_1/U_2/RX_CRC ;
  wire   [15:0] \U_1/U_2/U_2/cache_1 ;
  wire   [3:0] \U_1/U_2/U_5/nextstate ;
  wire   [3:0] \U_1/U_2/U_7/nextcount ;
  wire   [7:0] \U_1/U_3/send_data ;
  wire   [15:0] \U_1/U_3/TX_CRC ;
  wire   [3:0] \U_1/U_3/U_0/nextstate ;
  wire   [7:1] \U_1/U_3/U_2/present_val ;
  wire   [7:0] \U_1/U_3/U_3/current_send_data ;
  wire   [7:0] \U_1/U_3/U_3/flop_data ;
  wire   [2:0] \U_1/U_3/U_3/nextstate ;
  wire   [3:0] \U_1/U_3/U_4/nextcount ;
  tri   \U_0/U_0/U_0/nfdata[0] ;
  tri   \U_0/U_0/U_0/nfdata[1] ;
  tri   \U_0/U_0/U_0/nfdata[2] ;
  tri   \U_0/U_0/U_0/nfdata[3] ;
  tri   \U_0/U_0/U_0/nfdata[4] ;
  tri   \U_0/U_0/U_0/nfdata[5] ;
  tri   \U_0/U_0/U_0/nfdata[6] ;
  tri   \U_0/U_0/U_0/nfdata[7] ;
  tri   \U_0/U_0/U_0/nfaddr[0] ;
  tri   \U_0/U_0/U_0/nfaddr[1] ;
  tri   \U_0/U_0/U_0/nfaddr[2] ;
  tri   \U_0/U_0/U_0/nfaddr[3] ;
  tri   \U_0/U_0/U_0/nfaddr[4] ;
  tri   \U_0/U_0/U_0/nfaddr[5] ;
  tri   \U_0/U_0/U_0/nfaddr[6] ;
  tri   \U_0/U_0/U_0/nfaddr[7] ;
  tri   \U_1/U_0/U_0/nfdata[0] ;
  tri   \U_1/U_0/U_0/nfdata[1] ;
  tri   \U_1/U_0/U_0/nfdata[2] ;
  tri   \U_1/U_0/U_0/nfdata[3] ;
  tri   \U_1/U_0/U_0/nfdata[4] ;
  tri   \U_1/U_0/U_0/nfdata[5] ;
  tri   \U_1/U_0/U_0/nfdata[6] ;
  tri   \U_1/U_0/U_0/nfdata[7] ;
  tri   \U_1/U_0/U_0/nfaddr[0] ;
  tri   \U_1/U_0/U_0/nfaddr[1] ;
  tri   \U_1/U_0/U_0/nfaddr[2] ;
  tri   \U_1/U_0/U_0/nfaddr[3] ;
  tri   \U_1/U_0/U_0/nfaddr[4] ;
  tri   \U_1/U_0/U_0/nfaddr[5] ;
  tri   \U_1/U_0/U_0/nfaddr[6] ;
  tri   \U_1/U_0/U_0/nfaddr[7] ;

  DFFSR \U_0/U_0/U_1/U_0/Q_int_reg  ( .D(SERIAL_IN), .CLK(CLK), .R(n9500), .S(
        1'b1), .Q(\U_0/U_0/U_1/U_0/Q_int ) );
  DFFSR \U_0/U_0/U_1/U_0/Q_int2_reg  ( .D(\U_0/U_0/U_1/U_0/Q_int ), .CLK(CLK), 
        .R(n9489), .S(1'b1), .Q(\U_0/U_0/U_1/U_0/Q_int2 ) );
  DFFSR \U_0/U_0/U_1/U_7/nextState_reg[7]  ( .D(n9162), .CLK(CLK), .R(n9506), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_7/nextState[7] ) );
  DFFSR \U_0/U_0/U_1/U_7/state_reg[7]  ( .D(\U_0/U_0/U_1/U_7/nextState[7] ), 
        .CLK(CLK), .R(n9499), .S(1'b1), .Q(\U_0/U_0/U_1/U_7/state[7] ) );
  DFFSR \U_0/U_0/U_1/U_7/nextState_reg[6]  ( .D(n9161), .CLK(CLK), .R(n9499), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_7/nextState[6] ) );
  DFFSR \U_0/U_0/U_1/U_7/state_reg[6]  ( .D(\U_0/U_0/U_1/U_7/nextState[6] ), 
        .CLK(CLK), .R(n9499), .S(1'b1), .Q(\U_0/U_0/U_1/U_7/state[6] ) );
  DFFSR \U_0/U_0/U_1/U_7/nextState_reg[5]  ( .D(n9160), .CLK(CLK), .R(n9499), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_7/nextState[5] ) );
  DFFSR \U_0/U_0/U_1/U_7/state_reg[5]  ( .D(\U_0/U_0/U_1/U_7/nextState[5] ), 
        .CLK(CLK), .R(n9499), .S(1'b1), .Q(\U_0/U_0/U_1/U_7/state[5] ) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[9]  ( .D(n9154), .CLK(CLK), .R(n9499), 
        .S(1'b1), .Q(\U_0/U_0/U_1/STOP_DATA [1]) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[8]  ( .D(n9153), .CLK(CLK), .R(n9499), 
        .S(1'b1), .Q(\U_0/U_0/U_1/STOP_DATA [0]) );
  DFFSR \U_0/U_0/U_1/U_5/SB_DETECT_reg  ( .D(\U_0/U_0/U_1/U_5/sb_detect_flag ), 
        .CLK(CLK), .R(n9499), .S(1'b1), .Q(\U_0/U_0/U_1/SB_DETECT ) );
  DFFSR \U_0/U_0/U_1/U_2/state_reg[0]  ( .D(\U_0/U_0/U_1/U_2/nextState[0] ), 
        .CLK(CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/state[0] ) );
  DFFSR \U_0/U_0/U_1/U_2/timerRunning_reg  ( .D(n9152), .CLK(CLK), .R(n9500), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_2/timerRunning ) );
  DFFSR \U_0/U_0/U_1/U_2/nextCount_reg[1]  ( .D(\U_0/U_0/U_1/U_2/N32 ), .CLK(
        CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/nextCount [1]) );
  DFFSR \U_0/U_0/U_1/U_2/count_reg[1]  ( .D(\U_0/U_0/U_1/U_2/nextCount [1]), 
        .CLK(CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/count[1] ) );
  DFFSR \U_0/U_0/U_1/U_2/nextCount_reg[0]  ( .D(\U_0/U_0/U_1/U_2/N31 ), .CLK(
        CLK), .R(1'b1), .S(n9521), .Q(\U_0/U_0/U_1/U_2/nextCount [0]) );
  DFFSR \U_0/U_0/U_1/U_2/count_reg[0]  ( .D(\U_0/U_0/U_1/U_2/nextCount [0]), 
        .CLK(CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/N23 ) );
  DFFSR \U_0/U_0/U_1/U_2/nextCount_reg[2]  ( .D(\U_0/U_0/U_1/U_2/N33 ), .CLK(
        CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/nextCount [2]) );
  DFFSR \U_0/U_0/U_1/U_2/count_reg[2]  ( .D(\U_0/U_0/U_1/U_2/nextCount [2]), 
        .CLK(CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/count[2] ) );
  DFFSR \U_0/U_0/U_1/U_2/nextCount_reg[3]  ( .D(\U_0/U_0/U_1/U_2/N34 ), .CLK(
        CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/nextCount [3]) );
  DFFSR \U_0/U_0/U_1/U_2/count_reg[3]  ( .D(\U_0/U_0/U_1/U_2/nextCount [3]), 
        .CLK(CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/count[3] ) );
  DFFSR \U_0/U_0/U_1/U_2/nextCount_reg[4]  ( .D(\U_0/U_0/U_1/U_2/N35 ), .CLK(
        CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/nextCount [4]) );
  DFFSR \U_0/U_0/U_1/U_2/count_reg[4]  ( .D(\U_0/U_0/U_1/U_2/nextCount [4]), 
        .CLK(CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/count[4] ) );
  DFFSR \U_0/U_0/U_1/U_2/nextCount_reg[5]  ( .D(\U_0/U_0/U_1/U_2/N36 ), .CLK(
        CLK), .R(n9500), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/nextCount [5]) );
  DFFSR \U_0/U_0/U_1/U_2/count_reg[5]  ( .D(\U_0/U_0/U_1/U_2/nextCount [5]), 
        .CLK(CLK), .R(n9501), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/count[5] ) );
  DFFSR \U_0/U_0/U_1/U_2/nextCount_reg[6]  ( .D(\U_0/U_0/U_1/U_2/N37 ), .CLK(
        CLK), .R(n9501), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/nextCount [6]) );
  DFFSR \U_0/U_0/U_1/U_2/count_reg[6]  ( .D(\U_0/U_0/U_1/U_2/nextCount [6]), 
        .CLK(CLK), .R(n9501), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/count[6] ) );
  DFFSR \U_0/U_0/U_1/U_2/nextCount_reg[7]  ( .D(\U_0/U_0/U_1/U_2/N38 ), .CLK(
        CLK), .R(n9501), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/nextCount [7]) );
  DFFSR \U_0/U_0/U_1/U_2/count_reg[7]  ( .D(\U_0/U_0/U_1/U_2/nextCount [7]), 
        .CLK(CLK), .R(n9501), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/count[7] ) );
  DFFSR \U_0/U_0/U_1/U_2/state_reg[1]  ( .D(\U_0/U_0/U_1/U_2/nextState[1] ), 
        .CLK(CLK), .R(n9501), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/state[1] ) );
  DFFSR \U_0/U_0/U_1/U_2/state_reg[2]  ( .D(\U_0/U_0/U_1/U_2/nextState[2] ), 
        .CLK(CLK), .R(n9501), .S(1'b1), .Q(\U_0/U_0/U_1/U_2/state[2] ) );
  DFFSR \U_0/U_0/U_1/U_2/RBUF_LOAD_reg  ( .D(n9149), .CLK(CLK), .R(n9501), .S(
        1'b1), .Q(\U_0/U_0/U_1/RBUF_LOAD ) );
  DFFSR \U_0/U_0/U_1/U_2/SET_RBUF_FULL_reg  ( .D(n9146), .CLK(CLK), .R(n9501), 
        .S(1'b1), .Q(\U_0/U_0/U_1/SET_RBUF_FULL ) );
  DFFSR \U_0/U_0/U_1/U_2/CHK_ERROR_reg  ( .D(n9150), .CLK(CLK), .R(n9501), .S(
        1'b1), .Q(\U_0/U_0/U_1/CHK_ERROR ) );
  DFFSR \U_0/U_0/U_1/U_2/SBC_CLR_reg  ( .D(n9147), .CLK(CLK), .R(n9501), .S(
        1'b1), .Q(\U_0/U_0/U_1/SBC_CLR ) );
  DFFSR \U_0/U_0/U_1/U_2/TIMER_TRIG_reg  ( .D(n9148), .CLK(CLK), .R(n9501), 
        .S(1'b1), .Q(\U_0/U_0/U_1/TIMER_TRIG ) );
  DFFSR \U_0/U_0/U_1/U_7/nextState_reg[0]  ( .D(n9155), .CLK(CLK), .R(n9502), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_7/nextState[0] ) );
  DFFSR \U_0/U_0/U_1/U_7/state_reg[0]  ( .D(\U_0/U_0/U_1/U_7/nextState[0] ), 
        .CLK(CLK), .R(n9502), .S(1'b1), .Q(\U_0/U_0/U_1/U_7/state[0] ) );
  DFFSR \U_0/U_0/U_1/U_7/nextState_reg[1]  ( .D(n9156), .CLK(CLK), .R(n9502), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_7/nextState[1] ) );
  DFFSR \U_0/U_0/U_1/U_7/state_reg[1]  ( .D(\U_0/U_0/U_1/U_7/nextState[1] ), 
        .CLK(CLK), .R(n9502), .S(1'b1), .Q(\U_0/U_0/U_1/U_7/state[1] ) );
  DFFSR \U_0/U_0/U_1/U_7/nextState_reg[2]  ( .D(n9157), .CLK(CLK), .R(n9502), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_7/nextState[2] ) );
  DFFSR \U_0/U_0/U_1/U_7/state_reg[2]  ( .D(\U_0/U_0/U_1/U_7/nextState[2] ), 
        .CLK(CLK), .R(n9502), .S(1'b1), .Q(\U_0/U_0/U_1/U_7/state[2] ) );
  DFFSR \U_0/U_0/U_1/U_7/nextState_reg[3]  ( .D(n9158), .CLK(CLK), .R(n9502), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_7/nextState[3] ) );
  DFFSR \U_0/U_0/U_1/U_7/state_reg[3]  ( .D(\U_0/U_0/U_1/U_7/nextState[3] ), 
        .CLK(CLK), .R(n9502), .S(1'b1), .Q(\U_0/U_0/U_1/U_7/state[3] ) );
  DFFSR \U_0/U_0/U_1/U_7/nextState_reg[4]  ( .D(n9159), .CLK(CLK), .R(n9502), 
        .S(1'b1), .Q(\U_0/U_0/U_1/U_7/nextState[4] ) );
  DFFSR \U_0/U_0/U_1/U_7/state_reg[4]  ( .D(\U_0/U_0/U_1/U_7/nextState[4] ), 
        .CLK(CLK), .R(n9502), .S(1'b1), .Q(\U_0/U_0/U_1/U_7/state[4] ) );
  DFFSR \U_0/U_0/U_1/U_2/SBC_EN_reg  ( .D(n9151), .CLK(CLK), .R(n9502), .S(
        1'b1), .Q(\U_0/U_0/U_1/SBC_EN ) );
  DFFSR \U_0/U_0/U_1/U_5/SBE_reg  ( .D(\U_0/U_0/U_1/U_5/SBE_prime ), .CLK(CLK), 
        .R(n9502), .S(1'b1), .Q(\U_0/U_0/U_1/SBE ) );
  DFFSR \U_0/U_0/U_1/U_8/state_reg[0]  ( .D(n9144), .CLK(CLK), .R(n9503), .S(
        1'b1), .Q(\U_0/U_0/U_1/U_8/state[0] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/keyCount_reg[1]  ( .D(n9140), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/keyCount[1] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/keyCount_reg[2]  ( .D(n9139), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/keyCount[2] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/keyCount_reg[3]  ( .D(n9138), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/keyCount[3] ) );
  DFFSR \U_0/U_0/U_1/U_8/state_reg[2]  ( .D(n9145), .CLK(CLK), .R(n9503), .S(
        1'b1), .Q(\U_0/U_0/U_1/U_8/state[2] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/keyCount_reg[0]  ( .D(n9141), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/keyCount[0] ) );
  DFFSR \U_0/U_0/U_1/U_8/state_reg[3]  ( .D(n9143), .CLK(CLK), .R(n9503), .S(
        1'b1), .Q(\U_0/U_0/U_1/U_8/state[3] ) );
  DFFSR \U_0/U_0/U_1/U_8/state_reg[1]  ( .D(n9142), .CLK(CLK), .R(n9503), .S(
        1'b1), .Q(\U_0/U_0/U_1/U_8/state[1] ) );
  DFFSR \U_0/U_0/U_1/U_4/Q_int_reg  ( .D(n7691), .CLK(CLK), .R(n7748), .S(1'b1), .Q(\U_0/RBUF_FULL ) );
  DFFSR \U_0/U_0/U_1/U_1/OE_reg  ( .D(\U_0/U_0/U_1/U_1/OE_prime ), .CLK(CLK), 
        .R(n9503), .S(1'b1), .Q(\U_0/U_0/U_1/OE ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/address_reg[0]  ( .D(n9130), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/address[0] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/address_reg[1]  ( .D(n9131), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/address[1] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/address_reg[2]  ( .D(n9132), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/address[2] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/address_reg[6]  ( .D(n9136), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/address[6] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/address_reg[7]  ( .D(n9137), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/address[7] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/address_reg[3]  ( .D(n9133), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/address[3] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/address_reg[5]  ( .D(n9135), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/address[5] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/address_reg[4]  ( .D(n9134), .CLK(CLK), .Q(
        \U_0/U_0/U_1/U_8/address[4] ) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[7]  ( .D(n9129), .CLK(CLK), .R(n9503), 
        .S(1'b1), .Q(\U_0/U_0/U_1/LOAD_DATA [7]) );
  DFFSR \U_0/U_0/U_1/U_3/Q_int_reg[7]  ( .D(n7687), .CLK(CLK), .R(n9503), .S(
        1'b1), .Q(\U_0/U_0/U_1/RCV_DATA [7]) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[6]  ( .D(n9128), .CLK(CLK), .R(n9503), 
        .S(1'b1), .Q(\U_0/U_0/U_1/LOAD_DATA [6]) );
  DFFSR \U_0/U_0/U_1/U_3/Q_int_reg[6]  ( .D(n10575), .CLK(CLK), .R(n9503), .S(
        1'b1), .Q(\U_0/U_0/U_1/RCV_DATA [6]) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[5]  ( .D(n9127), .CLK(CLK), .R(n9503), 
        .S(1'b1), .Q(\U_0/U_0/U_1/LOAD_DATA [5]) );
  DFFSR \U_0/U_0/U_1/U_3/Q_int_reg[5]  ( .D(n7681), .CLK(CLK), .R(n9503), .S(
        1'b1), .Q(\U_0/U_0/U_1/RCV_DATA [5]) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[4]  ( .D(n9126), .CLK(CLK), .R(n9503), 
        .S(1'b1), .Q(\U_0/U_0/U_1/LOAD_DATA [4]) );
  DFFSR \U_0/U_0/U_1/U_3/Q_int_reg[4]  ( .D(n7678), .CLK(CLK), .R(n9504), .S(
        1'b1), .Q(\U_0/U_0/U_1/RCV_DATA [4]) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[3]  ( .D(n9125), .CLK(CLK), .R(n9504), 
        .S(1'b1), .Q(\U_0/U_0/U_1/LOAD_DATA [3]) );
  DFFSR \U_0/U_0/U_1/U_3/Q_int_reg[3]  ( .D(n7675), .CLK(CLK), .R(n9504), .S(
        1'b1), .Q(\U_0/U_0/U_1/RCV_DATA [3]) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[2]  ( .D(n9124), .CLK(CLK), .R(n9504), 
        .S(1'b1), .Q(\U_0/U_0/U_1/LOAD_DATA [2]) );
  DFFSR \U_0/U_0/U_1/U_3/Q_int_reg[2]  ( .D(n7672), .CLK(CLK), .R(n9504), .S(
        1'b1), .Q(\U_0/U_0/U_1/RCV_DATA [2]) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[1]  ( .D(n9123), .CLK(CLK), .R(n9504), 
        .S(1'b1), .Q(\U_0/U_0/U_1/LOAD_DATA [1]) );
  DFFSR \U_0/U_0/U_1/U_3/Q_int_reg[1]  ( .D(n7669), .CLK(CLK), .R(n9504), .S(
        1'b1), .Q(\U_0/U_0/U_1/RCV_DATA [1]) );
  DFFSR \U_0/U_0/U_1/U_6/present_val_reg[0]  ( .D(n9122), .CLK(CLK), .R(n9504), 
        .S(1'b1), .Q(\U_0/U_0/U_1/LOAD_DATA [0]) );
  DFFSR \U_0/U_0/U_1/U_3/Q_int_reg[0]  ( .D(n7666), .CLK(CLK), .R(n9504), .S(
        1'b1), .Q(\U_0/U_0/U_1/RCV_DATA [0]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/parityAccumulator_reg[0]  ( .D(n9121), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/parityAccumulator[0] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/parityAccumulator_reg[1]  ( .D(n9120), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/parityAccumulator[1] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/parityAccumulator_reg[2]  ( .D(n9119), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/parityAccumulator[2] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/parityAccumulator_reg[3]  ( .D(n9118), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/parityAccumulator[3] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/parityAccumulator_reg[4]  ( .D(n9117), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/parityAccumulator[4] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/parityAccumulator_reg[5]  ( .D(n9116), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/parityAccumulator[5] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/parityAccumulator_reg[6]  ( .D(n9115), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/parityAccumulator[6] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/parityAccumulator_reg[7]  ( .D(n9114), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/parityAccumulator[7] ) );
  DFFSR \U_0/U_0/U_1/U_8/PARITY_ERROR_reg  ( .D(
        \U_0/U_0/U_1/U_8/nextParityError ), .CLK(CLK), .R(n9504), .S(1'b1), 
        .Q(PARITY_ERROR) );
  DFFSR \U_0/U_0/U_1/U_8/parityError_reg  ( .D(
        \U_0/U_0/U_1/U_8/nextParityError ), .CLK(CLK), .R(n9504), .S(1'b1), 
        .Q(\U_0/U_0/U_1/U_8/parityError ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[0]  ( .D(n9113), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[0] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[0]  ( .D(n7662), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [0]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[1]  ( .D(n9112), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[1] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[1]  ( .D(n7661), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [1]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[2]  ( .D(n9111), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[2] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[2]  ( .D(n7660), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [2]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[3]  ( .D(n9110), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[3] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[3]  ( .D(n7659), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [3]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[4]  ( .D(n9109), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[4] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[4]  ( .D(n10344), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [4]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[5]  ( .D(n9108), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[5] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[5]  ( .D(n10345), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [5]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[6]  ( .D(n9107), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[6] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[6]  ( .D(n10346), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [6]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[7]  ( .D(n9106), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[7] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[7]  ( .D(n10347), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [7]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[8]  ( .D(n9105), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[8] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[8]  ( .D(n10348), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [8]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[9]  ( .D(n9104), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[9] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[9]  ( .D(n10349), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [9]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[10]  ( .D(n9103), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[10] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[10]  ( .D(n10350), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [10]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[11]  ( .D(n9102), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[11] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[11]  ( .D(n10351), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [11]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[12]  ( .D(n9101), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[12] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[12]  ( .D(n10352), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [12]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[13]  ( .D(n9100), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[13] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[13]  ( .D(n10353), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [13]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[14]  ( .D(n9099), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[14] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[14]  ( .D(n10354), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [14]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[15]  ( .D(n9098), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[15] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[15]  ( .D(n10355), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [15]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[16]  ( .D(n9097), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[16] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[16]  ( .D(n10356), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [16]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[17]  ( .D(n9096), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[17] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[17]  ( .D(n10357), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [17]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[18]  ( .D(n9095), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[18] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[18]  ( .D(n10358), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [18]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[19]  ( .D(n9094), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[19] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[19]  ( .D(n10359), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [19]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[20]  ( .D(n9093), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[20] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[20]  ( .D(n10360), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [20]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[21]  ( .D(n9092), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[21] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[21]  ( .D(n10361), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [21]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[22]  ( .D(n9091), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[22] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[22]  ( .D(n10362), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [22]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[23]  ( .D(n9090), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[23] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[23]  ( .D(n10363), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [23]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[24]  ( .D(n9089), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[24] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[24]  ( .D(n10364), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [24]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[25]  ( .D(n9088), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[25] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[25]  ( .D(n10365), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [25]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[26]  ( .D(n9087), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[26] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[26]  ( .D(n10366), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [26]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[27]  ( .D(n9086), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[27] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[27]  ( .D(n10367), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [27]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[28]  ( .D(n9085), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[28] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[28]  ( .D(n10368), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [28]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[29]  ( .D(n9084), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[29] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[29]  ( .D(n10369), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [29]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[30]  ( .D(n9083), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[30] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[30]  ( .D(n10370), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [30]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[31]  ( .D(n9082), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[31] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[31]  ( .D(n10371), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [31]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[32]  ( .D(n9081), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[32] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[32]  ( .D(n10372), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [32]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[33]  ( .D(n9080), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[33] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[33]  ( .D(n10373), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [33]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[34]  ( .D(n9079), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[34] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[34]  ( .D(n10374), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [34]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[35]  ( .D(n9078), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[35] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[35]  ( .D(n10375), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [35]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[36]  ( .D(n9077), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[36] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[36]  ( .D(n10376), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [36]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[37]  ( .D(n9076), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[37] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[37]  ( .D(n10377), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [37]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[38]  ( .D(n9075), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[38] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[38]  ( .D(n10378), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [38]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[39]  ( .D(n9074), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[39] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[39]  ( .D(n10379), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [39]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[40]  ( .D(n9073), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[40] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[40]  ( .D(n10380), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [40]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[41]  ( .D(n9072), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[41] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[41]  ( .D(n10381), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [41]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[42]  ( .D(n9071), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[42] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[42]  ( .D(n10382), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [42]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[43]  ( .D(n9070), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[43] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[43]  ( .D(n10383), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [43]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[44]  ( .D(n9069), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[44] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[44]  ( .D(n10384), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [44]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[45]  ( .D(n9068), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[45] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[45]  ( .D(n10385), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [45]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[46]  ( .D(n9067), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[46] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[46]  ( .D(n10386), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [46]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[47]  ( .D(n9066), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[47] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[47]  ( .D(n10387), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [47]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[48]  ( .D(n9065), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[48] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[48]  ( .D(n10388), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [48]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[49]  ( .D(n9064), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[49] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[49]  ( .D(n10389), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [49]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[50]  ( .D(n9063), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[50] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[50]  ( .D(n10390), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [50]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[51]  ( .D(n9062), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[51] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[51]  ( .D(n10391), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [51]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[52]  ( .D(n9061), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[52] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[52]  ( .D(n10392), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [52]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[53]  ( .D(n9060), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[53] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[53]  ( .D(n10393), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [53]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[54]  ( .D(n9059), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[54] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[54]  ( .D(n10394), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [54]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[55]  ( .D(n9058), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[55] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[55]  ( .D(n10395), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [55]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[56]  ( .D(n9057), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[56] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[56]  ( .D(n10396), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [56]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[57]  ( .D(n9056), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[57] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[57]  ( .D(n10397), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [57]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[58]  ( .D(n9055), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[58] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[58]  ( .D(n10398), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [58]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[59]  ( .D(n9054), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[59] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[59]  ( .D(n10399), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [59]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[60]  ( .D(n9053), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[60] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[60]  ( .D(n10400), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [60]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[61]  ( .D(n9052), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[61] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[61]  ( .D(n10401), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [61]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[62]  ( .D(n9051), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[62] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[62]  ( .D(n10402), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [62]) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/currentPlainKey_reg[63]  ( .D(n9050), .CLK(CLK), 
        .Q(\U_0/U_0/U_1/U_8/currentPlainKey[63] ) );
  DFFPOSX1 \U_0/U_0/U_1/U_8/PLAINKEY_reg[63]  ( .D(n7599), .CLK(CLK), .Q(
        \U_0/U_0/PLAINKEY [63]) );
  DFFSR \U_0/U_1/U_1/state_reg  ( .D(1'b1), .CLK(CLK), .R(n9504), .S(1'b1), 
        .Q(\U_0/U_1/U_1/state ) );
  DFFSR \U_0/U_2/U_0/DP_hold1_reg  ( .D(DPRH), .CLK(CLK), .R(1'b1), .S(n9521), 
        .Q(\U_0/U_2/U_0/DP_hold1 ) );
  DFFSR \U_0/U_2/U_0/DP_hold2_reg  ( .D(\U_0/U_2/U_0/DP_hold1 ), .CLK(CLK), 
        .R(1'b1), .S(n9521), .Q(\U_0/U_2/U_0/DP_hold2 ) );
  DFFSR \U_0/U_2/U_5/state_reg[0]  ( .D(\U_0/U_2/U_5/nextstate [0]), .CLK(CLK), 
        .R(n9505), .S(1'b1), .Q(\U_0/U_2/U_5/state[0] ) );
  DFFSR \U_0/U_2/U_5/state_reg[3]  ( .D(\U_0/U_2/U_5/nextstate [3]), .CLK(CLK), 
        .R(n9505), .S(1'b1), .Q(\U_0/U_2/U_5/state[3] ) );
  DFFSR \U_0/U_2/U_7/state_reg  ( .D(n10794), .CLK(CLK), .R(n9505), .S(1'b1), 
        .Q(\U_0/U_2/U_7/state ) );
  DFFSR \U_0/U_2/U_7/count_reg[2]  ( .D(\U_0/U_2/U_7/nextcount [2]), .CLK(CLK), 
        .R(n9505), .S(1'b1), .Q(\U_0/U_2/U_7/count[2] ) );
  DFFSR \U_0/U_2/U_7/count_reg[3]  ( .D(\U_0/U_2/U_7/nextcount [3]), .CLK(CLK), 
        .R(n9505), .S(1'b1), .Q(\U_0/U_2/U_7/count[3] ) );
  DFFSR \U_0/U_2/U_1/state_reg[0]  ( .D(\U_0/U_2/U_1/N29 ), .CLK(CLK), .R(
        n9505), .S(1'b1), .Q(\U_0/U_2/U_1/state[0] ) );
  DFFSR \U_0/U_2/U_1/DP_hold2_reg  ( .D(n9049), .CLK(CLK), .R(1'b1), .S(n9521), 
        .Q(\U_0/U_2/U_1/DP_hold2 ) );
  DFFSR \U_0/U_2/U_1/state_reg[3]  ( .D(\U_0/U_2/U_1/N32 ), .CLK(CLK), .R(
        n9505), .S(1'b1), .Q(\U_0/U_2/U_1/state[3] ) );
  DFFSR \U_0/U_2/U_1/state_reg[2]  ( .D(\U_0/U_2/U_1/N31 ), .CLK(CLK), .R(
        n9505), .S(1'b1), .Q(\U_0/U_2/U_1/state[2] ) );
  DFFSR \U_0/U_2/U_1/state_reg[1]  ( .D(n9687), .CLK(CLK), .R(n9505), .S(1'b1), 
        .Q(\U_0/U_2/U_1/state[1] ) );
  DFFSR \U_0/U_2/U_1/DP_hold1_reg  ( .D(n9048), .CLK(CLK), .R(1'b1), .S(n9521), 
        .Q(\U_0/U_2/U_1/DP_hold1 ) );
  DFFSR \U_0/U_2/U_6/present_val_reg[7]  ( .D(n9047), .CLK(CLK), .R(n9505), 
        .S(1'b1), .Q(\U_0/RCV_DATA [7]) );
  DFFSR \U_0/U_2/U_6/present_val_reg[6]  ( .D(n9046), .CLK(CLK), .R(n9505), 
        .S(1'b1), .Q(\U_0/RCV_DATA [6]) );
  DFFSR \U_0/U_2/U_6/present_val_reg[5]  ( .D(n9045), .CLK(CLK), .R(n9505), 
        .S(1'b1), .Q(\U_0/RCV_DATA [5]) );
  DFFSR \U_0/U_2/U_6/present_val_reg[4]  ( .D(n9044), .CLK(CLK), .R(n9506), 
        .S(1'b1), .Q(\U_0/RCV_DATA [4]) );
  DFFSR \U_0/U_2/U_6/present_val_reg[3]  ( .D(n9043), .CLK(CLK), .R(n9506), 
        .S(1'b1), .Q(\U_0/RCV_DATA [3]) );
  DFFSR \U_0/U_2/U_6/present_val_reg[2]  ( .D(n9042), .CLK(CLK), .R(n9506), 
        .S(1'b1), .Q(\U_0/RCV_DATA [2]) );
  DFFSR \U_0/U_2/U_6/present_val_reg[1]  ( .D(n9041), .CLK(CLK), .R(n9506), 
        .S(1'b1), .Q(\U_0/RCV_DATA [1]) );
  DFFSR \U_0/U_2/U_6/present_val_reg[0]  ( .D(n9040), .CLK(CLK), .R(n9506), 
        .S(1'b1), .Q(\U_0/RCV_DATA [0]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[7]  ( .D(n8979), .CLK(CLK), .R(
        n9506), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [7]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[15]  ( .D(n8971), .CLK(CLK), .R(
        n9506), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [15]) );
  DFFSR \U_0/U_2/U_5/state_reg[2]  ( .D(\U_0/U_2/U_5/nextstate [2]), .CLK(CLK), 
        .R(n9506), .S(1'b1), .Q(\U_0/U_2/U_5/state[2] ) );
  DFFSR \U_0/U_2/U_5/count_reg[0]  ( .D(n9033), .CLK(CLK), .R(n9506), .S(1'b1), 
        .Q(\U_0/U_2/U_5/count[0] ) );
  DFFSR \U_0/U_2/U_5/count_reg[1]  ( .D(n9034), .CLK(CLK), .R(n9506), .S(1'b1), 
        .Q(\U_0/U_2/U_5/count[1] ) );
  DFFSR \U_0/U_2/U_5/count_reg[2]  ( .D(n9035), .CLK(CLK), .R(n9506), .S(1'b1), 
        .Q(\U_0/U_2/U_5/count[2] ) );
  DFFSR \U_0/U_2/U_5/count_reg[3]  ( .D(n9036), .CLK(CLK), .R(n9507), .S(1'b1), 
        .Q(\U_0/U_2/U_5/count[3] ) );
  DFFSR \U_0/U_2/U_5/state_reg[1]  ( .D(\U_0/U_2/U_5/nextstate [1]), .CLK(CLK), 
        .R(n9507), .S(1'b1), .Q(\U_0/U_2/U_5/state[1] ) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[15]  ( .D(n9039), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[15] ) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[0]  ( .D(n9031), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[0] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[0]  ( .D(n9030), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [0]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[0]  ( .D(n9029), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [0]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[8]  ( .D(n9007), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[8] ) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[2]  ( .D(n9025), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[2] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[2]  ( .D(n9024), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [2]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[2]  ( .D(n9023), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [2]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[10]  ( .D(n9001), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[10] ) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[3]  ( .D(n9022), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[3] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[3]  ( .D(n9021), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [3]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[3]  ( .D(n9020), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [3]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[11]  ( .D(n8998), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[11] ) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[4]  ( .D(n9019), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[4] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[4]  ( .D(n9018), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [4]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[4]  ( .D(n9017), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [4]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[12]  ( .D(n8995), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[12] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[12]  ( .D(n8994), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [12]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[12]  ( .D(n8993), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [12]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[5]  ( .D(n9016), .CLK(CLK), .R(n9507), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[5] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[5]  ( .D(n9015), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [5]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[5]  ( .D(n9014), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [5]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[13]  ( .D(n8992), .CLK(CLK), .R(n9508), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[13] ) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[6]  ( .D(n9013), .CLK(CLK), .R(n9508), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[6] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[6]  ( .D(n9012), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [6]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[6]  ( .D(n9011), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [6]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[14]  ( .D(n8989), .CLK(CLK), .R(n9508), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[14] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[14]  ( .D(n8988), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [14]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[14]  ( .D(n8987), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [14]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[7]  ( .D(n9010), .CLK(CLK), .R(n9508), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[7] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[7]  ( .D(n9009), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [7]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[7]  ( .D(n9008), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [7]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[13]  ( .D(n8991), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [13]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[13]  ( .D(n8990), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [13]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[11]  ( .D(n8997), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [11]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[11]  ( .D(n8996), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [11]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[1]  ( .D(n9028), .CLK(CLK), .R(n9508), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[1] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[1]  ( .D(n9027), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [1]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[1]  ( .D(n9026), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [1]) );
  DFFSR \U_0/U_2/U_2/current_crc_reg[9]  ( .D(n9004), .CLK(CLK), .R(n9508), 
        .S(1'b1), .Q(\U_0/U_2/U_2/current_crc[9] ) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[9]  ( .D(n9003), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [9]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[9]  ( .D(n9002), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [9]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[10]  ( .D(n9000), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [10]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[10]  ( .D(n8999), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [10]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[8]  ( .D(n9006), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [8]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[8]  ( .D(n9005), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [8]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_1_reg[15]  ( .D(n9038), .CLK(CLK), .Q(
        \U_0/U_2/U_2/cache_1 [15]) );
  DFFPOSX1 \U_0/U_2/U_2/cache_2_reg[15]  ( .D(n9037), .CLK(CLK), .Q(
        \U_0/U_2/RX_CRC [15]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[0]  ( .D(n8986), .CLK(CLK), .R(
        n9508), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [0]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[8]  ( .D(n8978), .CLK(CLK), .R(
        n9508), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [8]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[1]  ( .D(n8985), .CLK(CLK), .R(
        n9508), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [1]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[9]  ( .D(n8977), .CLK(CLK), .R(
        n9508), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [9]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[2]  ( .D(n8984), .CLK(CLK), .R(
        n9508), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [2]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[10]  ( .D(n8976), .CLK(CLK), .R(
        n9508), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [10]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[3]  ( .D(n8983), .CLK(CLK), .R(
        n9509), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [3]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[11]  ( .D(n8975), .CLK(CLK), .R(
        n9509), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [11]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[4]  ( .D(n8982), .CLK(CLK), .R(
        n9509), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [4]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[12]  ( .D(n8974), .CLK(CLK), .R(
        n9509), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [12]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[5]  ( .D(n8981), .CLK(CLK), .R(
        n9509), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [5]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[13]  ( .D(n8973), .CLK(CLK), .R(
        n9509), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [13]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[6]  ( .D(n8980), .CLK(CLK), .R(
        n9509), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [6]) );
  DFFSR \U_0/U_2/U_3/present_CHECK_CRC_reg[14]  ( .D(n8972), .CLK(CLK), .R(
        n9509), .S(1'b1), .Q(\U_0/U_2/rx_CHECK_CRC [14]) );
  DFFSR \U_0/U_2/U_7/count_reg[0]  ( .D(\U_0/U_2/U_7/nextcount [0]), .CLK(CLK), 
        .R(n9509), .S(1'b1), .Q(\U_0/U_2/U_7/count[0] ) );
  DFFSR \U_0/U_2/U_7/count_reg[1]  ( .D(\U_0/U_2/U_7/nextcount [1]), .CLK(CLK), 
        .R(n9509), .S(1'b1), .Q(\U_0/U_2/U_7/count[1] ) );
  DFFPOSX1 \U_0/U_2/U_5/curR_ERROR_reg  ( .D(n9032), .CLK(CLK), .Q(
        \U_0/U_2/U_5/curR_ERROR ) );
  DFFSR \U_0/U_2/U_5/R_ERROR_reg  ( .D(n9688), .CLK(CLK), .R(n9509), .S(1'b1), 
        .Q(RE_H) );
  DFFPOSX1 \U_0/U_2/U_5/curCRC_ERROR_reg  ( .D(n8970), .CLK(CLK), .Q(
        \U_0/U_2/U_5/curCRC_ERROR ) );
  DFFPOSX1 \U_0/U_2/U_5/CRC_ERROR_reg  ( .D(n8969), .CLK(CLK), .Q(CRCE_H) );
  DFFSR \U_0/U_3/U_0/dp_tx_out_reg  ( .D(\U_0/U_3/U_0/DE_holdout_nxt ), .CLK(
        CLK), .R(1'b1), .S(n9521), .Q(DPTS) );
  DFFSR \U_0/U_3/U_0/state_reg[3]  ( .D(\U_0/U_3/U_0/nextstate [3]), .CLK(CLK), 
        .R(n9509), .S(1'b1), .Q(\U_0/U_3/U_0/state[3] ) );
  DFFSR \U_0/U_3/U_0/DE_holdout_reg  ( .D(\U_0/U_3/U_0/DE_holdout_nxt ), .CLK(
        CLK), .R(1'b1), .S(n9521), .Q(\U_0/U_3/U_0/DE_holdout ) );
  DFFPOSX1 \U_0/U_3/U_0/DE_holdout_last_reg  ( .D(n7532), .CLK(CLK), .Q(
        \U_0/U_3/U_0/DE_holdout_last ) );
  DFFSR \U_0/U_3/U_4/SHIFT_ENABLE_E_reg  ( .D(n7754), .CLK(CLK), .R(n9510), 
        .S(1'b1), .Q(\U_0/U_3/SHIFT_ENABLE_E ) );
  DFFSR \U_0/U_3/U_0/state_reg[2]  ( .D(\U_0/U_3/U_0/nextstate [2]), .CLK(CLK), 
        .R(n9510), .S(1'b1), .Q(\U_0/U_3/U_0/state[2] ) );
  DFFSR \U_0/U_3/U_0/state_reg[0]  ( .D(\U_0/U_3/U_0/nextstate [0]), .CLK(CLK), 
        .R(n9510), .S(1'b1), .Q(\U_0/U_3/U_0/state[0] ) );
  DFFSR \U_0/U_3/U_0/state_reg[1]  ( .D(\U_0/U_3/U_0/nextstate [1]), .CLK(CLK), 
        .R(n9510), .S(1'b1), .Q(\U_0/U_3/U_0/state[1] ) );
  DFFSR \U_0/U_3/U_3/count_reg[6]  ( .D(n8495), .CLK(CLK), .R(n9510), .S(1'b1), 
        .Q(\U_0/U_3/U_3/N188 ) );
  DFFSR \U_0/U_3/U_3/state_reg[1]  ( .D(\U_0/U_3/U_3/nextstate [1]), .CLK(CLK), 
        .R(n9510), .S(1'b1), .Q(\U_0/U_3/U_3/state[1] ) );
  DFFSR \U_0/U_3/U_3/state_reg[2]  ( .D(\U_0/U_3/U_3/nextstate [2]), .CLK(CLK), 
        .R(n9510), .S(1'b1), .Q(\U_0/U_3/U_3/state[2] ) );
  DFFSR \U_0/U_3/U_3/state_reg[0]  ( .D(\U_0/U_3/U_3/nextstate [0]), .CLK(CLK), 
        .R(n9510), .S(1'b1), .Q(\U_0/U_3/U_3/state[0] ) );
  DFFSR \U_0/U_1/U_0/state_reg[2]  ( .D(\U_0/U_1/U_0/nextState [2]), .CLK(CLK), 
        .R(n9510), .S(1'b1), .Q(\U_0/U_1/U_0/state[2] ) );
  DFFPOSX1 \U_0/U_1/U_0/R_ENABLE_reg  ( .D(n7522), .CLK(CLK), .Q(
        \U_0/U_1/R_ENABLE ) );
  DFFSR \U_0/U_1/U_1/readptr_reg[0]  ( .D(\U_0/U_1/U_1/N343 ), .CLK(CLK), .R(
        n9510), .S(1'b1), .Q(\U_0/U_1/U_1/readptr[0] ) );
  DFFSR \U_0/U_1/U_1/readptr_reg[1]  ( .D(\U_0/U_1/U_1/N344 ), .CLK(CLK), .R(
        n9510), .S(1'b1), .Q(\U_0/U_1/U_1/readptr[1] ) );
  DFFSR \U_0/U_1/U_1/readptr_reg[2]  ( .D(\U_0/U_1/U_1/N345 ), .CLK(CLK), .R(
        n9510), .S(1'b1), .Q(\U_0/U_1/U_1/readptr[2] ) );
  DFFSR \U_0/U_1/U_1/readptr_reg[3]  ( .D(\U_0/U_1/U_1/N346 ), .CLK(CLK), .R(
        n9511), .S(1'b1), .Q(\U_0/U_1/U_1/readptr[3] ) );
  DFFSR \U_0/U_1/U_1/readptr_reg[4]  ( .D(\U_0/U_1/U_1/N347 ), .CLK(CLK), .R(
        n9511), .S(1'b1), .Q(\U_0/U_1/U_1/readptr[4] ) );
  DFFSR \U_0/U_1/U_1/writeptr_reg[4]  ( .D(n8967), .CLK(CLK), .R(n9511), .S(
        1'b1), .Q(\U_0/U_1/U_1/writeptr[4] ) );
  DFFSR \U_0/U_1/U_1/writeptr_reg[3]  ( .D(n8963), .CLK(CLK), .R(n9511), .S(
        1'b1), .Q(\U_0/U_1/U_1/writeptr[3] ) );
  DFFSR \U_0/U_1/U_1/writeptr_reg[0]  ( .D(n8966), .CLK(CLK), .R(n9511), .S(
        1'b1), .Q(\U_0/U_1/U_1/writeptr[0] ) );
  DFFSR \U_0/U_1/U_1/writeptr_reg[1]  ( .D(n8965), .CLK(CLK), .R(n9511), .S(
        1'b1), .Q(\U_0/U_1/U_1/writeptr[1] ) );
  DFFSR \U_0/U_1/U_1/writeptr_reg[2]  ( .D(n8964), .CLK(CLK), .R(n9511), .S(
        1'b1), .Q(\U_0/U_1/U_1/writeptr[2] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[0][0]  ( .D(n9741), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[0][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[0][1]  ( .D(n9740), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[0][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[0][0]  ( .D(n9948), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[0][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[0][1]  ( .D(n9947), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[0][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[0][2]  ( .D(n9946), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[0][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[0][3]  ( .D(n9945), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[0][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[0][4]  ( .D(n9944), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[0][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[0][5]  ( .D(n9943), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[0][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[0][6]  ( .D(n9942), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[0][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[0][7]  ( .D(n9941), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[0][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[1][0]  ( .D(n9738), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[1][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[1][1]  ( .D(n9737), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[1][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[1][0]  ( .D(n9939), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[1][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[1][1]  ( .D(n9938), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[1][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[1][2]  ( .D(n9937), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[1][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[1][3]  ( .D(n9936), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[1][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[1][4]  ( .D(n9935), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[1][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[1][5]  ( .D(n9934), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[1][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[1][6]  ( .D(n9933), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[1][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[1][7]  ( .D(n9932), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[1][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[2][0]  ( .D(n9735), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[2][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[2][1]  ( .D(n9734), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[2][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[2][0]  ( .D(n9930), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[2][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[2][1]  ( .D(n9929), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[2][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[2][2]  ( .D(n9928), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[2][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[2][3]  ( .D(n9927), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[2][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[2][4]  ( .D(n9926), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[2][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[2][5]  ( .D(n9925), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[2][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[2][6]  ( .D(n9924), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[2][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[2][7]  ( .D(n9923), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[2][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[3][0]  ( .D(n9732), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[3][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[3][1]  ( .D(n9731), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[3][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[3][0]  ( .D(n9921), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[3][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[3][1]  ( .D(n9920), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[3][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[3][2]  ( .D(n9919), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[3][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[3][3]  ( .D(n9918), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[3][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[3][4]  ( .D(n9917), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[3][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[3][5]  ( .D(n9916), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[3][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[3][6]  ( .D(n9915), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[3][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[3][7]  ( .D(n9914), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[3][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[4][0]  ( .D(n8908), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[4][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[4][1]  ( .D(n8907), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[4][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[4][0]  ( .D(n8682), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[4][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[4][1]  ( .D(n8681), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[4][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[4][2]  ( .D(n8680), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[4][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[4][3]  ( .D(n8679), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[4][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[4][4]  ( .D(n8678), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[4][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[4][5]  ( .D(n8677), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[4][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[4][6]  ( .D(n8676), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[4][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[4][7]  ( .D(n8675), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[4][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[5][0]  ( .D(n8910), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[5][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[5][1]  ( .D(n8909), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[5][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[5][0]  ( .D(n8690), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[5][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[5][1]  ( .D(n8689), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[5][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[5][2]  ( .D(n8688), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[5][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[5][3]  ( .D(n8687), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[5][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[5][4]  ( .D(n8686), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[5][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[5][5]  ( .D(n8685), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[5][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[5][6]  ( .D(n8684), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[5][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[5][7]  ( .D(n8683), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[5][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[6][0]  ( .D(n8698), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[6][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[6][1]  ( .D(n8697), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[6][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[6][2]  ( .D(n8696), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[6][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[6][3]  ( .D(n8695), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[6][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[6][4]  ( .D(n8694), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[6][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[6][5]  ( .D(n8693), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[6][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[6][6]  ( .D(n8692), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[6][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[6][7]  ( .D(n8691), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[6][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[7][6]  ( .D(n8706), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[7][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[7][7]  ( .D(n8705), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[7][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[7][0]  ( .D(n8704), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[7][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[7][1]  ( .D(n8703), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[7][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[7][2]  ( .D(n8702), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[7][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[7][3]  ( .D(n8701), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[7][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[7][4]  ( .D(n8700), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[7][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[7][5]  ( .D(n8699), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[7][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[11][1]  ( .D(n8922), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[11][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[11][0]  ( .D(n8921), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[11][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[6][0]  ( .D(n8912), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[6][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[6][1]  ( .D(n8911), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[6][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[7][0]  ( .D(n8914), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[7][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[7][1]  ( .D(n8913), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[7][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[11][0]  ( .D(n8738), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[11][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[11][1]  ( .D(n8737), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[11][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[11][2]  ( .D(n8736), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[11][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[11][3]  ( .D(n8735), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[11][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[11][4]  ( .D(n8734), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[11][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[11][5]  ( .D(n8733), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[11][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[11][6]  ( .D(n8732), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[11][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[11][7]  ( .D(n8731), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[11][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[8][0]  ( .D(n8916), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[8][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[8][1]  ( .D(n8915), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[8][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[8][0]  ( .D(n8714), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[8][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[8][1]  ( .D(n8713), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[8][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[8][2]  ( .D(n8712), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[8][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[8][3]  ( .D(n8711), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[8][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[8][4]  ( .D(n8710), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[8][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[8][5]  ( .D(n8709), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[8][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[8][6]  ( .D(n8708), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[8][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[8][7]  ( .D(n8707), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[8][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[9][0]  ( .D(n8918), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[9][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[9][1]  ( .D(n8917), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[9][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[9][0]  ( .D(n8722), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[9][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[9][1]  ( .D(n8721), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[9][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[9][2]  ( .D(n8720), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[9][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[9][3]  ( .D(n8719), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[9][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[9][4]  ( .D(n8718), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[9][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[9][5]  ( .D(n8717), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[9][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[9][6]  ( .D(n8716), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[9][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[9][7]  ( .D(n8715), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[9][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[10][0]  ( .D(n8920), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[10][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[10][1]  ( .D(n8919), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[10][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[10][0]  ( .D(n8730), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[10][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[10][1]  ( .D(n8729), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[10][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[10][2]  ( .D(n8728), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[10][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[10][3]  ( .D(n8727), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[10][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[10][4]  ( .D(n8726), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[10][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[10][5]  ( .D(n8725), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[10][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[10][6]  ( .D(n8724), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[10][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[10][7]  ( .D(n8723), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[10][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[12][0]  ( .D(n9783), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[12][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[12][1]  ( .D(n9782), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[12][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[12][0]  ( .D(n9904), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[12][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[12][1]  ( .D(n9903), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[12][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[12][2]  ( .D(n9902), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[12][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[12][3]  ( .D(n9901), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[12][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[12][4]  ( .D(n9900), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[12][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[12][5]  ( .D(n9899), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[12][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[12][6]  ( .D(n9898), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[12][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[12][7]  ( .D(n9897), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[12][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[13][0]  ( .D(n9780), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[13][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[13][1]  ( .D(n9779), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[13][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[13][0]  ( .D(n9895), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[13][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[13][1]  ( .D(n9894), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[13][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[13][2]  ( .D(n9893), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[13][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[13][3]  ( .D(n9892), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[13][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[13][4]  ( .D(n9891), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[13][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[13][5]  ( .D(n9890), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[13][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[13][6]  ( .D(n9889), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[13][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[13][7]  ( .D(n9888), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[13][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[14][0]  ( .D(n9886), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[14][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[14][1]  ( .D(n9885), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[14][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[14][2]  ( .D(n9884), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[14][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[14][3]  ( .D(n9883), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[14][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[14][4]  ( .D(n9882), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[14][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[14][5]  ( .D(n9881), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[14][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[14][6]  ( .D(n9880), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[14][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[14][7]  ( .D(n9879), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[14][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[15][0]  ( .D(n9877), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[15][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[15][1]  ( .D(n9876), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[15][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[15][2]  ( .D(n9875), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[15][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[15][3]  ( .D(n9874), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[15][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[15][4]  ( .D(n9873), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[15][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[15][5]  ( .D(n9872), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[15][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[15][6]  ( .D(n9871), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[15][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[15][7]  ( .D(n9870), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[15][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[24][0]  ( .D(n9755), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[24][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[24][1]  ( .D(n9754), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[24][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[24][0]  ( .D(n9828), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[24][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[24][1]  ( .D(n9827), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[24][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[24][2]  ( .D(n9826), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[24][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[24][3]  ( .D(n9825), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[24][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[24][4]  ( .D(n9824), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[24][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[24][5]  ( .D(n9823), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[24][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[24][6]  ( .D(n9822), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[24][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[24][7]  ( .D(n9821), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[24][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[25][0]  ( .D(n9752), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[25][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[25][1]  ( .D(n9751), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[25][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[25][0]  ( .D(n9819), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[25][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[25][1]  ( .D(n9818), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[25][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[25][2]  ( .D(n9817), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[25][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[25][3]  ( .D(n9816), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[25][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[25][4]  ( .D(n9815), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[25][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[25][5]  ( .D(n9814), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[25][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[25][6]  ( .D(n9813), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[25][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[25][7]  ( .D(n9812), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[25][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[26][0]  ( .D(n9749), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[26][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[26][1]  ( .D(n9748), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[26][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[26][0]  ( .D(n9810), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[26][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[26][1]  ( .D(n9809), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[26][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[26][2]  ( .D(n9808), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[26][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[26][3]  ( .D(n9807), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[26][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[26][4]  ( .D(n9806), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[26][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[26][5]  ( .D(n9805), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[26][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[26][6]  ( .D(n9804), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[26][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[26][7]  ( .D(n9803), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[26][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[27][0]  ( .D(n9746), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[27][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[27][1]  ( .D(n9745), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[27][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[27][0]  ( .D(n9801), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[27][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[27][1]  ( .D(n9800), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[27][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[27][2]  ( .D(n9799), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[27][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[27][3]  ( .D(n9798), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[27][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[27][4]  ( .D(n9797), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[27][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[27][5]  ( .D(n9796), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[27][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[27][6]  ( .D(n9795), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[27][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[27][7]  ( .D(n9794), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[27][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[28][0]  ( .D(n8956), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[28][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[28][1]  ( .D(n8955), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[28][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[28][0]  ( .D(n8874), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[28][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[28][1]  ( .D(n8873), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[28][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[28][2]  ( .D(n8872), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[28][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[28][3]  ( .D(n8871), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[28][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[28][4]  ( .D(n8870), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[28][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[28][5]  ( .D(n8869), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[28][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[28][6]  ( .D(n8868), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[28][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[28][7]  ( .D(n8867), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[28][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[29][0]  ( .D(n8958), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[29][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[29][1]  ( .D(n8957), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[29][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[29][0]  ( .D(n8882), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[29][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[29][1]  ( .D(n8881), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[29][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[29][2]  ( .D(n8880), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[29][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[29][3]  ( .D(n8879), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[29][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[29][4]  ( .D(n8878), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[29][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[29][5]  ( .D(n8877), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[29][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[29][6]  ( .D(n8876), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[29][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[29][7]  ( .D(n8875), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[29][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[30][0]  ( .D(n8960), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[30][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[30][1]  ( .D(n8959), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[30][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[30][0]  ( .D(n8890), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[30][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[30][1]  ( .D(n8889), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[30][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[30][2]  ( .D(n8888), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[30][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[30][3]  ( .D(n8887), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[30][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[30][4]  ( .D(n8886), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[30][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[30][5]  ( .D(n8885), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[30][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[30][6]  ( .D(n8884), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[30][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[30][7]  ( .D(n8883), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[30][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[31][0]  ( .D(n8962), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[31][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[31][1]  ( .D(n8961), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[31][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[31][0]  ( .D(n8898), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[31][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[31][1]  ( .D(n8897), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[31][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[31][2]  ( .D(n8896), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[31][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[31][3]  ( .D(n8895), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[31][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[31][4]  ( .D(n8894), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[31][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[31][5]  ( .D(n8893), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[31][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[31][6]  ( .D(n8892), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[31][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[31][7]  ( .D(n8891), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[31][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[14][0]  ( .D(n9777), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[14][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[14][1]  ( .D(n9776), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[14][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[15][0]  ( .D(n9774), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[15][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[15][1]  ( .D(n9773), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[15][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[16][0]  ( .D(n8932), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[16][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[16][1]  ( .D(n8931), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[16][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[16][0]  ( .D(n8778), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[16][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[16][1]  ( .D(n8777), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[16][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[16][2]  ( .D(n8776), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[16][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[16][3]  ( .D(n8775), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[16][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[16][4]  ( .D(n8774), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[16][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[16][5]  ( .D(n8773), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[16][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[16][6]  ( .D(n8772), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[16][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[16][7]  ( .D(n8771), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[16][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[17][0]  ( .D(n8934), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[17][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[17][1]  ( .D(n8933), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[17][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[17][0]  ( .D(n8786), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[17][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[17][1]  ( .D(n8785), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[17][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[17][2]  ( .D(n8784), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[17][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[17][3]  ( .D(n8783), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[17][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[17][4]  ( .D(n8782), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[17][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[17][5]  ( .D(n8781), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[17][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[17][6]  ( .D(n8780), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[17][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[17][7]  ( .D(n8779), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[17][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[18][0]  ( .D(n8936), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[18][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[18][1]  ( .D(n8935), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[18][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[18][0]  ( .D(n8794), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[18][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[18][1]  ( .D(n8793), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[18][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[18][2]  ( .D(n8792), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[18][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[18][3]  ( .D(n8791), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[18][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[18][4]  ( .D(n8790), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[18][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[18][5]  ( .D(n8789), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[18][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[18][6]  ( .D(n8788), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[18][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[18][7]  ( .D(n8787), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[18][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[19][0]  ( .D(n8938), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[19][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[19][1]  ( .D(n8937), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[19][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[19][3]  ( .D(n8802), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[19][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[19][4]  ( .D(n8801), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[19][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[19][5]  ( .D(n8800), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[19][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[19][6]  ( .D(n8799), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[19][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[19][7]  ( .D(n8798), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[19][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[19][0]  ( .D(n8797), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[19][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[19][1]  ( .D(n8796), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[19][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[19][2]  ( .D(n8795), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[19][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[20][0]  ( .D(n9767), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[20][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[20][1]  ( .D(n9766), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[20][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[20][0]  ( .D(n9864), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[20][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[20][1]  ( .D(n9863), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[20][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[20][2]  ( .D(n9862), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[20][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[20][3]  ( .D(n9861), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[20][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[20][4]  ( .D(n9860), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[20][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[20][5]  ( .D(n9859), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[20][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[20][6]  ( .D(n9858), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[20][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[20][7]  ( .D(n9857), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[20][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[21][0]  ( .D(n9764), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[21][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[21][1]  ( .D(n9763), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[21][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[21][0]  ( .D(n9855), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[21][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[21][1]  ( .D(n9854), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[21][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[21][2]  ( .D(n9853), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[21][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[21][3]  ( .D(n9852), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[21][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[21][4]  ( .D(n9851), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[21][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[21][5]  ( .D(n9850), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[21][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[21][6]  ( .D(n9849), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[21][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[21][7]  ( .D(n9848), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[21][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[22][0]  ( .D(n9761), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[22][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[22][1]  ( .D(n9760), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[22][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[22][0]  ( .D(n9846), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[22][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[22][1]  ( .D(n9845), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[22][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[22][2]  ( .D(n9844), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[22][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[22][3]  ( .D(n9843), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[22][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[22][4]  ( .D(n9842), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[22][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[22][5]  ( .D(n9841), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[22][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[22][6]  ( .D(n9840), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[22][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[22][7]  ( .D(n9839), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[22][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[23][0]  ( .D(n9758), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[23][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/opcode_reg[23][1]  ( .D(n9757), .CLK(CLK), .Q(
        \U_0/U_1/U_1/opcode[23][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[23][0]  ( .D(n9837), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[23][0] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[23][1]  ( .D(n9836), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[23][1] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[23][2]  ( .D(n9835), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[23][2] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[23][3]  ( .D(n9834), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[23][3] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[23][4]  ( .D(n9833), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[23][4] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[23][5]  ( .D(n9832), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[23][5] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[23][6]  ( .D(n9831), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[23][6] ) );
  DFFPOSX1 \U_0/U_1/U_1/memory_reg[23][7]  ( .D(n9830), .CLK(CLK), .Q(
        \U_0/U_1/U_1/memory[23][7] ) );
  DFFPOSX1 \U_0/U_1/U_1/FULL_reg  ( .D(n10403), .CLK(CLK), .Q(FULL_H) );
  DFFPOSX1 \U_0/U_1/U_1/EMPTY_reg  ( .D(n10404), .CLK(CLK), .Q(EMPTY_H) );
  DFFSR \U_0/U_1/U_1/BYTE_COUNT_reg[0]  ( .D(\U_0/U_1/U_1/N338 ), .CLK(CLK), 
        .R(n9511), .S(1'b1), .Q(\U_0/U_1/BYTE_COUNT [0]) );
  DFFSR \U_0/U_1/U_1/BYTE_COUNT_reg[1]  ( .D(\U_0/U_1/U_1/N339 ), .CLK(CLK), 
        .R(n9511), .S(1'b1), .Q(\U_0/U_1/BYTE_COUNT [1]) );
  DFFSR \U_0/U_1/U_1/BYTE_COUNT_reg[2]  ( .D(\U_0/U_1/U_1/N340 ), .CLK(CLK), 
        .R(n9511), .S(1'b1), .Q(\U_0/U_1/BYTE_COUNT [2]) );
  DFFSR \U_0/U_1/U_1/BYTE_COUNT_reg[3]  ( .D(\U_0/U_1/U_1/N341 ), .CLK(CLK), 
        .R(n9511), .S(1'b1), .Q(\U_0/U_1/BYTE_COUNT [3]) );
  DFFSR \U_0/U_1/U_1/BYTE_COUNT_reg[4]  ( .D(\U_0/U_1/U_1/N342 ), .CLK(CLK), 
        .R(n9511), .S(1'b1), .Q(\U_0/U_1/U_0/N39 ) );
  DFFPOSX1 \U_0/U_1/U_1/DATA_reg[0]  ( .D(n8642), .CLK(CLK), .Q(
        \U_0/U_1/DATA [0]) );
  DFFPOSX1 \U_0/U_1/U_1/DATA_reg[1]  ( .D(n8641), .CLK(CLK), .Q(
        \U_0/U_1/DATA [1]) );
  DFFPOSX1 \U_0/U_1/U_1/DATA_reg[2]  ( .D(n8640), .CLK(CLK), .Q(
        \U_0/U_1/DATA [2]) );
  DFFPOSX1 \U_0/U_1/U_1/DATA_reg[3]  ( .D(n8639), .CLK(CLK), .Q(
        \U_0/U_1/DATA [3]) );
  DFFPOSX1 \U_0/U_1/U_1/DATA_reg[4]  ( .D(n8638), .CLK(CLK), .Q(
        \U_0/U_1/DATA [4]) );
  DFFPOSX1 \U_0/U_1/U_1/DATA_reg[5]  ( .D(n8637), .CLK(CLK), .Q(
        \U_0/U_1/DATA [5]) );
  DFFPOSX1 \U_0/U_1/U_1/DATA_reg[6]  ( .D(n8636), .CLK(CLK), .Q(
        \U_0/U_1/DATA [6]) );
  DFFPOSX1 \U_0/U_1/U_1/DATA_reg[7]  ( .D(n8635), .CLK(CLK), .Q(
        \U_0/U_1/DATA [7]) );
  DFFPOSX1 \U_0/U_1/U_1/OUT_OPCODE_reg[0]  ( .D(n8634), .CLK(CLK), .Q(
        \U_0/U_1/OUT_OPCODE [0]) );
  DFFPOSX1 \U_0/U_1/U_1/OUT_OPCODE_reg[1]  ( .D(n8633), .CLK(CLK), .Q(
        \U_0/U_1/OUT_OPCODE [1]) );
  DFFSR \U_0/U_1/U_0/state_reg[0]  ( .D(\U_0/U_1/U_0/nextState [0]), .CLK(CLK), 
        .R(n9512), .S(1'b1), .Q(\U_0/U_1/U_0/state[0] ) );
  DFFSR \U_0/U_1/U_0/state_reg[1]  ( .D(\U_0/U_1/U_0/nextState [1]), .CLK(CLK), 
        .R(n9512), .S(1'b1), .Q(\U_0/U_1/U_0/state[1] ) );
  DFFPOSX1 \U_0/U_1/U_0/B_READY_reg  ( .D(n7502), .CLK(CLK), .Q(\U_0/B_READY )
         );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_OPCODE_reg[0]  ( .D(n7501), .CLK(CLK), .Q(
        \U_0/PRGA_OPCODE[0] ) );
  DFFPOSX1 \U_0/U_1/U_0/tempOpcode_reg[0]  ( .D(n7500), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempOpcode [0]) );
  DFFPOSX1 \U_0/U_1/U_0/tempData_reg[7]  ( .D(n7499), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempData [7]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_IN_reg[7]  ( .D(n7498), .CLK(CLK), .Q(
        \U_0/PRGA_IN [7]) );
  DFFPOSX1 \U_0/U_1/U_0/tempData_reg[6]  ( .D(n7497), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempData [6]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_IN_reg[6]  ( .D(n7496), .CLK(CLK), .Q(
        \U_0/PRGA_IN [6]) );
  DFFPOSX1 \U_0/U_1/U_0/tempData_reg[5]  ( .D(n7495), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempData [5]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_IN_reg[5]  ( .D(n7494), .CLK(CLK), .Q(
        \U_0/PRGA_IN [5]) );
  DFFPOSX1 \U_0/U_1/U_0/tempData_reg[4]  ( .D(n7493), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempData [4]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_IN_reg[4]  ( .D(n7492), .CLK(CLK), .Q(
        \U_0/PRGA_IN [4]) );
  DFFPOSX1 \U_0/U_1/U_0/tempData_reg[3]  ( .D(n7491), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempData [3]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_IN_reg[3]  ( .D(n7490), .CLK(CLK), .Q(
        \U_0/PRGA_IN [3]) );
  DFFPOSX1 \U_0/U_1/U_0/tempData_reg[2]  ( .D(n7489), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempData [2]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_IN_reg[2]  ( .D(n7488), .CLK(CLK), .Q(
        \U_0/PRGA_IN [2]) );
  DFFPOSX1 \U_0/U_1/U_0/tempData_reg[1]  ( .D(n7487), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempData [1]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_IN_reg[1]  ( .D(n7486), .CLK(CLK), .Q(
        \U_0/PRGA_IN [1]) );
  DFFPOSX1 \U_0/U_1/U_0/tempData_reg[0]  ( .D(n7485), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempData [0]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_IN_reg[0]  ( .D(n7484), .CLK(CLK), .Q(
        \U_0/PRGA_IN [0]) );
  DFFPOSX1 \U_0/U_1/U_0/PRGA_OPCODE_reg[1]  ( .D(n7483), .CLK(CLK), .Q(
        \U_0/PRGA_OPCODE[1] ) );
  DFFSR \U_0/U_3/U_3/count_reg[0]  ( .D(n8968), .CLK(CLK), .R(n9512), .S(1'b1), 
        .Q(\U_0/U_3/U_3/count[0] ) );
  DFFSR \U_0/U_3/U_3/count_reg[5]  ( .D(n8496), .CLK(CLK), .R(n9512), .S(1'b1), 
        .Q(\U_0/U_3/U_3/count[5] ) );
  DFFSR \U_0/U_3/U_3/count_reg[1]  ( .D(n8500), .CLK(CLK), .R(n9512), .S(1'b1), 
        .Q(\U_0/U_3/U_3/count[1] ) );
  DFFSR \U_0/U_3/U_3/count_reg[2]  ( .D(n8499), .CLK(CLK), .R(n9512), .S(1'b1), 
        .Q(\U_0/U_3/U_3/count[2] ) );
  DFFSR \U_0/U_3/U_3/count_reg[3]  ( .D(n8498), .CLK(CLK), .R(n9512), .S(1'b1), 
        .Q(\U_0/U_3/U_3/count[3] ) );
  DFFSR \U_0/U_3/U_3/count_reg[4]  ( .D(n8497), .CLK(CLK), .R(n9512), .S(1'b1), 
        .Q(\U_0/U_3/U_3/count[4] ) );
  DFFSR \U_0/U_0/U_0/state_reg[0]  ( .D(\U_0/U_0/U_0/nextState [0]), .CLK(CLK), 
        .R(n9512), .S(1'b1), .Q(\U_0/U_0/U_0/state[0] ) );
  DFFPOSX1 \U_0/U_0/U_0/permuteComplete_reg  ( .D(n8509), .CLK(CLK), .Q(
        \U_0/U_0/U_0/permuteComplete ) );
  DFFSR \U_0/U_0/U_0/state_reg[3]  ( .D(\U_0/U_0/U_0/nextState [3]), .CLK(CLK), 
        .R(n9512), .S(1'b1), .Q(\U_0/U_0/U_0/state[3] ) );
  DFFSR \U_0/U_0/U_0/state_reg[4]  ( .D(\U_0/U_0/U_0/nextState [4]), .CLK(CLK), 
        .R(n9512), .S(1'b1), .Q(\U_0/U_0/U_0/state[4] ) );
  DFFPOSX1 \U_0/U_0/U_0/prefillCounter_reg[7]  ( .D(n8501), .CLK(CLK), .Q(
        \U_0/U_0/U_0/prefillCounter[7] ) );
  DFFSR \U_0/U_0/U_0/state_reg[1]  ( .D(\U_0/U_0/U_0/nextState [1]), .CLK(CLK), 
        .R(n9512), .S(1'b1), .Q(\U_0/U_0/U_0/state[1] ) );
  DFFSR \U_0/U_0/U_0/state_reg[2]  ( .D(\U_0/U_0/U_0/nextState [2]), .CLK(CLK), 
        .R(n9518), .S(1'b1), .Q(\U_0/U_0/U_0/state[2] ) );
  DFFPOSX1 \U_0/U_0/U_0/prefillCounter_reg[0]  ( .D(n8508), .CLK(CLK), .Q(
        \U_0/U_0/U_0/prefillCounter[0] ) );
  DFFPOSX1 \U_0/U_0/U_0/prefillCounter_reg[1]  ( .D(n8507), .CLK(CLK), .Q(
        \U_0/U_0/U_0/prefillCounter[1] ) );
  DFFPOSX1 \U_0/U_0/U_0/prefillCounter_reg[2]  ( .D(n8506), .CLK(CLK), .Q(
        \U_0/U_0/U_0/prefillCounter[2] ) );
  DFFPOSX1 \U_0/U_0/U_0/prefillCounter_reg[3]  ( .D(n8505), .CLK(CLK), .Q(
        \U_0/U_0/U_0/prefillCounter[3] ) );
  DFFPOSX1 \U_0/U_0/U_0/prefillCounter_reg[4]  ( .D(n8504), .CLK(CLK), .Q(
        \U_0/U_0/U_0/prefillCounter[4] ) );
  DFFPOSX1 \U_0/U_0/U_0/prefillCounter_reg[5]  ( .D(n8503), .CLK(CLK), .Q(
        \U_0/U_0/U_0/prefillCounter[5] ) );
  DFFPOSX1 \U_0/U_0/U_0/prefillCounter_reg[6]  ( .D(n8502), .CLK(CLK), .Q(
        \U_0/U_0/U_0/prefillCounter[6] ) );
  DFFSR \U_0/U_0/U_0/PDATA_READY_reg  ( .D(n11145), .CLK(CLK), .R(n9519), .S(
        1'b1), .Q(\U_0/PDATA_READY ) );
  DFFPOSX1 \U_0/U_0/U_0/intj_reg[7]  ( .D(n8537), .CLK(CLK), .Q(
        \U_0/U_0/U_0/intj[7] ) );
  DFFPOSX1 \U_0/U_0/U_0/intj_reg[0]  ( .D(n8544), .CLK(CLK), .Q(
        \U_0/U_0/U_0/intj[0] ) );
  DFFPOSX1 \U_0/U_0/U_0/intj_reg[1]  ( .D(n8543), .CLK(CLK), .Q(
        \U_0/U_0/U_0/intj[1] ) );
  DFFPOSX1 \U_0/U_0/U_0/intj_reg[2]  ( .D(n8542), .CLK(CLK), .Q(
        \U_0/U_0/U_0/intj[2] ) );
  DFFPOSX1 \U_0/U_0/U_0/intj_reg[3]  ( .D(n8541), .CLK(CLK), .Q(
        \U_0/U_0/U_0/intj[3] ) );
  DFFPOSX1 \U_0/U_0/U_0/intj_reg[4]  ( .D(n8540), .CLK(CLK), .Q(
        \U_0/U_0/U_0/intj[4] ) );
  DFFPOSX1 \U_0/U_0/U_0/intj_reg[5]  ( .D(n8539), .CLK(CLK), .Q(
        \U_0/U_0/U_0/intj[5] ) );
  DFFPOSX1 \U_0/U_0/U_0/intj_reg[6]  ( .D(n8538), .CLK(CLK), .Q(
        \U_0/U_0/U_0/intj[6] ) );
  DFFPOSX1 \U_0/U_0/U_0/inti_reg[0]  ( .D(n10013), .CLK(CLK), .Q(
        \U_0/U_0/U_0/inti[0] ) );
  DFFPOSX1 \U_0/U_0/U_0/inti_reg[1]  ( .D(n10014), .CLK(CLK), .Q(
        \U_0/U_0/U_0/inti[1] ) );
  DFFPOSX1 \U_0/U_0/U_0/inti_reg[2]  ( .D(n10015), .CLK(CLK), .Q(
        \U_0/U_0/U_0/inti[2] ) );
  DFFPOSX1 \U_0/U_0/U_0/inti_reg[3]  ( .D(n10016), .CLK(CLK), .Q(
        \U_0/U_0/U_0/inti[3] ) );
  DFFPOSX1 \U_0/U_0/U_0/inti_reg[4]  ( .D(n10017), .CLK(CLK), .Q(
        \U_0/U_0/U_0/inti[4] ) );
  DFFPOSX1 \U_0/U_0/U_0/inti_reg[5]  ( .D(n10018), .CLK(CLK), .Q(
        \U_0/U_0/U_0/inti[5] ) );
  DFFPOSX1 \U_0/U_0/U_0/inti_reg[6]  ( .D(n10019), .CLK(CLK), .Q(
        \U_0/U_0/U_0/inti[6] ) );
  DFFPOSX1 \U_0/U_0/U_0/inti_reg[7]  ( .D(n10020), .CLK(CLK), .Q(
        \U_0/U_0/U_0/inti[7] ) );
  DFFPOSX1 \U_0/U_0/U_0/extratemp_reg[7]  ( .D(n10039), .CLK(CLK), .Q(
        \U_0/U_0/U_0/extratemp[7] ) );
  DFFPOSX1 \U_0/U_0/U_0/extratemp_reg[6]  ( .D(n10038), .CLK(CLK), .Q(
        \U_0/U_0/U_0/extratemp[6] ) );
  DFFPOSX1 \U_0/U_0/U_0/extratemp_reg[5]  ( .D(n10037), .CLK(CLK), .Q(
        \U_0/U_0/U_0/extratemp[5] ) );
  DFFPOSX1 \U_0/U_0/U_0/extratemp_reg[4]  ( .D(n10036), .CLK(CLK), .Q(
        \U_0/U_0/U_0/extratemp[4] ) );
  DFFPOSX1 \U_0/U_0/U_0/extratemp_reg[3]  ( .D(n10035), .CLK(CLK), .Q(
        \U_0/U_0/U_0/extratemp[3] ) );
  DFFPOSX1 \U_0/U_0/U_0/extratemp_reg[2]  ( .D(n10034), .CLK(CLK), .Q(
        \U_0/U_0/U_0/extratemp[2] ) );
  DFFPOSX1 \U_0/U_0/U_0/extratemp_reg[1]  ( .D(n10033), .CLK(CLK), .Q(
        \U_0/U_0/U_0/extratemp[1] ) );
  DFFPOSX1 \U_0/U_0/U_0/extratemp_reg[0]  ( .D(n10032), .CLK(CLK), .Q(
        \U_0/U_0/U_0/extratemp[0] ) );
  DFFPOSX1 \U_0/U_0/U_0/delaydata_reg[7]  ( .D(n10029), .CLK(CLK), .Q(
        \U_0/U_0/U_0/delaydata [7]) );
  DFFPOSX1 \U_0/U_0/U_0/delaydata_reg[0]  ( .D(n10028), .CLK(CLK), .Q(
        \U_0/U_0/U_0/delaydata [0]) );
  DFFPOSX1 \U_0/U_0/U_0/delaydata_reg[1]  ( .D(n10027), .CLK(CLK), .Q(
        \U_0/U_0/U_0/delaydata [1]) );
  DFFPOSX1 \U_0/U_0/U_0/delaydata_reg[2]  ( .D(n10026), .CLK(CLK), .Q(
        \U_0/U_0/U_0/delaydata [2]) );
  DFFPOSX1 \U_0/U_0/U_0/delaydata_reg[3]  ( .D(n10025), .CLK(CLK), .Q(
        \U_0/U_0/U_0/delaydata [3]) );
  DFFPOSX1 \U_0/U_0/U_0/delaydata_reg[4]  ( .D(n10024), .CLK(CLK), .Q(
        \U_0/U_0/U_0/delaydata [4]) );
  DFFPOSX1 \U_0/U_0/U_0/delaydata_reg[5]  ( .D(n10023), .CLK(CLK), .Q(
        \U_0/U_0/U_0/delaydata [5]) );
  DFFPOSX1 \U_0/U_0/U_0/delaydata_reg[6]  ( .D(n10022), .CLK(CLK), .Q(
        \U_0/U_0/U_0/delaydata [6]) );
  DFFSR \U_0/U_0/U_0/sj_reg[7]  ( .D(n8528), .CLK(CLK), .R(n9513), .S(1'b1), 
        .Q(\U_0/U_0/U_0/sj[7] ) );
  DFFSR \U_0/U_0/U_0/sj_reg[6]  ( .D(n8527), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_0/U_0/U_0/sj[6] ) );
  DFFSR \U_0/U_0/U_0/sj_reg[5]  ( .D(n8526), .CLK(CLK), .R(n9514), .S(1'b1), 
        .Q(\U_0/U_0/U_0/sj[5] ) );
  DFFSR \U_0/U_0/U_0/sj_reg[4]  ( .D(n8525), .CLK(CLK), .R(n9520), .S(1'b1), 
        .Q(\U_0/U_0/U_0/sj[4] ) );
  DFFSR \U_0/U_0/U_0/sj_reg[3]  ( .D(n8524), .CLK(CLK), .R(n9490), .S(1'b1), 
        .Q(\U_0/U_0/U_0/sj[3] ) );
  DFFSR \U_0/U_0/U_0/sj_reg[2]  ( .D(n8523), .CLK(CLK), .R(n9524), .S(1'b1), 
        .Q(\U_0/U_0/U_0/sj[2] ) );
  DFFSR \U_0/U_0/U_0/sj_reg[1]  ( .D(n8522), .CLK(CLK), .R(n9526), .S(1'b1), 
        .Q(\U_0/U_0/U_0/sj[1] ) );
  DFFSR \U_0/U_0/U_0/sj_reg[0]  ( .D(n8521), .CLK(CLK), .R(n9523), .S(1'b1), 
        .Q(\U_0/U_0/U_0/sj[0] ) );
  DFFPOSX1 \U_0/U_0/U_0/fw_enable_reg  ( .D(n7462), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fw_enable ) );
  DFFPOSX1 \U_0/U_0/U_0/W_ENABLE_reg  ( .D(n7461), .CLK(CLK), .Q(W_ENABLE_H)
         );
  DFFPOSX1 \U_0/U_0/U_0/temp_reg[6]  ( .D(n8552), .CLK(CLK), .Q(
        \U_0/U_0/U_0/temp[6] ) );
  DFFPOSX1 \U_0/U_0/U_0/temp_reg[0]  ( .D(n8551), .CLK(CLK), .Q(
        \U_0/U_0/U_0/temp[0] ) );
  DFFPOSX1 \U_0/U_0/U_0/temp_reg[1]  ( .D(n8550), .CLK(CLK), .Q(
        \U_0/U_0/U_0/temp[1] ) );
  DFFPOSX1 \U_0/U_0/U_0/temp_reg[2]  ( .D(n8549), .CLK(CLK), .Q(
        \U_0/U_0/U_0/temp[2] ) );
  DFFPOSX1 \U_0/U_0/U_0/temp_reg[3]  ( .D(n8548), .CLK(CLK), .Q(
        \U_0/U_0/U_0/temp[3] ) );
  DFFPOSX1 \U_0/U_0/U_0/temp_reg[4]  ( .D(n8547), .CLK(CLK), .Q(
        \U_0/U_0/U_0/temp[4] ) );
  DFFPOSX1 \U_0/U_0/U_0/temp_reg[5]  ( .D(n8546), .CLK(CLK), .Q(
        \U_0/U_0/U_0/temp[5] ) );
  DFFPOSX1 \U_0/U_0/U_0/temp_reg[7]  ( .D(n8545), .CLK(CLK), .Q(
        \U_0/U_0/U_0/temp[7] ) );
  DFFSR \U_0/U_0/U_0/currentProcessedData_reg[7]  ( .D(
        \U_0/U_0/U_0/nextProcessedData[7] ), .CLK(CLK), .R(n9533), .S(1'b1), 
        .Q(\U_0/U_0/U_0/currentProcessedData [7]) );
  DFFPOSX1 \U_0/U_0/U_0/PROCESSED_DATA_reg[7]  ( .D(n10405), .CLK(CLK), .Q(
        \U_0/PROCESSED_DATA [7]) );
  DFFSR \U_0/U_0/U_0/currentProcessedData_reg[6]  ( .D(
        \U_0/U_0/U_0/nextProcessedData[6] ), .CLK(CLK), .R(n9532), .S(1'b1), 
        .Q(\U_0/U_0/U_0/currentProcessedData [6]) );
  DFFPOSX1 \U_0/U_0/U_0/PROCESSED_DATA_reg[6]  ( .D(n10406), .CLK(CLK), .Q(
        \U_0/PROCESSED_DATA [6]) );
  DFFSR \U_0/U_0/U_0/currentProcessedData_reg[5]  ( .D(
        \U_0/U_0/U_0/nextProcessedData[5] ), .CLK(CLK), .R(n9521), .S(1'b1), 
        .Q(\U_0/U_0/U_0/currentProcessedData [5]) );
  DFFPOSX1 \U_0/U_0/U_0/PROCESSED_DATA_reg[5]  ( .D(n10407), .CLK(CLK), .Q(
        \U_0/PROCESSED_DATA [5]) );
  DFFSR \U_0/U_0/U_0/currentProcessedData_reg[4]  ( .D(
        \U_0/U_0/U_0/nextProcessedData[4] ), .CLK(CLK), .R(n9522), .S(1'b1), 
        .Q(\U_0/U_0/U_0/currentProcessedData [4]) );
  DFFPOSX1 \U_0/U_0/U_0/PROCESSED_DATA_reg[4]  ( .D(n10408), .CLK(CLK), .Q(
        \U_0/PROCESSED_DATA [4]) );
  DFFSR \U_0/U_0/U_0/currentProcessedData_reg[3]  ( .D(
        \U_0/U_0/U_0/nextProcessedData[3] ), .CLK(CLK), .R(n9531), .S(1'b1), 
        .Q(\U_0/U_0/U_0/currentProcessedData [3]) );
  DFFPOSX1 \U_0/U_0/U_0/PROCESSED_DATA_reg[3]  ( .D(n10409), .CLK(CLK), .Q(
        \U_0/PROCESSED_DATA [3]) );
  DFFSR \U_0/U_0/U_0/currentProcessedData_reg[2]  ( .D(
        \U_0/U_0/U_0/nextProcessedData[2] ), .CLK(CLK), .R(n9534), .S(1'b1), 
        .Q(\U_0/U_0/U_0/currentProcessedData [2]) );
  DFFPOSX1 \U_0/U_0/U_0/PROCESSED_DATA_reg[2]  ( .D(n10410), .CLK(CLK), .Q(
        \U_0/PROCESSED_DATA [2]) );
  DFFSR \U_0/U_0/U_0/currentProcessedData_reg[1]  ( .D(
        \U_0/U_0/U_0/nextProcessedData[1] ), .CLK(CLK), .R(n9488), .S(1'b1), 
        .Q(\U_0/U_0/U_0/currentProcessedData [1]) );
  DFFPOSX1 \U_0/U_0/U_0/PROCESSED_DATA_reg[1]  ( .D(n10411), .CLK(CLK), .Q(
        \U_0/PROCESSED_DATA [1]) );
  DFFSR \U_0/U_0/U_0/currentProcessedData_reg[0]  ( .D(
        \U_0/U_0/U_0/nextProcessedData[0] ), .CLK(CLK), .R(n9527), .S(1'b1), 
        .Q(\U_0/U_0/U_0/currentProcessedData [0]) );
  DFFPOSX1 \U_0/U_0/U_0/PROCESSED_DATA_reg[0]  ( .D(n10412), .CLK(CLK), .Q(
        \U_0/PROCESSED_DATA [0]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[15]  ( .D(n8472), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [15]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[1]  ( .D(n8486), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [1]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[9]  ( .D(n8478), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [9]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[2]  ( .D(n8485), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [2]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[10]  ( .D(n8477), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [10]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[3]  ( .D(n8484), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [3]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[11]  ( .D(n8476), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [11]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[4]  ( .D(n8483), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [4]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[12]  ( .D(n8475), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [12]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[5]  ( .D(n8482), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [5]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[13]  ( .D(n8474), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [13]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[6]  ( .D(n8481), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [6]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[14]  ( .D(n8473), .CLK(CLK), .R(n9489), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [14]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[7]  ( .D(n8480), .CLK(CLK), .R(n9489), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [7]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[0]  ( .D(n8487), .CLK(CLK), .R(n9489), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [0]) );
  DFFSR \U_0/U_3/U_1/current_crc_reg[8]  ( .D(n8479), .CLK(CLK), .R(n9489), 
        .S(1'b1), .Q(\U_0/U_3/TX_CRC [8]) );
  DFFPOSX1 \U_0/U_0/U_0/fdata_reg[6]  ( .D(n7428), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fdata [6]) );
  DFFPOSX1 \U_0/U_0/U_0/DATA_reg[6]  ( .D(n7427), .CLK(CLK), .Q(DATA_H[6]) );
  DFFPOSX1 \U_0/U_0/U_0/fdata_reg[5]  ( .D(n7426), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fdata [5]) );
  DFFPOSX1 \U_0/U_0/U_0/DATA_reg[5]  ( .D(n7425), .CLK(CLK), .Q(DATA_H[5]) );
  DFFPOSX1 \U_0/U_0/U_0/fdata_reg[4]  ( .D(n7424), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fdata [4]) );
  DFFPOSX1 \U_0/U_0/U_0/DATA_reg[4]  ( .D(n7423), .CLK(CLK), .Q(DATA_H[4]) );
  DFFPOSX1 \U_0/U_0/U_0/fdata_reg[3]  ( .D(n7422), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fdata [3]) );
  DFFPOSX1 \U_0/U_0/U_0/DATA_reg[3]  ( .D(n7421), .CLK(CLK), .Q(DATA_H[3]) );
  DFFPOSX1 \U_0/U_0/U_0/fdata_reg[2]  ( .D(n7420), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fdata [2]) );
  DFFPOSX1 \U_0/U_0/U_0/DATA_reg[2]  ( .D(n7419), .CLK(CLK), .Q(DATA_H[2]) );
  DFFPOSX1 \U_0/U_0/U_0/fdata_reg[1]  ( .D(n7418), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fdata [1]) );
  DFFPOSX1 \U_0/U_0/U_0/DATA_reg[1]  ( .D(n7417), .CLK(CLK), .Q(DATA_H[1]) );
  DFFPOSX1 \U_0/U_0/U_0/fdata_reg[0]  ( .D(n7416), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fdata [0]) );
  DFFPOSX1 \U_0/U_0/U_0/DATA_reg[0]  ( .D(n7415), .CLK(CLK), .Q(DATA_H[0]) );
  DFFPOSX1 \U_0/U_0/U_0/fr_enable_reg  ( .D(n7414), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fr_enable ) );
  DFFPOSX1 \U_0/U_0/U_0/R_ENABLE_reg  ( .D(n7413), .CLK(CLK), .Q(R_ENABLE_H)
         );
  DFFSR \U_0/U_0/U_0/si_reg[7]  ( .D(n8510), .CLK(CLK), .R(n9489), .S(1'b1), 
        .Q(\U_0/U_0/U_0/si[7] ) );
  DFFSR \U_0/U_0/U_0/si_reg[0]  ( .D(n8520), .CLK(CLK), .R(n9489), .S(1'b1), 
        .Q(\U_0/U_0/U_0/si[0] ) );
  DFFSR \U_0/U_0/U_0/si_reg[1]  ( .D(n8518), .CLK(CLK), .R(n9489), .S(1'b1), 
        .Q(\U_0/U_0/U_0/si[1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyi_reg[1]  ( .D(n8517), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyi[1] ) );
  DFFSR \U_0/U_0/U_0/si_reg[2]  ( .D(n8516), .CLK(CLK), .R(n9489), .S(1'b1), 
        .Q(\U_0/U_0/U_0/si[2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyi_reg[2]  ( .D(n8515), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyi[2] ) );
  DFFSR \U_0/U_0/U_0/si_reg[3]  ( .D(n8514), .CLK(CLK), .R(n9489), .S(1'b1), 
        .Q(\U_0/U_0/U_0/si[3] ) );
  DFFSR \U_0/U_0/U_0/si_reg[4]  ( .D(n8513), .CLK(CLK), .R(n9489), .S(1'b1), 
        .Q(\U_0/U_0/U_0/si[4] ) );
  DFFSR \U_0/U_0/U_0/si_reg[5]  ( .D(n8512), .CLK(CLK), .R(n9489), .S(1'b1), 
        .Q(\U_0/U_0/U_0/si[5] ) );
  DFFSR \U_0/U_0/U_0/si_reg[6]  ( .D(n8511), .CLK(CLK), .R(n9489), .S(1'b1), 
        .Q(\U_0/U_0/U_0/si[6] ) );
  DFFPOSX1 \U_0/U_0/U_0/ADDR_reg[0]  ( .D(n7404), .CLK(CLK), .Q(ADDR_H[0]) );
  DFFPOSX1 \U_0/U_0/U_0/faddr_reg[0]  ( .D(n10413), .CLK(CLK), .Q(
        \U_0/U_0/U_0/faddr [0]) );
  DFFPOSX1 \U_0/U_0/U_0/ADDR_reg[1]  ( .D(n7402), .CLK(CLK), .Q(ADDR_H[1]) );
  DFFPOSX1 \U_0/U_0/U_0/faddr_reg[1]  ( .D(n10414), .CLK(CLK), .Q(
        \U_0/U_0/U_0/faddr [1]) );
  DFFPOSX1 \U_0/U_0/U_0/ADDR_reg[2]  ( .D(n7400), .CLK(CLK), .Q(ADDR_H[2]) );
  DFFPOSX1 \U_0/U_0/U_0/faddr_reg[2]  ( .D(n10415), .CLK(CLK), .Q(
        \U_0/U_0/U_0/faddr [2]) );
  DFFPOSX1 \U_0/U_0/U_0/ADDR_reg[3]  ( .D(n7398), .CLK(CLK), .Q(ADDR_H[3]) );
  DFFPOSX1 \U_0/U_0/U_0/faddr_reg[3]  ( .D(n10416), .CLK(CLK), .Q(
        \U_0/U_0/U_0/faddr [3]) );
  DFFPOSX1 \U_0/U_0/U_0/ADDR_reg[4]  ( .D(n7396), .CLK(CLK), .Q(ADDR_H[4]) );
  DFFPOSX1 \U_0/U_0/U_0/faddr_reg[4]  ( .D(n10417), .CLK(CLK), .Q(
        \U_0/U_0/U_0/faddr [4]) );
  DFFPOSX1 \U_0/U_0/U_0/ADDR_reg[5]  ( .D(n7394), .CLK(CLK), .Q(ADDR_H[5]) );
  DFFPOSX1 \U_0/U_0/U_0/faddr_reg[5]  ( .D(n10418), .CLK(CLK), .Q(
        \U_0/U_0/U_0/faddr [5]) );
  DFFPOSX1 \U_0/U_0/U_0/ADDR_reg[6]  ( .D(n7392), .CLK(CLK), .Q(ADDR_H[6]) );
  DFFPOSX1 \U_0/U_0/U_0/faddr_reg[6]  ( .D(n10419), .CLK(CLK), .Q(
        \U_0/U_0/U_0/faddr [6]) );
  DFFPOSX1 \U_0/U_0/U_0/ADDR_reg[7]  ( .D(n7390), .CLK(CLK), .Q(ADDR_H[7]) );
  DFFPOSX1 \U_0/U_0/U_0/faddr_reg[7]  ( .D(n10420), .CLK(CLK), .Q(
        \U_0/U_0/U_0/faddr [7]) );
  DFFPOSX1 \U_0/U_0/U_0/keyi_reg[0]  ( .D(n8519), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyi[0] ) );
  DFFPOSX1 \U_0/U_0/U_0/fdata_reg[7]  ( .D(n7388), .CLK(CLK), .Q(
        \U_0/U_0/U_0/fdata [7]) );
  DFFPOSX1 \U_0/U_0/U_0/DATA_reg[7]  ( .D(n7387), .CLK(CLK), .Q(DATA_H[7]) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[0][6]  ( .D(n9952), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[0][6] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[0][5]  ( .D(n9953), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[0][5] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[0][4]  ( .D(n9954), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[0][4] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[0][3]  ( .D(n8564), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[0][3] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[0][2]  ( .D(n8565), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[0][2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[0][1]  ( .D(n8566), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[0][1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[0][0]  ( .D(n8567), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[0][0] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[1][7]  ( .D(n9955), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[1][7] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[0][7]  ( .D(n9956), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[0][7] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[7][0]  ( .D(n9957), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[7][0] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[7][1]  ( .D(n9958), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[7][1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[7][2]  ( .D(n9959), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[7][2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[7][3]  ( .D(n9960), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[7][3] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[7][4]  ( .D(n9961), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[7][4] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[7][5]  ( .D(n9962), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[7][5] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[7][6]  ( .D(n9963), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[7][6] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[7][7]  ( .D(n9964), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[7][7] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[6][0]  ( .D(n9965), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[6][0] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[6][1]  ( .D(n9966), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[6][1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[6][2]  ( .D(n9967), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[6][2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[6][3]  ( .D(n9968), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[6][3] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[6][4]  ( .D(n9969), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[6][4] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[6][5]  ( .D(n9970), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[6][5] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[6][6]  ( .D(n9971), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[6][6] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[6][7]  ( .D(n9972), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[6][7] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[5][0]  ( .D(n9973), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[5][0] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[5][1]  ( .D(n9974), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[5][1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[5][2]  ( .D(n9975), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[5][2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[5][3]  ( .D(n9976), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[5][3] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[5][4]  ( .D(n9977), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[5][4] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[5][5]  ( .D(n9978), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[5][5] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[5][6]  ( .D(n9979), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[5][6] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[5][7]  ( .D(n9980), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[5][7] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[4][0]  ( .D(n9981), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[4][0] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[4][1]  ( .D(n9982), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[4][1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[4][2]  ( .D(n9983), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[4][2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[4][3]  ( .D(n9984), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[4][3] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[4][4]  ( .D(n9985), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[4][4] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[4][5]  ( .D(n9986), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[4][5] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[4][6]  ( .D(n9987), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[4][6] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[4][7]  ( .D(n9988), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[4][7] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[3][0]  ( .D(n9989), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[3][0] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[3][1]  ( .D(n9990), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[3][1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[3][2]  ( .D(n9991), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[3][2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[3][3]  ( .D(n9992), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[3][3] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[3][4]  ( .D(n9993), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[3][4] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[3][5]  ( .D(n9994), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[3][5] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[3][6]  ( .D(n9995), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[3][6] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[3][7]  ( .D(n9996), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[3][7] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[2][0]  ( .D(n9997), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[2][0] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[2][1]  ( .D(n9998), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[2][1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[2][2]  ( .D(n9999), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[2][2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[2][3]  ( .D(n10000), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[2][3] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[2][4]  ( .D(n10001), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[2][4] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[2][5]  ( .D(n10002), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[2][5] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[2][6]  ( .D(n10003), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[2][6] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[2][7]  ( .D(n10004), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[2][7] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[1][0]  ( .D(n10005), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[1][0] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[1][1]  ( .D(n10006), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[1][1] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[1][2]  ( .D(n10007), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[1][2] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[1][3]  ( .D(n10008), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[1][3] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[1][4]  ( .D(n10009), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[1][4] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[1][5]  ( .D(n10010), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[1][5] ) );
  DFFPOSX1 \U_0/U_0/U_0/keyTable_reg[1][6]  ( .D(n10011), .CLK(CLK), .Q(
        \U_0/U_0/U_0/keyTable[1][6] ) );
  DFFPOSX1 \U_0/U_1/U_0/tempOpcode_reg[1]  ( .D(n7386), .CLK(CLK), .Q(
        \U_0/U_1/U_0/tempOpcode [1]) );
  DFFPOSX1 \U_0/U_3/U_3/flop_data_reg[7]  ( .D(n7750), .CLK(CLK), .Q(
        \U_0/U_3/U_3/flop_data [7]) );
  DFFPOSX1 \U_0/U_3/U_3/flop_data_reg[0]  ( .D(n10050), .CLK(CLK), .Q(
        \U_0/U_3/U_3/flop_data [0]) );
  DFFPOSX1 \U_0/U_3/U_3/flop_data_reg[1]  ( .D(n10049), .CLK(CLK), .Q(
        \U_0/U_3/U_3/flop_data [1]) );
  DFFPOSX1 \U_0/U_3/U_3/flop_data_reg[2]  ( .D(n10048), .CLK(CLK), .Q(
        \U_0/U_3/U_3/flop_data [2]) );
  DFFPOSX1 \U_0/U_3/U_3/flop_data_reg[3]  ( .D(n10047), .CLK(CLK), .Q(
        \U_0/U_3/U_3/flop_data [3]) );
  DFFPOSX1 \U_0/U_3/U_3/flop_data_reg[4]  ( .D(n10046), .CLK(CLK), .Q(
        \U_0/U_3/U_3/flop_data [4]) );
  DFFPOSX1 \U_0/U_3/U_3/flop_data_reg[5]  ( .D(n10045), .CLK(CLK), .Q(
        \U_0/U_3/U_3/flop_data [5]) );
  DFFPOSX1 \U_0/U_3/U_3/flop_data_reg[6]  ( .D(n10044), .CLK(CLK), .Q(
        \U_0/U_3/U_3/flop_data [6]) );
  DFFPOSX1 \U_0/U_3/U_3/current_send_data_reg[6]  ( .D(n7385), .CLK(CLK), .Q(
        \U_0/U_3/U_3/current_send_data [6]) );
  DFFPOSX1 \U_0/U_3/U_3/send_data_reg[6]  ( .D(n7384), .CLK(CLK), .Q(
        \U_0/U_3/send_data [6]) );
  DFFPOSX1 \U_0/U_3/U_3/current_send_data_reg[5]  ( .D(n7383), .CLK(CLK), .Q(
        \U_0/U_3/U_3/current_send_data [5]) );
  DFFPOSX1 \U_0/U_3/U_3/send_data_reg[5]  ( .D(n7382), .CLK(CLK), .Q(
        \U_0/U_3/send_data [5]) );
  DFFPOSX1 \U_0/U_3/U_3/current_send_data_reg[4]  ( .D(n7381), .CLK(CLK), .Q(
        \U_0/U_3/U_3/current_send_data [4]) );
  DFFPOSX1 \U_0/U_3/U_3/send_data_reg[4]  ( .D(n7380), .CLK(CLK), .Q(
        \U_0/U_3/send_data [4]) );
  DFFPOSX1 \U_0/U_3/U_3/current_send_data_reg[3]  ( .D(n7379), .CLK(CLK), .Q(
        \U_0/U_3/U_3/current_send_data [3]) );
  DFFPOSX1 \U_0/U_3/U_3/send_data_reg[3]  ( .D(n7378), .CLK(CLK), .Q(
        \U_0/U_3/send_data [3]) );
  DFFPOSX1 \U_0/U_3/U_3/current_send_data_reg[2]  ( .D(n7377), .CLK(CLK), .Q(
        \U_0/U_3/U_3/current_send_data [2]) );
  DFFPOSX1 \U_0/U_3/U_3/send_data_reg[2]  ( .D(n7376), .CLK(CLK), .Q(
        \U_0/U_3/send_data [2]) );
  DFFPOSX1 \U_0/U_3/U_3/current_send_data_reg[1]  ( .D(n7375), .CLK(CLK), .Q(
        \U_0/U_3/U_3/current_send_data [1]) );
  DFFPOSX1 \U_0/U_3/U_3/send_data_reg[1]  ( .D(n7374), .CLK(CLK), .Q(
        \U_0/U_3/send_data [1]) );
  DFFPOSX1 \U_0/U_3/U_3/current_send_data_reg[0]  ( .D(n7373), .CLK(CLK), .Q(
        \U_0/U_3/U_3/current_send_data [0]) );
  DFFPOSX1 \U_0/U_3/U_3/send_data_reg[0]  ( .D(n7372), .CLK(CLK), .Q(
        \U_0/U_3/send_data [0]) );
  DFFPOSX1 \U_0/U_3/U_3/current_send_data_reg[7]  ( .D(n7371), .CLK(CLK), .Q(
        \U_0/U_3/U_3/current_send_data [7]) );
  DFFPOSX1 \U_0/U_3/U_3/send_data_reg[7]  ( .D(n7370), .CLK(CLK), .Q(
        \U_0/U_3/send_data [7]) );
  DFFSR \U_0/U_3/U_4/state_reg  ( .D(host_is_sending), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_0/U_3/U_4/state ) );
  DFFSR \U_0/U_3/U_4/count_reg[0]  ( .D(\U_0/U_3/U_4/nextcount [0]), .CLK(CLK), 
        .R(n9490), .S(1'b1), .Q(\U_0/U_3/U_4/count[0] ) );
  DFFSR \U_0/U_3/U_4/count_reg[2]  ( .D(\U_0/U_3/U_4/nextcount [2]), .CLK(CLK), 
        .R(n9490), .S(1'b1), .Q(\U_0/U_3/U_4/count[2] ) );
  DFFSR \U_0/U_3/U_4/count_reg[3]  ( .D(\U_0/U_3/U_4/nextcount [3]), .CLK(CLK), 
        .R(n9490), .S(1'b1), .Q(\U_0/U_3/U_4/count[3] ) );
  DFFSR \U_0/U_3/U_4/count_reg[1]  ( .D(\U_0/U_3/U_4/nextcount [1]), .CLK(CLK), 
        .R(n9490), .S(1'b1), .Q(\U_0/U_3/U_4/count[1] ) );
  DFFSR \U_0/U_3/U_2/count_reg[1]  ( .D(n8470), .CLK(CLK), .R(1'b1), .S(n9521), 
        .Q(\U_0/U_3/U_2/count[1] ) );
  DFFSR \U_0/U_3/U_2/count_reg[2]  ( .D(n8469), .CLK(CLK), .R(1'b1), .S(n9521), 
        .Q(\U_0/U_3/U_2/count[2] ) );
  DFFSR \U_0/U_3/U_2/count_reg[0]  ( .D(n10873), .CLK(CLK), .R(1'b1), .S(n9521), .Q(\U_0/U_3/U_2/count[0] ) );
  DFFSR \U_0/U_3/U_2/present_val_reg[7]  ( .D(n10874), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_0/U_3/U_2/present_val [7]) );
  DFFSR \U_0/U_3/U_2/present_val_reg[6]  ( .D(n8462), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_0/U_3/U_2/present_val [6]) );
  DFFSR \U_0/U_3/U_2/present_val_reg[5]  ( .D(n8463), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_0/U_3/U_2/present_val [5]) );
  DFFSR \U_0/U_3/U_2/present_val_reg[4]  ( .D(n8464), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_0/U_3/U_2/present_val [4]) );
  DFFSR \U_0/U_3/U_2/present_val_reg[3]  ( .D(n8465), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_0/U_3/U_2/present_val [3]) );
  DFFSR \U_0/U_3/U_2/present_val_reg[2]  ( .D(n8466), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_0/U_3/U_2/present_val [2]) );
  DFFSR \U_0/U_3/U_2/present_val_reg[1]  ( .D(n8467), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_0/U_3/U_2/present_val [1]) );
  DFFSR \U_0/U_3/U_2/present_val_reg[0]  ( .D(n8468), .CLK(CLK), .R(n9491), 
        .S(1'b1), .Q(\U_0/U_3/d_encode ) );
  DFFSR \U_0/U_3/U_0/DE_holdout_BS_reg  ( .D(n8460), .CLK(CLK), .R(n9491), .S(
        1'b1), .Q(\U_0/U_3/U_0/DE_holdout_BS ) );
  DFFSR \U_0/U_3/U_0/dm_tx_out_reg  ( .D(\U_0/U_3/U_0/dm_tx_nxt ), .CLK(CLK), 
        .R(n9491), .S(1'b1), .Q(DMTS) );
  DFFSR \U_1/U_0/U_1/U_0/Q_int_reg  ( .D(SERIAL_IN), .CLK(CLK), .R(n9491), .S(
        1'b1), .Q(\U_1/U_0/U_1/U_0/Q_int ) );
  DFFSR \U_1/U_0/U_1/U_0/Q_int2_reg  ( .D(\U_1/U_0/U_1/U_0/Q_int ), .CLK(CLK), 
        .R(n9491), .S(1'b1), .Q(\U_1/U_0/U_1/U_0/Q_int2 ) );
  DFFSR \U_1/U_0/U_1/U_7/nextState_reg[7]  ( .D(n8459), .CLK(CLK), .R(n9491), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_7/nextState[7] ) );
  DFFSR \U_1/U_0/U_1/U_7/state_reg[7]  ( .D(\U_1/U_0/U_1/U_7/nextState[7] ), 
        .CLK(CLK), .R(n9491), .S(1'b1), .Q(\U_1/U_0/U_1/U_7/state[7] ) );
  DFFSR \U_1/U_0/U_1/U_7/nextState_reg[6]  ( .D(n8458), .CLK(CLK), .R(n9491), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_7/nextState[6] ) );
  DFFSR \U_1/U_0/U_1/U_7/state_reg[6]  ( .D(\U_1/U_0/U_1/U_7/nextState[6] ), 
        .CLK(CLK), .R(n9491), .S(1'b1), .Q(\U_1/U_0/U_1/U_7/state[6] ) );
  DFFSR \U_1/U_0/U_1/U_7/nextState_reg[5]  ( .D(n8457), .CLK(CLK), .R(n9491), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_7/nextState[5] ) );
  DFFSR \U_1/U_0/U_1/U_7/state_reg[5]  ( .D(\U_1/U_0/U_1/U_7/nextState[5] ), 
        .CLK(CLK), .R(n9491), .S(1'b1), .Q(\U_1/U_0/U_1/U_7/state[5] ) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[9]  ( .D(n8451), .CLK(CLK), .R(n9491), 
        .S(1'b1), .Q(\U_1/U_0/U_1/STOP_DATA [1]) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[8]  ( .D(n8450), .CLK(CLK), .R(n9492), 
        .S(1'b1), .Q(\U_1/U_0/U_1/STOP_DATA [0]) );
  DFFSR \U_1/U_0/U_1/U_5/SB_DETECT_reg  ( .D(\U_1/U_0/U_1/U_5/sb_detect_flag ), 
        .CLK(CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/SB_DETECT ) );
  DFFSR \U_1/U_0/U_1/U_2/state_reg[0]  ( .D(\U_1/U_0/U_1/U_2/nextState[0] ), 
        .CLK(CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/state[0] ) );
  DFFSR \U_1/U_0/U_1/U_2/timerRunning_reg  ( .D(n8449), .CLK(CLK), .R(n9492), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_2/timerRunning ) );
  DFFSR \U_1/U_0/U_1/U_2/nextCount_reg[1]  ( .D(\U_1/U_0/U_1/U_2/N32 ), .CLK(
        CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/nextCount [1]) );
  DFFSR \U_1/U_0/U_1/U_2/count_reg[1]  ( .D(\U_1/U_0/U_1/U_2/nextCount [1]), 
        .CLK(CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/count[1] ) );
  DFFSR \U_1/U_0/U_1/U_2/nextCount_reg[0]  ( .D(\U_1/U_0/U_1/U_2/N31 ), .CLK(
        CLK), .R(1'b1), .S(n9522), .Q(\U_1/U_0/U_1/U_2/nextCount [0]) );
  DFFSR \U_1/U_0/U_1/U_2/count_reg[0]  ( .D(\U_1/U_0/U_1/U_2/nextCount [0]), 
        .CLK(CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/N23 ) );
  DFFSR \U_1/U_0/U_1/U_2/nextCount_reg[2]  ( .D(\U_1/U_0/U_1/U_2/N33 ), .CLK(
        CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/nextCount [2]) );
  DFFSR \U_1/U_0/U_1/U_2/count_reg[2]  ( .D(\U_1/U_0/U_1/U_2/nextCount [2]), 
        .CLK(CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/count[2] ) );
  DFFSR \U_1/U_0/U_1/U_2/nextCount_reg[3]  ( .D(\U_1/U_0/U_1/U_2/N34 ), .CLK(
        CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/nextCount [3]) );
  DFFSR \U_1/U_0/U_1/U_2/count_reg[3]  ( .D(\U_1/U_0/U_1/U_2/nextCount [3]), 
        .CLK(CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/count[3] ) );
  DFFSR \U_1/U_0/U_1/U_2/nextCount_reg[4]  ( .D(\U_1/U_0/U_1/U_2/N35 ), .CLK(
        CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/nextCount [4]) );
  DFFSR \U_1/U_0/U_1/U_2/count_reg[4]  ( .D(\U_1/U_0/U_1/U_2/nextCount [4]), 
        .CLK(CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/count[4] ) );
  DFFSR \U_1/U_0/U_1/U_2/nextCount_reg[5]  ( .D(\U_1/U_0/U_1/U_2/N36 ), .CLK(
        CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/nextCount [5]) );
  DFFSR \U_1/U_0/U_1/U_2/count_reg[5]  ( .D(\U_1/U_0/U_1/U_2/nextCount [5]), 
        .CLK(CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/count[5] ) );
  DFFSR \U_1/U_0/U_1/U_2/nextCount_reg[6]  ( .D(\U_1/U_0/U_1/U_2/N37 ), .CLK(
        CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/nextCount [6]) );
  DFFSR \U_1/U_0/U_1/U_2/count_reg[6]  ( .D(\U_1/U_0/U_1/U_2/nextCount [6]), 
        .CLK(CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/count[6] ) );
  DFFSR \U_1/U_0/U_1/U_2/nextCount_reg[7]  ( .D(\U_1/U_0/U_1/U_2/N38 ), .CLK(
        CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/nextCount [7]) );
  DFFSR \U_1/U_0/U_1/U_2/count_reg[7]  ( .D(\U_1/U_0/U_1/U_2/nextCount [7]), 
        .CLK(CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/count[7] ) );
  DFFSR \U_1/U_0/U_1/U_2/state_reg[1]  ( .D(\U_1/U_0/U_1/U_2/nextState[1] ), 
        .CLK(CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/state[1] ) );
  DFFSR \U_1/U_0/U_1/U_2/state_reg[2]  ( .D(\U_1/U_0/U_1/U_2/nextState[2] ), 
        .CLK(CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_2/state[2] ) );
  DFFSR \U_1/U_0/U_1/U_2/RBUF_LOAD_reg  ( .D(n8446), .CLK(CLK), .R(n9493), .S(
        1'b1), .Q(\U_1/U_0/U_1/RBUF_LOAD ) );
  DFFSR \U_1/U_0/U_1/U_2/SET_RBUF_FULL_reg  ( .D(n8443), .CLK(CLK), .R(n9493), 
        .S(1'b1), .Q(\U_1/U_0/U_1/SET_RBUF_FULL ) );
  DFFSR \U_1/U_0/U_1/U_2/CHK_ERROR_reg  ( .D(n8447), .CLK(CLK), .R(n9493), .S(
        1'b1), .Q(\U_1/U_0/U_1/CHK_ERROR ) );
  DFFSR \U_1/U_0/U_1/U_2/SBC_CLR_reg  ( .D(n8444), .CLK(CLK), .R(n9489), .S(
        1'b1), .Q(\U_1/U_0/U_1/SBC_CLR ) );
  DFFSR \U_1/U_0/U_1/U_2/TIMER_TRIG_reg  ( .D(n8445), .CLK(CLK), .R(n9530), 
        .S(1'b1), .Q(\U_1/U_0/U_1/TIMER_TRIG ) );
  DFFSR \U_1/U_0/U_1/U_7/nextState_reg[0]  ( .D(n8452), .CLK(CLK), .R(n9525), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_7/nextState[0] ) );
  DFFSR \U_1/U_0/U_1/U_7/state_reg[0]  ( .D(\U_1/U_0/U_1/U_7/nextState[0] ), 
        .CLK(CLK), .R(n9491), .S(1'b1), .Q(\U_1/U_0/U_1/U_7/state[0] ) );
  DFFSR \U_1/U_0/U_1/U_7/nextState_reg[1]  ( .D(n8453), .CLK(CLK), .R(n9488), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_7/nextState[1] ) );
  DFFSR \U_1/U_0/U_1/U_7/state_reg[1]  ( .D(\U_1/U_0/U_1/U_7/nextState[1] ), 
        .CLK(CLK), .R(n9492), .S(1'b1), .Q(\U_1/U_0/U_1/U_7/state[1] ) );
  DFFSR \U_1/U_0/U_1/U_7/nextState_reg[2]  ( .D(n8454), .CLK(CLK), .R(n9533), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_7/nextState[2] ) );
  DFFSR \U_1/U_0/U_1/U_7/state_reg[2]  ( .D(\U_1/U_0/U_1/U_7/nextState[2] ), 
        .CLK(CLK), .R(n9493), .S(1'b1), .Q(\U_1/U_0/U_1/U_7/state[2] ) );
  DFFSR \U_1/U_0/U_1/U_7/nextState_reg[3]  ( .D(n8455), .CLK(CLK), .R(n9521), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_7/nextState[3] ) );
  DFFSR \U_1/U_0/U_1/U_7/state_reg[3]  ( .D(\U_1/U_0/U_1/U_7/nextState[3] ), 
        .CLK(CLK), .R(n9494), .S(1'b1), .Q(\U_1/U_0/U_1/U_7/state[3] ) );
  DFFSR \U_1/U_0/U_1/U_7/nextState_reg[4]  ( .D(n8456), .CLK(CLK), .R(n9532), 
        .S(1'b1), .Q(\U_1/U_0/U_1/U_7/nextState[4] ) );
  DFFSR \U_1/U_0/U_1/U_7/state_reg[4]  ( .D(\U_1/U_0/U_1/U_7/nextState[4] ), 
        .CLK(CLK), .R(n9494), .S(1'b1), .Q(\U_1/U_0/U_1/U_7/state[4] ) );
  DFFSR \U_1/U_0/U_1/U_2/SBC_EN_reg  ( .D(n8448), .CLK(CLK), .R(n9494), .S(
        1'b1), .Q(\U_1/U_0/U_1/SBC_EN ) );
  DFFSR \U_1/U_0/U_1/U_5/SBE_reg  ( .D(\U_1/U_0/U_1/U_5/SBE_prime ), .CLK(CLK), 
        .R(n9494), .S(1'b1), .Q(\U_1/U_0/U_1/SBE ) );
  DFFSR \U_1/U_0/U_1/U_8/state_reg[0]  ( .D(n8441), .CLK(CLK), .R(n9494), .S(
        1'b1), .Q(\U_1/U_0/U_1/U_8/state[0] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/keyCount_reg[1]  ( .D(n8437), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/keyCount[1] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/keyCount_reg[2]  ( .D(n8436), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/keyCount[2] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/keyCount_reg[3]  ( .D(n8435), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/keyCount[3] ) );
  DFFSR \U_1/U_0/U_1/U_8/state_reg[2]  ( .D(n8442), .CLK(CLK), .R(n9494), .S(
        1'b1), .Q(\U_1/U_0/U_1/U_8/state[2] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/keyCount_reg[0]  ( .D(n8438), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/keyCount[0] ) );
  DFFSR \U_1/U_0/U_1/U_8/state_reg[3]  ( .D(n8440), .CLK(CLK), .R(n9494), .S(
        1'b1), .Q(\U_1/U_0/U_1/U_8/state[3] ) );
  DFFSR \U_1/U_0/U_1/U_8/state_reg[1]  ( .D(n8439), .CLK(CLK), .R(n9494), .S(
        1'b1), .Q(\U_1/U_0/U_1/U_8/state[1] ) );
  DFFSR \U_1/U_0/U_1/U_4/Q_int_reg  ( .D(n7299), .CLK(CLK), .R(n7749), .S(1'b1), .Q(\U_1/RBUF_FULL ) );
  DFFSR \U_1/U_0/U_1/U_1/OE_reg  ( .D(\U_1/U_0/U_1/U_1/OE_prime ), .CLK(CLK), 
        .R(n9494), .S(1'b1), .Q(\U_1/U_0/U_1/OE ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/address_reg[0]  ( .D(n8427), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/address[0] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/address_reg[1]  ( .D(n8428), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/address[1] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/address_reg[2]  ( .D(n8429), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/address[2] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/address_reg[6]  ( .D(n8433), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/address[6] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/address_reg[7]  ( .D(n8434), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/address[7] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/address_reg[3]  ( .D(n8430), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/address[3] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/address_reg[5]  ( .D(n8432), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/address[5] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/address_reg[4]  ( .D(n8431), .CLK(CLK), .Q(
        \U_1/U_0/U_1/U_8/address[4] ) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[7]  ( .D(n8426), .CLK(CLK), .R(n9494), 
        .S(1'b1), .Q(\U_1/U_0/U_1/LOAD_DATA [7]) );
  DFFSR \U_1/U_0/U_1/U_3/Q_int_reg[7]  ( .D(n7295), .CLK(CLK), .R(n9494), .S(
        1'b1), .Q(\U_1/U_0/U_1/RCV_DATA [7]) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[6]  ( .D(n8425), .CLK(CLK), .R(n9494), 
        .S(1'b1), .Q(\U_1/U_0/U_1/LOAD_DATA [6]) );
  DFFSR \U_1/U_0/U_1/U_3/Q_int_reg[6]  ( .D(n11327), .CLK(CLK), .R(n9494), .S(
        1'b1), .Q(\U_1/U_0/U_1/RCV_DATA [6]) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[5]  ( .D(n8424), .CLK(CLK), .R(n9495), 
        .S(1'b1), .Q(\U_1/U_0/U_1/LOAD_DATA [5]) );
  DFFSR \U_1/U_0/U_1/U_3/Q_int_reg[5]  ( .D(n7289), .CLK(CLK), .R(n9495), .S(
        1'b1), .Q(\U_1/U_0/U_1/RCV_DATA [5]) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[4]  ( .D(n8423), .CLK(CLK), .R(n9495), 
        .S(1'b1), .Q(\U_1/U_0/U_1/LOAD_DATA [4]) );
  DFFSR \U_1/U_0/U_1/U_3/Q_int_reg[4]  ( .D(n7286), .CLK(CLK), .R(n9495), .S(
        1'b1), .Q(\U_1/U_0/U_1/RCV_DATA [4]) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[3]  ( .D(n8422), .CLK(CLK), .R(n9495), 
        .S(1'b1), .Q(\U_1/U_0/U_1/LOAD_DATA [3]) );
  DFFSR \U_1/U_0/U_1/U_3/Q_int_reg[3]  ( .D(n7283), .CLK(CLK), .R(n9495), .S(
        1'b1), .Q(\U_1/U_0/U_1/RCV_DATA [3]) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[2]  ( .D(n8421), .CLK(CLK), .R(n9495), 
        .S(1'b1), .Q(\U_1/U_0/U_1/LOAD_DATA [2]) );
  DFFSR \U_1/U_0/U_1/U_3/Q_int_reg[2]  ( .D(n7280), .CLK(CLK), .R(n9495), .S(
        1'b1), .Q(\U_1/U_0/U_1/RCV_DATA [2]) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[1]  ( .D(n8420), .CLK(CLK), .R(n9495), 
        .S(1'b1), .Q(\U_1/U_0/U_1/LOAD_DATA [1]) );
  DFFSR \U_1/U_0/U_1/U_3/Q_int_reg[1]  ( .D(n7277), .CLK(CLK), .R(n9495), .S(
        1'b1), .Q(\U_1/U_0/U_1/RCV_DATA [1]) );
  DFFSR \U_1/U_0/U_1/U_6/present_val_reg[0]  ( .D(n8419), .CLK(CLK), .R(n9495), 
        .S(1'b1), .Q(\U_1/U_0/U_1/LOAD_DATA [0]) );
  DFFSR \U_1/U_0/U_1/U_3/Q_int_reg[0]  ( .D(n7274), .CLK(CLK), .R(n9495), .S(
        1'b1), .Q(\U_1/U_0/U_1/RCV_DATA [0]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/parityAccumulator_reg[0]  ( .D(n8418), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/parityAccumulator[0] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/parityAccumulator_reg[1]  ( .D(n8417), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/parityAccumulator[1] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/parityAccumulator_reg[2]  ( .D(n8416), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/parityAccumulator[2] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/parityAccumulator_reg[3]  ( .D(n8415), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/parityAccumulator[3] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/parityAccumulator_reg[4]  ( .D(n8414), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/parityAccumulator[4] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/parityAccumulator_reg[5]  ( .D(n8413), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/parityAccumulator[5] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/parityAccumulator_reg[6]  ( .D(n8412), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/parityAccumulator[6] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/parityAccumulator_reg[7]  ( .D(n8411), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/parityAccumulator[7] ) );
  DFFSR \U_1/U_0/U_1/U_8/PARITY_ERROR_reg  ( .D(
        \U_1/U_0/U_1/U_8/nextParityError ), .CLK(CLK), .R(n9496), .S(1'b1), 
        .Q(PARITY_ERROR1) );
  DFFSR \U_1/U_0/U_1/U_8/parityError_reg  ( .D(
        \U_1/U_0/U_1/U_8/nextParityError ), .CLK(CLK), .R(n9496), .S(1'b1), 
        .Q(\U_1/U_0/U_1/U_8/parityError ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[0]  ( .D(n8410), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[0] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[0]  ( .D(n7270), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [0]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[1]  ( .D(n8409), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[1] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[1]  ( .D(n7269), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [1]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[2]  ( .D(n8408), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[2] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[2]  ( .D(n7268), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [2]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[3]  ( .D(n8407), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[3] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[3]  ( .D(n7267), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [3]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[4]  ( .D(n8406), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[4] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[4]  ( .D(n10422), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [4]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[5]  ( .D(n8405), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[5] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[5]  ( .D(n10423), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [5]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[6]  ( .D(n8404), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[6] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[6]  ( .D(n10424), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [6]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[7]  ( .D(n8403), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[7] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[7]  ( .D(n10425), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [7]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[8]  ( .D(n8402), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[8] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[8]  ( .D(n10426), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [8]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[9]  ( .D(n8401), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[9] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[9]  ( .D(n10427), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [9]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[10]  ( .D(n8400), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[10] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[10]  ( .D(n10428), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [10]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[11]  ( .D(n8399), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[11] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[11]  ( .D(n10429), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [11]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[12]  ( .D(n8398), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[12] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[12]  ( .D(n10430), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [12]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[13]  ( .D(n8397), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[13] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[13]  ( .D(n10431), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [13]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[14]  ( .D(n8396), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[14] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[14]  ( .D(n10432), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [14]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[15]  ( .D(n8395), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[15] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[15]  ( .D(n10433), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [15]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[16]  ( .D(n8394), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[16] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[16]  ( .D(n10434), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [16]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[17]  ( .D(n8393), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[17] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[17]  ( .D(n10435), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [17]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[18]  ( .D(n8392), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[18] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[18]  ( .D(n10436), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [18]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[19]  ( .D(n8391), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[19] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[19]  ( .D(n10437), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [19]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[20]  ( .D(n8390), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[20] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[20]  ( .D(n10438), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [20]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[21]  ( .D(n8389), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[21] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[21]  ( .D(n10439), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [21]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[22]  ( .D(n8388), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[22] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[22]  ( .D(n10440), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [22]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[23]  ( .D(n8387), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[23] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[23]  ( .D(n10441), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [23]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[24]  ( .D(n8386), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[24] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[24]  ( .D(n10442), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [24]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[25]  ( .D(n8385), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[25] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[25]  ( .D(n10443), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [25]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[26]  ( .D(n8384), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[26] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[26]  ( .D(n10444), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [26]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[27]  ( .D(n8383), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[27] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[27]  ( .D(n10445), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [27]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[28]  ( .D(n8382), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[28] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[28]  ( .D(n10446), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [28]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[29]  ( .D(n8381), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[29] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[29]  ( .D(n10447), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [29]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[30]  ( .D(n8380), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[30] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[30]  ( .D(n10448), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [30]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[31]  ( .D(n8379), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[31] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[31]  ( .D(n10449), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [31]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[32]  ( .D(n8378), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[32] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[32]  ( .D(n10450), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [32]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[33]  ( .D(n8377), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[33] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[33]  ( .D(n10451), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [33]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[34]  ( .D(n8376), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[34] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[34]  ( .D(n10452), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [34]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[35]  ( .D(n8375), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[35] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[35]  ( .D(n10453), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [35]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[36]  ( .D(n8374), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[36] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[36]  ( .D(n10454), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [36]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[37]  ( .D(n8373), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[37] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[37]  ( .D(n10455), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [37]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[38]  ( .D(n8372), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[38] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[38]  ( .D(n10456), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [38]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[39]  ( .D(n8371), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[39] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[39]  ( .D(n10457), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [39]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[40]  ( .D(n8370), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[40] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[40]  ( .D(n10458), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [40]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[41]  ( .D(n8369), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[41] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[41]  ( .D(n10459), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [41]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[42]  ( .D(n8368), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[42] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[42]  ( .D(n10460), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [42]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[43]  ( .D(n8367), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[43] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[43]  ( .D(n10461), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [43]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[44]  ( .D(n8366), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[44] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[44]  ( .D(n10462), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [44]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[45]  ( .D(n8365), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[45] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[45]  ( .D(n10463), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [45]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[46]  ( .D(n8364), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[46] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[46]  ( .D(n10464), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [46]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[47]  ( .D(n8363), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[47] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[47]  ( .D(n10465), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [47]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[48]  ( .D(n8362), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[48] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[48]  ( .D(n10466), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [48]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[49]  ( .D(n8361), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[49] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[49]  ( .D(n10467), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [49]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[50]  ( .D(n8360), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[50] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[50]  ( .D(n10468), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [50]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[51]  ( .D(n8359), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[51] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[51]  ( .D(n10469), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [51]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[52]  ( .D(n8358), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[52] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[52]  ( .D(n10470), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [52]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[53]  ( .D(n8357), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[53] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[53]  ( .D(n10471), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [53]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[54]  ( .D(n8356), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[54] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[54]  ( .D(n10472), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [54]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[55]  ( .D(n8355), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[55] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[55]  ( .D(n10473), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [55]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[56]  ( .D(n8354), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[56] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[56]  ( .D(n10474), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [56]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[57]  ( .D(n8353), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[57] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[57]  ( .D(n10475), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [57]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[58]  ( .D(n8352), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[58] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[58]  ( .D(n10476), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [58]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[59]  ( .D(n8351), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[59] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[59]  ( .D(n10477), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [59]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[60]  ( .D(n8350), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[60] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[60]  ( .D(n10478), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [60]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[61]  ( .D(n8349), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[61] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[61]  ( .D(n10479), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [61]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[62]  ( .D(n8348), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[62] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[62]  ( .D(n10480), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [62]) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/currentPlainKey_reg[63]  ( .D(n8347), .CLK(CLK), 
        .Q(\U_1/U_0/U_1/U_8/currentPlainKey[63] ) );
  DFFPOSX1 \U_1/U_0/U_1/U_8/PLAINKEY_reg[63]  ( .D(n7207), .CLK(CLK), .Q(
        \U_1/U_0/PLAINKEY [63]) );
  DFFSR \U_1/U_1/U_1/state_reg  ( .D(1'b1), .CLK(CLK), .R(n9496), .S(1'b1), 
        .Q(\U_1/U_1/U_1/state ) );
  DFFSR \U_1/U_2/U_0/DP_hold1_reg  ( .D(DPRS), .CLK(CLK), .R(1'b1), .S(n9521), 
        .Q(\U_1/U_2/U_0/DP_hold1 ) );
  DFFSR \U_1/U_2/U_0/DP_hold2_reg  ( .D(\U_1/U_2/U_0/DP_hold1 ), .CLK(CLK), 
        .R(1'b1), .S(n9522), .Q(\U_1/U_2/U_0/DP_hold2 ) );
  DFFSR \U_1/U_2/U_5/state_reg[0]  ( .D(\U_1/U_2/U_5/nextstate [0]), .CLK(CLK), 
        .R(n9496), .S(1'b1), .Q(\U_1/U_2/U_5/state[0] ) );
  DFFSR \U_1/U_2/U_5/state_reg[3]  ( .D(\U_1/U_2/U_5/nextstate [3]), .CLK(CLK), 
        .R(n9496), .S(1'b1), .Q(\U_1/U_2/U_5/state[3] ) );
  DFFSR \U_1/U_2/U_7/state_reg  ( .D(n11546), .CLK(CLK), .R(n9496), .S(1'b1), 
        .Q(\U_1/U_2/U_7/state ) );
  DFFSR \U_1/U_2/U_7/count_reg[2]  ( .D(\U_1/U_2/U_7/nextcount [2]), .CLK(CLK), 
        .R(n9496), .S(1'b1), .Q(\U_1/U_2/U_7/count[2] ) );
  DFFSR \U_1/U_2/U_7/count_reg[3]  ( .D(\U_1/U_2/U_7/nextcount [3]), .CLK(CLK), 
        .R(n9496), .S(1'b1), .Q(\U_1/U_2/U_7/count[3] ) );
  DFFSR \U_1/U_2/U_1/state_reg[0]  ( .D(\U_1/U_2/U_1/N29 ), .CLK(CLK), .R(
        n9496), .S(1'b1), .Q(\U_1/U_2/U_1/state[0] ) );
  DFFSR \U_1/U_2/U_1/DP_hold2_reg  ( .D(n8346), .CLK(CLK), .R(1'b1), .S(n9522), 
        .Q(\U_1/U_2/U_1/DP_hold2 ) );
  DFFSR \U_1/U_2/U_1/state_reg[3]  ( .D(\U_1/U_2/U_1/N32 ), .CLK(CLK), .R(
        n9496), .S(1'b1), .Q(\U_1/U_2/U_1/state[3] ) );
  DFFSR \U_1/U_2/U_1/state_reg[2]  ( .D(\U_1/U_2/U_1/N31 ), .CLK(CLK), .R(
        n9496), .S(1'b1), .Q(\U_1/U_2/U_1/state[2] ) );
  DFFSR \U_1/U_2/U_1/state_reg[1]  ( .D(n9695), .CLK(CLK), .R(n9496), .S(1'b1), 
        .Q(\U_1/U_2/U_1/state[1] ) );
  DFFSR \U_1/U_2/U_1/DP_hold1_reg  ( .D(n8345), .CLK(CLK), .R(1'b1), .S(n9522), 
        .Q(\U_1/U_2/U_1/DP_hold1 ) );
  DFFSR \U_1/U_2/U_6/present_val_reg[7]  ( .D(n8344), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/RCV_DATA [7]) );
  DFFSR \U_1/U_2/U_6/present_val_reg[6]  ( .D(n8343), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/RCV_DATA [6]) );
  DFFSR \U_1/U_2/U_6/present_val_reg[5]  ( .D(n8342), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/RCV_DATA [5]) );
  DFFSR \U_1/U_2/U_6/present_val_reg[4]  ( .D(n8341), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/RCV_DATA [4]) );
  DFFSR \U_1/U_2/U_6/present_val_reg[3]  ( .D(n8340), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/RCV_DATA [3]) );
  DFFSR \U_1/U_2/U_6/present_val_reg[2]  ( .D(n8339), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/RCV_DATA [2]) );
  DFFSR \U_1/U_2/U_6/present_val_reg[1]  ( .D(n8338), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/RCV_DATA [1]) );
  DFFSR \U_1/U_2/U_6/present_val_reg[0]  ( .D(n8337), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/RCV_DATA [0]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[7]  ( .D(n8276), .CLK(CLK), .R(
        n9497), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [7]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[15]  ( .D(n8268), .CLK(CLK), .R(
        n9497), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [15]) );
  DFFSR \U_1/U_2/U_5/state_reg[2]  ( .D(\U_1/U_2/U_5/nextstate [2]), .CLK(CLK), 
        .R(n9497), .S(1'b1), .Q(\U_1/U_2/U_5/state[2] ) );
  DFFSR \U_1/U_2/U_5/count_reg[0]  ( .D(n8330), .CLK(CLK), .R(n9497), .S(1'b1), 
        .Q(\U_1/U_2/U_5/count[0] ) );
  DFFSR \U_1/U_2/U_5/count_reg[1]  ( .D(n8331), .CLK(CLK), .R(n9498), .S(1'b1), 
        .Q(\U_1/U_2/U_5/count[1] ) );
  DFFSR \U_1/U_2/U_5/count_reg[2]  ( .D(n8332), .CLK(CLK), .R(n9498), .S(1'b1), 
        .Q(\U_1/U_2/U_5/count[2] ) );
  DFFSR \U_1/U_2/U_5/count_reg[3]  ( .D(n8333), .CLK(CLK), .R(n9498), .S(1'b1), 
        .Q(\U_1/U_2/U_5/count[3] ) );
  DFFSR \U_1/U_2/U_5/state_reg[1]  ( .D(\U_1/U_2/U_5/nextstate [1]), .CLK(CLK), 
        .R(n9498), .S(1'b1), .Q(\U_1/U_2/U_5/state[1] ) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[15]  ( .D(n8336), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[15] ) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[0]  ( .D(n8328), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[0] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[0]  ( .D(n8327), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [0]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[0]  ( .D(n8326), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [0]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[8]  ( .D(n8304), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[8] ) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[2]  ( .D(n8322), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[2] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[2]  ( .D(n8321), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [2]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[2]  ( .D(n8320), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [2]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[10]  ( .D(n8298), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[10] ) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[3]  ( .D(n8319), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[3] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[3]  ( .D(n8318), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [3]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[3]  ( .D(n8317), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [3]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[11]  ( .D(n8295), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[11] ) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[4]  ( .D(n8316), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[4] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[4]  ( .D(n8315), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [4]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[4]  ( .D(n8314), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [4]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[12]  ( .D(n8292), .CLK(CLK), .R(n9491), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[12] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[12]  ( .D(n8291), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [12]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[12]  ( .D(n8290), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [12]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[5]  ( .D(n8313), .CLK(CLK), .R(n9492), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[5] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[5]  ( .D(n8312), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [5]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[5]  ( .D(n8311), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [5]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[13]  ( .D(n8289), .CLK(CLK), .R(n9493), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[13] ) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[6]  ( .D(n8310), .CLK(CLK), .R(n9495), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[6] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[6]  ( .D(n8309), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [6]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[6]  ( .D(n8308), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [6]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[14]  ( .D(n8286), .CLK(CLK), .R(n9494), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[14] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[14]  ( .D(n8285), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [14]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[14]  ( .D(n8284), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [14]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[7]  ( .D(n8307), .CLK(CLK), .R(n9496), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[7] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[7]  ( .D(n8306), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [7]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[7]  ( .D(n8305), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [7]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[13]  ( .D(n8288), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [13]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[13]  ( .D(n8287), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [13]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[11]  ( .D(n8294), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [11]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[11]  ( .D(n8293), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [11]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[1]  ( .D(n8325), .CLK(CLK), .R(n9495), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[1] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[1]  ( .D(n8324), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [1]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[1]  ( .D(n8323), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [1]) );
  DFFSR \U_1/U_2/U_2/current_crc_reg[9]  ( .D(n8301), .CLK(CLK), .R(n9490), 
        .S(1'b1), .Q(\U_1/U_2/U_2/current_crc[9] ) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[9]  ( .D(n8300), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [9]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[9]  ( .D(n8299), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [9]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[10]  ( .D(n8297), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [10]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[10]  ( .D(n8296), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [10]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[8]  ( .D(n8303), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [8]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[8]  ( .D(n8302), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [8]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_1_reg[15]  ( .D(n8335), .CLK(CLK), .Q(
        \U_1/U_2/U_2/cache_1 [15]) );
  DFFPOSX1 \U_1/U_2/U_2/cache_2_reg[15]  ( .D(n8334), .CLK(CLK), .Q(
        \U_1/U_2/RX_CRC [15]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[0]  ( .D(n8283), .CLK(CLK), .R(
        n9517), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [0]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[8]  ( .D(n8275), .CLK(CLK), .R(
        n9497), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [8]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[1]  ( .D(n8282), .CLK(CLK), .R(
        n9498), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [1]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[9]  ( .D(n8274), .CLK(CLK), .R(
        n9499), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [9]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[2]  ( .D(n8281), .CLK(CLK), .R(
        n9499), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [2]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[10]  ( .D(n8273), .CLK(CLK), .R(
        n9499), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [10]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[3]  ( .D(n8280), .CLK(CLK), .R(
        n9499), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [3]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[11]  ( .D(n8272), .CLK(CLK), .R(
        n9499), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [11]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[4]  ( .D(n8279), .CLK(CLK), .R(
        n9521), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [4]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[12]  ( .D(n8271), .CLK(CLK), .R(
        n9520), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [12]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[5]  ( .D(n8278), .CLK(CLK), .R(
        n9521), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [5]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[13]  ( .D(n8270), .CLK(CLK), .R(
        n9520), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [13]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[6]  ( .D(n8277), .CLK(CLK), .R(
        n9520), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [6]) );
  DFFSR \U_1/U_2/U_3/present_CHECK_CRC_reg[14]  ( .D(n8269), .CLK(CLK), .R(
        n9520), .S(1'b1), .Q(\U_1/U_2/rx_CHECK_CRC [14]) );
  DFFSR \U_1/U_2/U_7/count_reg[0]  ( .D(\U_1/U_2/U_7/nextcount [0]), .CLK(CLK), 
        .R(n9520), .S(1'b1), .Q(\U_1/U_2/U_7/count[0] ) );
  DFFSR \U_1/U_2/U_7/count_reg[1]  ( .D(\U_1/U_2/U_7/nextcount [1]), .CLK(CLK), 
        .R(n9520), .S(1'b1), .Q(\U_1/U_2/U_7/count[1] ) );
  DFFPOSX1 \U_1/U_2/U_5/curR_ERROR_reg  ( .D(n8329), .CLK(CLK), .Q(
        \U_1/U_2/U_5/curR_ERROR ) );
  DFFSR \U_1/U_2/U_5/R_ERROR_reg  ( .D(n9696), .CLK(CLK), .R(n9520), .S(1'b1), 
        .Q(RE_S) );
  DFFPOSX1 \U_1/U_2/U_5/curCRC_ERROR_reg  ( .D(n8267), .CLK(CLK), .Q(
        \U_1/U_2/U_5/curCRC_ERROR ) );
  DFFPOSX1 \U_1/U_2/U_5/CRC_ERROR_reg  ( .D(n8266), .CLK(CLK), .Q(CRCE_S) );
  DFFSR \U_1/U_3/U_0/dp_tx_out_reg  ( .D(\U_1/U_3/U_0/DE_holdout_nxt ), .CLK(
        CLK), .R(1'b1), .S(n9522), .Q(DPTH) );
  DFFSR \U_1/U_3/U_0/state_reg[3]  ( .D(\U_1/U_3/U_0/nextstate [3]), .CLK(CLK), 
        .R(n9520), .S(1'b1), .Q(\U_1/U_3/U_0/state[3] ) );
  DFFSR \U_1/U_3/U_0/DE_holdout_reg  ( .D(\U_1/U_3/U_0/DE_holdout_nxt ), .CLK(
        CLK), .R(1'b1), .S(n9522), .Q(\U_1/U_3/U_0/DE_holdout ) );
  DFFPOSX1 \U_1/U_3/U_0/DE_holdout_last_reg  ( .D(n7140), .CLK(CLK), .Q(
        \U_1/U_3/U_0/DE_holdout_last ) );
  DFFSR \U_1/U_3/U_4/SHIFT_ENABLE_E_reg  ( .D(n7756), .CLK(CLK), .R(n9520), 
        .S(1'b1), .Q(\U_1/U_3/SHIFT_ENABLE_E ) );
  DFFSR \U_1/U_3/U_0/state_reg[2]  ( .D(\U_1/U_3/U_0/nextstate [2]), .CLK(CLK), 
        .R(n9520), .S(1'b1), .Q(\U_1/U_3/U_0/state[2] ) );
  DFFSR \U_1/U_3/U_0/state_reg[0]  ( .D(\U_1/U_3/U_0/nextstate [0]), .CLK(CLK), 
        .R(n9520), .S(1'b1), .Q(\U_1/U_3/U_0/state[0] ) );
  DFFSR \U_1/U_3/U_0/state_reg[1]  ( .D(\U_1/U_3/U_0/nextstate [1]), .CLK(CLK), 
        .R(n9519), .S(1'b1), .Q(\U_1/U_3/U_0/state[1] ) );
  DFFSR \U_1/U_3/U_3/count_reg[6]  ( .D(n7792), .CLK(CLK), .R(n9520), .S(1'b1), 
        .Q(\U_1/U_3/U_3/N188 ) );
  DFFSR \U_1/U_3/U_3/state_reg[1]  ( .D(\U_1/U_3/U_3/nextstate [1]), .CLK(CLK), 
        .R(n9519), .S(1'b1), .Q(\U_1/U_3/U_3/state[1] ) );
  DFFSR \U_1/U_3/U_3/state_reg[2]  ( .D(\U_1/U_3/U_3/nextstate [2]), .CLK(CLK), 
        .R(n9519), .S(1'b1), .Q(\U_1/U_3/U_3/state[2] ) );
  DFFSR \U_1/U_3/U_3/state_reg[0]  ( .D(\U_1/U_3/U_3/nextstate [0]), .CLK(CLK), 
        .R(n9519), .S(1'b1), .Q(\U_1/U_3/U_3/state[0] ) );
  DFFSR \U_1/U_1/U_0/state_reg[2]  ( .D(\U_1/U_1/U_0/nextState [2]), .CLK(CLK), 
        .R(n9519), .S(1'b1), .Q(\U_1/U_1/U_0/state[2] ) );
  DFFPOSX1 \U_1/U_1/U_0/R_ENABLE_reg  ( .D(n7130), .CLK(CLK), .Q(
        \U_1/U_1/R_ENABLE ) );
  DFFSR \U_1/U_1/U_1/readptr_reg[0]  ( .D(\U_1/U_1/U_1/N343 ), .CLK(CLK), .R(
        n9519), .S(1'b1), .Q(\U_1/U_1/U_1/readptr[0] ) );
  DFFSR \U_1/U_1/U_1/readptr_reg[1]  ( .D(\U_1/U_1/U_1/N344 ), .CLK(CLK), .R(
        n9519), .S(1'b1), .Q(\U_1/U_1/U_1/readptr[1] ) );
  DFFSR \U_1/U_1/U_1/readptr_reg[2]  ( .D(\U_1/U_1/U_1/N345 ), .CLK(CLK), .R(
        n9519), .S(1'b1), .Q(\U_1/U_1/U_1/readptr[2] ) );
  DFFSR \U_1/U_1/U_1/readptr_reg[3]  ( .D(\U_1/U_1/U_1/N346 ), .CLK(CLK), .R(
        n9519), .S(1'b1), .Q(\U_1/U_1/U_1/readptr[3] ) );
  DFFSR \U_1/U_1/U_1/readptr_reg[4]  ( .D(\U_1/U_1/U_1/N347 ), .CLK(CLK), .R(
        n9518), .S(1'b1), .Q(\U_1/U_1/U_1/readptr[4] ) );
  DFFSR \U_1/U_1/U_1/writeptr_reg[4]  ( .D(n8264), .CLK(CLK), .R(n9519), .S(
        1'b1), .Q(\U_1/U_1/U_1/writeptr[4] ) );
  DFFSR \U_1/U_1/U_1/writeptr_reg[3]  ( .D(n8260), .CLK(CLK), .R(n9519), .S(
        1'b1), .Q(\U_1/U_1/U_1/writeptr[3] ) );
  DFFSR \U_1/U_1/U_1/writeptr_reg[0]  ( .D(n8263), .CLK(CLK), .R(n9519), .S(
        1'b1), .Q(\U_1/U_1/U_1/writeptr[0] ) );
  DFFSR \U_1/U_1/U_1/writeptr_reg[1]  ( .D(n8262), .CLK(CLK), .R(n9518), .S(
        1'b1), .Q(\U_1/U_1/U_1/writeptr[1] ) );
  DFFSR \U_1/U_1/U_1/writeptr_reg[2]  ( .D(n8261), .CLK(CLK), .R(n9518), .S(
        1'b1), .Q(\U_1/U_1/U_1/writeptr[2] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[0][0]  ( .D(n10072), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[0][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[0][1]  ( .D(n10071), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[0][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[0][0]  ( .D(n10279), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[0][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[0][1]  ( .D(n10278), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[0][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[0][2]  ( .D(n10277), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[0][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[0][3]  ( .D(n10276), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[0][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[0][4]  ( .D(n10275), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[0][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[0][5]  ( .D(n10274), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[0][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[0][6]  ( .D(n10273), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[0][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[0][7]  ( .D(n10272), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[0][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[1][0]  ( .D(n10069), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[1][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[1][1]  ( .D(n10068), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[1][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[1][0]  ( .D(n10270), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[1][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[1][1]  ( .D(n10269), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[1][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[1][2]  ( .D(n10268), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[1][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[1][3]  ( .D(n10267), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[1][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[1][4]  ( .D(n10266), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[1][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[1][5]  ( .D(n10265), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[1][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[1][6]  ( .D(n10264), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[1][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[1][7]  ( .D(n10263), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[1][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[2][0]  ( .D(n10066), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[2][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[2][1]  ( .D(n10065), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[2][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[2][0]  ( .D(n10261), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[2][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[2][1]  ( .D(n10260), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[2][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[2][2]  ( .D(n10259), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[2][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[2][3]  ( .D(n10258), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[2][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[2][4]  ( .D(n10257), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[2][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[2][5]  ( .D(n10256), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[2][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[2][6]  ( .D(n10255), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[2][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[2][7]  ( .D(n10254), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[2][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[3][0]  ( .D(n10063), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[3][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[3][1]  ( .D(n10062), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[3][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[3][0]  ( .D(n10252), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[3][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[3][1]  ( .D(n10251), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[3][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[3][2]  ( .D(n10250), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[3][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[3][3]  ( .D(n10249), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[3][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[3][4]  ( .D(n10248), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[3][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[3][5]  ( .D(n10247), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[3][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[3][6]  ( .D(n10246), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[3][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[3][7]  ( .D(n10245), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[3][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[4][0]  ( .D(n8205), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[4][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[4][1]  ( .D(n8204), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[4][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[4][0]  ( .D(n7979), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[4][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[4][1]  ( .D(n7978), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[4][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[4][2]  ( .D(n7977), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[4][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[4][3]  ( .D(n7976), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[4][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[4][4]  ( .D(n7975), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[4][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[4][5]  ( .D(n7974), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[4][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[4][6]  ( .D(n7973), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[4][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[4][7]  ( .D(n7972), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[4][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[5][0]  ( .D(n8207), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[5][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[5][1]  ( .D(n8206), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[5][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[5][0]  ( .D(n7987), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[5][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[5][1]  ( .D(n7986), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[5][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[5][2]  ( .D(n7985), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[5][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[5][3]  ( .D(n7984), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[5][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[5][4]  ( .D(n7983), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[5][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[5][5]  ( .D(n7982), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[5][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[5][6]  ( .D(n7981), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[5][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[5][7]  ( .D(n7980), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[5][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[6][0]  ( .D(n7995), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[6][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[6][1]  ( .D(n7994), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[6][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[6][2]  ( .D(n7993), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[6][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[6][3]  ( .D(n7992), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[6][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[6][4]  ( .D(n7991), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[6][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[6][5]  ( .D(n7990), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[6][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[6][6]  ( .D(n7989), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[6][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[6][7]  ( .D(n7988), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[6][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[7][6]  ( .D(n8003), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[7][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[7][7]  ( .D(n8002), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[7][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[7][0]  ( .D(n8001), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[7][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[7][1]  ( .D(n8000), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[7][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[7][2]  ( .D(n7999), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[7][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[7][3]  ( .D(n7998), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[7][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[7][4]  ( .D(n7997), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[7][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[7][5]  ( .D(n7996), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[7][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[11][1]  ( .D(n8219), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[11][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[11][0]  ( .D(n8218), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[11][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[6][0]  ( .D(n8209), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[6][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[6][1]  ( .D(n8208), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[6][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[7][0]  ( .D(n8211), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[7][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[7][1]  ( .D(n8210), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[7][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[11][0]  ( .D(n8035), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[11][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[11][1]  ( .D(n8034), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[11][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[11][2]  ( .D(n8033), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[11][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[11][3]  ( .D(n8032), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[11][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[11][4]  ( .D(n8031), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[11][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[11][5]  ( .D(n8030), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[11][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[11][6]  ( .D(n8029), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[11][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[11][7]  ( .D(n8028), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[11][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[8][0]  ( .D(n8213), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[8][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[8][1]  ( .D(n8212), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[8][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[8][0]  ( .D(n8011), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[8][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[8][1]  ( .D(n8010), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[8][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[8][2]  ( .D(n8009), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[8][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[8][3]  ( .D(n8008), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[8][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[8][4]  ( .D(n8007), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[8][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[8][5]  ( .D(n8006), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[8][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[8][6]  ( .D(n8005), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[8][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[8][7]  ( .D(n8004), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[8][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[9][0]  ( .D(n8215), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[9][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[9][1]  ( .D(n8214), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[9][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[9][0]  ( .D(n8019), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[9][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[9][1]  ( .D(n8018), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[9][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[9][2]  ( .D(n8017), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[9][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[9][3]  ( .D(n8016), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[9][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[9][4]  ( .D(n8015), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[9][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[9][5]  ( .D(n8014), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[9][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[9][6]  ( .D(n8013), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[9][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[9][7]  ( .D(n8012), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[9][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[10][0]  ( .D(n8217), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[10][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[10][1]  ( .D(n8216), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[10][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[10][0]  ( .D(n8027), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[10][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[10][1]  ( .D(n8026), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[10][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[10][2]  ( .D(n8025), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[10][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[10][3]  ( .D(n8024), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[10][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[10][4]  ( .D(n8023), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[10][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[10][5]  ( .D(n8022), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[10][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[10][6]  ( .D(n8021), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[10][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[10][7]  ( .D(n8020), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[10][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[12][0]  ( .D(n10114), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[12][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[12][1]  ( .D(n10113), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[12][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[12][0]  ( .D(n10235), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[12][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[12][1]  ( .D(n10234), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[12][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[12][2]  ( .D(n10233), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[12][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[12][3]  ( .D(n10232), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[12][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[12][4]  ( .D(n10231), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[12][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[12][5]  ( .D(n10230), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[12][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[12][6]  ( .D(n10229), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[12][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[12][7]  ( .D(n10228), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[12][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[13][0]  ( .D(n10111), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[13][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[13][1]  ( .D(n10110), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[13][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[13][0]  ( .D(n10226), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[13][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[13][1]  ( .D(n10225), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[13][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[13][2]  ( .D(n10224), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[13][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[13][3]  ( .D(n10223), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[13][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[13][4]  ( .D(n10222), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[13][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[13][5]  ( .D(n10221), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[13][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[13][6]  ( .D(n10220), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[13][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[13][7]  ( .D(n10219), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[13][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[14][0]  ( .D(n10217), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[14][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[14][1]  ( .D(n10216), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[14][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[14][2]  ( .D(n10215), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[14][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[14][3]  ( .D(n10214), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[14][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[14][4]  ( .D(n10213), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[14][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[14][5]  ( .D(n10212), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[14][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[14][6]  ( .D(n10211), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[14][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[14][7]  ( .D(n10210), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[14][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[15][0]  ( .D(n10208), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[15][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[15][1]  ( .D(n10207), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[15][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[15][2]  ( .D(n10206), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[15][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[15][3]  ( .D(n10205), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[15][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[15][4]  ( .D(n10204), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[15][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[15][5]  ( .D(n10203), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[15][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[15][6]  ( .D(n10202), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[15][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[15][7]  ( .D(n10201), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[15][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[24][0]  ( .D(n10086), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[24][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[24][1]  ( .D(n10085), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[24][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[24][0]  ( .D(n10159), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[24][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[24][1]  ( .D(n10158), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[24][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[24][2]  ( .D(n10157), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[24][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[24][3]  ( .D(n10156), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[24][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[24][4]  ( .D(n10155), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[24][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[24][5]  ( .D(n10154), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[24][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[24][6]  ( .D(n10153), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[24][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[24][7]  ( .D(n10152), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[24][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[25][0]  ( .D(n10083), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[25][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[25][1]  ( .D(n10082), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[25][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[25][0]  ( .D(n10150), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[25][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[25][1]  ( .D(n10149), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[25][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[25][2]  ( .D(n10148), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[25][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[25][3]  ( .D(n10147), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[25][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[25][4]  ( .D(n10146), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[25][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[25][5]  ( .D(n10145), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[25][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[25][6]  ( .D(n10144), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[25][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[25][7]  ( .D(n10143), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[25][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[26][0]  ( .D(n10080), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[26][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[26][1]  ( .D(n10079), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[26][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[26][0]  ( .D(n10141), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[26][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[26][1]  ( .D(n10140), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[26][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[26][2]  ( .D(n10139), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[26][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[26][3]  ( .D(n10138), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[26][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[26][4]  ( .D(n10137), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[26][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[26][5]  ( .D(n10136), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[26][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[26][6]  ( .D(n10135), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[26][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[26][7]  ( .D(n10134), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[26][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[27][0]  ( .D(n10077), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[27][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[27][1]  ( .D(n10076), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[27][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[27][0]  ( .D(n10132), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[27][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[27][1]  ( .D(n10131), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[27][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[27][2]  ( .D(n10130), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[27][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[27][3]  ( .D(n10129), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[27][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[27][4]  ( .D(n10128), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[27][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[27][5]  ( .D(n10127), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[27][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[27][6]  ( .D(n10126), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[27][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[27][7]  ( .D(n10125), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[27][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[28][0]  ( .D(n8253), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[28][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[28][1]  ( .D(n8252), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[28][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[28][0]  ( .D(n8171), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[28][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[28][1]  ( .D(n8170), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[28][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[28][2]  ( .D(n8169), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[28][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[28][3]  ( .D(n8168), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[28][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[28][4]  ( .D(n8167), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[28][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[28][5]  ( .D(n8166), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[28][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[28][6]  ( .D(n8165), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[28][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[28][7]  ( .D(n8164), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[28][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[29][0]  ( .D(n8255), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[29][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[29][1]  ( .D(n8254), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[29][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[29][0]  ( .D(n8179), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[29][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[29][1]  ( .D(n8178), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[29][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[29][2]  ( .D(n8177), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[29][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[29][3]  ( .D(n8176), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[29][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[29][4]  ( .D(n8175), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[29][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[29][5]  ( .D(n8174), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[29][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[29][6]  ( .D(n8173), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[29][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[29][7]  ( .D(n8172), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[29][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[30][0]  ( .D(n8257), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[30][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[30][1]  ( .D(n8256), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[30][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[30][0]  ( .D(n8187), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[30][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[30][1]  ( .D(n8186), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[30][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[30][2]  ( .D(n8185), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[30][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[30][3]  ( .D(n8184), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[30][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[30][4]  ( .D(n8183), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[30][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[30][5]  ( .D(n8182), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[30][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[30][6]  ( .D(n8181), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[30][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[30][7]  ( .D(n8180), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[30][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[31][0]  ( .D(n8259), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[31][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[31][1]  ( .D(n8258), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[31][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[31][0]  ( .D(n8195), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[31][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[31][1]  ( .D(n8194), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[31][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[31][2]  ( .D(n8193), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[31][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[31][3]  ( .D(n8192), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[31][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[31][4]  ( .D(n8191), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[31][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[31][5]  ( .D(n8190), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[31][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[31][6]  ( .D(n8189), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[31][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[31][7]  ( .D(n8188), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[31][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[14][0]  ( .D(n10108), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[14][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[14][1]  ( .D(n10107), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[14][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[15][0]  ( .D(n10105), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[15][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[15][1]  ( .D(n10104), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[15][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[16][0]  ( .D(n8229), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[16][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[16][1]  ( .D(n8228), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[16][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[16][0]  ( .D(n8075), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[16][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[16][1]  ( .D(n8074), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[16][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[16][2]  ( .D(n8073), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[16][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[16][3]  ( .D(n8072), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[16][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[16][4]  ( .D(n8071), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[16][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[16][5]  ( .D(n8070), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[16][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[16][6]  ( .D(n8069), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[16][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[16][7]  ( .D(n8068), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[16][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[17][0]  ( .D(n8231), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[17][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[17][1]  ( .D(n8230), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[17][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[17][0]  ( .D(n8083), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[17][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[17][1]  ( .D(n8082), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[17][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[17][2]  ( .D(n8081), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[17][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[17][3]  ( .D(n8080), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[17][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[17][4]  ( .D(n8079), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[17][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[17][5]  ( .D(n8078), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[17][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[17][6]  ( .D(n8077), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[17][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[17][7]  ( .D(n8076), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[17][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[18][0]  ( .D(n8233), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[18][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[18][1]  ( .D(n8232), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[18][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[18][0]  ( .D(n8091), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[18][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[18][1]  ( .D(n8090), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[18][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[18][2]  ( .D(n8089), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[18][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[18][3]  ( .D(n8088), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[18][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[18][4]  ( .D(n8087), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[18][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[18][5]  ( .D(n8086), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[18][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[18][6]  ( .D(n8085), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[18][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[18][7]  ( .D(n8084), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[18][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[19][0]  ( .D(n8235), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[19][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[19][1]  ( .D(n8234), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[19][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[19][3]  ( .D(n8099), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[19][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[19][4]  ( .D(n8098), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[19][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[19][5]  ( .D(n8097), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[19][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[19][6]  ( .D(n8096), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[19][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[19][7]  ( .D(n8095), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[19][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[19][0]  ( .D(n8094), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[19][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[19][1]  ( .D(n8093), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[19][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[19][2]  ( .D(n8092), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[19][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[20][0]  ( .D(n10098), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[20][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[20][1]  ( .D(n10097), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[20][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[20][0]  ( .D(n10195), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[20][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[20][1]  ( .D(n10194), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[20][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[20][2]  ( .D(n10193), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[20][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[20][3]  ( .D(n10192), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[20][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[20][4]  ( .D(n10191), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[20][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[20][5]  ( .D(n10190), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[20][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[20][6]  ( .D(n10189), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[20][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[20][7]  ( .D(n10188), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[20][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[21][0]  ( .D(n10095), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[21][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[21][1]  ( .D(n10094), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[21][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[21][0]  ( .D(n10186), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[21][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[21][1]  ( .D(n10185), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[21][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[21][2]  ( .D(n10184), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[21][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[21][3]  ( .D(n10183), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[21][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[21][4]  ( .D(n10182), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[21][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[21][5]  ( .D(n10181), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[21][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[21][6]  ( .D(n10180), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[21][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[21][7]  ( .D(n10179), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[21][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[22][0]  ( .D(n10092), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[22][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[22][1]  ( .D(n10091), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[22][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[22][0]  ( .D(n10177), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[22][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[22][1]  ( .D(n10176), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[22][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[22][2]  ( .D(n10175), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[22][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[22][3]  ( .D(n10174), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[22][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[22][4]  ( .D(n10173), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[22][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[22][5]  ( .D(n10172), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[22][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[22][6]  ( .D(n10171), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[22][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[22][7]  ( .D(n10170), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[22][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[23][0]  ( .D(n10089), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[23][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/opcode_reg[23][1]  ( .D(n10088), .CLK(CLK), .Q(
        \U_1/U_1/U_1/opcode[23][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[23][0]  ( .D(n10168), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[23][0] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[23][1]  ( .D(n10167), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[23][1] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[23][2]  ( .D(n10166), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[23][2] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[23][3]  ( .D(n10165), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[23][3] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[23][4]  ( .D(n10164), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[23][4] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[23][5]  ( .D(n10163), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[23][5] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[23][6]  ( .D(n10162), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[23][6] ) );
  DFFPOSX1 \U_1/U_1/U_1/memory_reg[23][7]  ( .D(n10161), .CLK(CLK), .Q(
        \U_1/U_1/U_1/memory[23][7] ) );
  DFFPOSX1 \U_1/U_1/U_1/FULL_reg  ( .D(n10481), .CLK(CLK), .Q(FULL_S) );
  DFFPOSX1 \U_1/U_1/U_1/EMPTY_reg  ( .D(n10482), .CLK(CLK), .Q(EMPTY_S) );
  DFFSR \U_1/U_1/U_1/BYTE_COUNT_reg[0]  ( .D(\U_1/U_1/U_1/N338 ), .CLK(CLK), 
        .R(n9518), .S(1'b1), .Q(\U_1/U_1/BYTE_COUNT [0]) );
  DFFSR \U_1/U_1/U_1/BYTE_COUNT_reg[1]  ( .D(\U_1/U_1/U_1/N339 ), .CLK(CLK), 
        .R(n9518), .S(1'b1), .Q(\U_1/U_1/BYTE_COUNT [1]) );
  DFFSR \U_1/U_1/U_1/BYTE_COUNT_reg[2]  ( .D(\U_1/U_1/U_1/N340 ), .CLK(CLK), 
        .R(n9518), .S(1'b1), .Q(\U_1/U_1/BYTE_COUNT [2]) );
  DFFSR \U_1/U_1/U_1/BYTE_COUNT_reg[3]  ( .D(\U_1/U_1/U_1/N341 ), .CLK(CLK), 
        .R(n9518), .S(1'b1), .Q(\U_1/U_1/BYTE_COUNT [3]) );
  DFFSR \U_1/U_1/U_1/BYTE_COUNT_reg[4]  ( .D(\U_1/U_1/U_1/N342 ), .CLK(CLK), 
        .R(n9518), .S(1'b1), .Q(\U_1/U_1/U_0/N39 ) );
  DFFPOSX1 \U_1/U_1/U_1/DATA_reg[0]  ( .D(n7939), .CLK(CLK), .Q(
        \U_1/U_1/DATA [0]) );
  DFFPOSX1 \U_1/U_1/U_1/DATA_reg[1]  ( .D(n7938), .CLK(CLK), .Q(
        \U_1/U_1/DATA [1]) );
  DFFPOSX1 \U_1/U_1/U_1/DATA_reg[2]  ( .D(n7937), .CLK(CLK), .Q(
        \U_1/U_1/DATA [2]) );
  DFFPOSX1 \U_1/U_1/U_1/DATA_reg[3]  ( .D(n7936), .CLK(CLK), .Q(
        \U_1/U_1/DATA [3]) );
  DFFPOSX1 \U_1/U_1/U_1/DATA_reg[4]  ( .D(n7935), .CLK(CLK), .Q(
        \U_1/U_1/DATA [4]) );
  DFFPOSX1 \U_1/U_1/U_1/DATA_reg[5]  ( .D(n7934), .CLK(CLK), .Q(
        \U_1/U_1/DATA [5]) );
  DFFPOSX1 \U_1/U_1/U_1/DATA_reg[6]  ( .D(n7933), .CLK(CLK), .Q(
        \U_1/U_1/DATA [6]) );
  DFFPOSX1 \U_1/U_1/U_1/DATA_reg[7]  ( .D(n7932), .CLK(CLK), .Q(
        \U_1/U_1/DATA [7]) );
  DFFPOSX1 \U_1/U_1/U_1/OUT_OPCODE_reg[0]  ( .D(n7931), .CLK(CLK), .Q(
        \U_1/U_1/OUT_OPCODE [0]) );
  DFFPOSX1 \U_1/U_1/U_1/OUT_OPCODE_reg[1]  ( .D(n7930), .CLK(CLK), .Q(
        \U_1/U_1/OUT_OPCODE [1]) );
  DFFSR \U_1/U_1/U_0/state_reg[0]  ( .D(\U_1/U_1/U_0/nextState [0]), .CLK(CLK), 
        .R(n9518), .S(1'b1), .Q(\U_1/U_1/U_0/state[0] ) );
  DFFSR \U_1/U_1/U_0/state_reg[1]  ( .D(\U_1/U_1/U_0/nextState [1]), .CLK(CLK), 
        .R(n9518), .S(1'b1), .Q(\U_1/U_1/U_0/state[1] ) );
  DFFPOSX1 \U_1/U_1/U_0/B_READY_reg  ( .D(n7110), .CLK(CLK), .Q(\U_1/B_READY )
         );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_OPCODE_reg[0]  ( .D(n7109), .CLK(CLK), .Q(
        \U_1/PRGA_OPCODE[0] ) );
  DFFPOSX1 \U_1/U_1/U_0/tempOpcode_reg[0]  ( .D(n7108), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempOpcode [0]) );
  DFFPOSX1 \U_1/U_1/U_0/tempData_reg[7]  ( .D(n7107), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempData [7]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_IN_reg[7]  ( .D(n7106), .CLK(CLK), .Q(
        \U_1/PRGA_IN [7]) );
  DFFPOSX1 \U_1/U_1/U_0/tempData_reg[6]  ( .D(n7105), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempData [6]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_IN_reg[6]  ( .D(n7104), .CLK(CLK), .Q(
        \U_1/PRGA_IN [6]) );
  DFFPOSX1 \U_1/U_1/U_0/tempData_reg[5]  ( .D(n7103), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempData [5]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_IN_reg[5]  ( .D(n7102), .CLK(CLK), .Q(
        \U_1/PRGA_IN [5]) );
  DFFPOSX1 \U_1/U_1/U_0/tempData_reg[4]  ( .D(n7101), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempData [4]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_IN_reg[4]  ( .D(n7100), .CLK(CLK), .Q(
        \U_1/PRGA_IN [4]) );
  DFFPOSX1 \U_1/U_1/U_0/tempData_reg[3]  ( .D(n7099), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempData [3]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_IN_reg[3]  ( .D(n7098), .CLK(CLK), .Q(
        \U_1/PRGA_IN [3]) );
  DFFPOSX1 \U_1/U_1/U_0/tempData_reg[2]  ( .D(n7097), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempData [2]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_IN_reg[2]  ( .D(n7096), .CLK(CLK), .Q(
        \U_1/PRGA_IN [2]) );
  DFFPOSX1 \U_1/U_1/U_0/tempData_reg[1]  ( .D(n7095), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempData [1]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_IN_reg[1]  ( .D(n7094), .CLK(CLK), .Q(
        \U_1/PRGA_IN [1]) );
  DFFPOSX1 \U_1/U_1/U_0/tempData_reg[0]  ( .D(n7093), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempData [0]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_IN_reg[0]  ( .D(n7092), .CLK(CLK), .Q(
        \U_1/PRGA_IN [0]) );
  DFFPOSX1 \U_1/U_1/U_0/PRGA_OPCODE_reg[1]  ( .D(n7091), .CLK(CLK), .Q(
        \U_1/PRGA_OPCODE[1] ) );
  DFFSR \U_1/U_3/U_3/count_reg[0]  ( .D(n8265), .CLK(CLK), .R(n9518), .S(1'b1), 
        .Q(\U_1/U_3/U_3/count[0] ) );
  DFFSR \U_1/U_3/U_3/count_reg[5]  ( .D(n7793), .CLK(CLK), .R(n9518), .S(1'b1), 
        .Q(\U_1/U_3/U_3/count[5] ) );
  DFFSR \U_1/U_3/U_3/count_reg[1]  ( .D(n7797), .CLK(CLK), .R(n9517), .S(1'b1), 
        .Q(\U_1/U_3/U_3/count[1] ) );
  DFFSR \U_1/U_3/U_3/count_reg[2]  ( .D(n7796), .CLK(CLK), .R(n9517), .S(1'b1), 
        .Q(\U_1/U_3/U_3/count[2] ) );
  DFFSR \U_1/U_3/U_3/count_reg[3]  ( .D(n7795), .CLK(CLK), .R(n9517), .S(1'b1), 
        .Q(\U_1/U_3/U_3/count[3] ) );
  DFFSR \U_1/U_3/U_3/count_reg[4]  ( .D(n7794), .CLK(CLK), .R(n9517), .S(1'b1), 
        .Q(\U_1/U_3/U_3/count[4] ) );
  DFFSR \U_1/U_0/U_0/state_reg[0]  ( .D(\U_1/U_0/U_0/nextState [0]), .CLK(CLK), 
        .R(n9517), .S(1'b1), .Q(\U_1/U_0/U_0/state[0] ) );
  DFFSR \U_1/U_0/U_0/si_reg[0]  ( .D(n7817), .CLK(CLK), .R(n9517), .S(1'b1), 
        .Q(\U_1/U_0/U_0/si[0] ) );
  DFFPOSX1 \U_1/U_0/U_0/permuteComplete_reg  ( .D(n7806), .CLK(CLK), .Q(
        \U_1/U_0/U_0/permuteComplete ) );
  DFFSR \U_1/U_0/U_0/state_reg[3]  ( .D(\U_1/U_0/U_0/nextState [3]), .CLK(CLK), 
        .R(n9517), .S(1'b1), .Q(\U_1/U_0/U_0/state[3] ) );
  DFFSR \U_1/U_0/U_0/state_reg[4]  ( .D(\U_1/U_0/U_0/nextState [4]), .CLK(CLK), 
        .R(n9517), .S(1'b1), .Q(\U_1/U_0/U_0/state[4] ) );
  DFFSR \U_1/U_0/U_0/state_reg[1]  ( .D(\U_1/U_0/U_0/nextState [1]), .CLK(CLK), 
        .R(n9517), .S(1'b1), .Q(\U_1/U_0/U_0/state[1] ) );
  DFFSR \U_1/U_0/U_0/PDATA_READY_reg  ( .D(n11882), .CLK(CLK), .R(n9517), .S(
        1'b1), .Q(\U_1/PDATA_READY ) );
  DFFSR \U_1/U_0/U_0/state_reg[2]  ( .D(\U_1/U_0/U_0/nextState [2]), .CLK(CLK), 
        .R(n9517), .S(1'b1), .Q(\U_1/U_0/U_0/state[2] ) );
  DFFPOSX1 \U_1/U_0/U_0/fr_enable_reg  ( .D(n7077), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fr_enable ) );
  DFFPOSX1 \U_1/U_0/U_0/R_ENABLE_reg  ( .D(n7076), .CLK(CLK), .Q(R_ENABLE_S)
         );
  DFFPOSX1 \U_1/U_0/U_0/fw_enable_reg  ( .D(n7075), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fw_enable ) );
  DFFPOSX1 \U_1/U_0/U_0/W_ENABLE_reg  ( .D(n7074), .CLK(CLK), .Q(W_ENABLE_S)
         );
  DFFPOSX1 \U_1/U_0/U_0/prefillCounter_reg[0]  ( .D(n7805), .CLK(CLK), .Q(
        \U_1/U_0/U_0/prefillCounter[0] ) );
  DFFPOSX1 \U_1/U_0/U_0/prefillCounter_reg[1]  ( .D(n7804), .CLK(CLK), .Q(
        \U_1/U_0/U_0/prefillCounter[1] ) );
  DFFPOSX1 \U_1/U_0/U_0/prefillCounter_reg[2]  ( .D(n7803), .CLK(CLK), .Q(
        \U_1/U_0/U_0/prefillCounter[2] ) );
  DFFPOSX1 \U_1/U_0/U_0/prefillCounter_reg[3]  ( .D(n7802), .CLK(CLK), .Q(
        \U_1/U_0/U_0/prefillCounter[3] ) );
  DFFPOSX1 \U_1/U_0/U_0/prefillCounter_reg[4]  ( .D(n7801), .CLK(CLK), .Q(
        \U_1/U_0/U_0/prefillCounter[4] ) );
  DFFPOSX1 \U_1/U_0/U_0/prefillCounter_reg[5]  ( .D(n7800), .CLK(CLK), .Q(
        \U_1/U_0/U_0/prefillCounter[5] ) );
  DFFPOSX1 \U_1/U_0/U_0/prefillCounter_reg[6]  ( .D(n7799), .CLK(CLK), .Q(
        \U_1/U_0/U_0/prefillCounter[6] ) );
  DFFPOSX1 \U_1/U_0/U_0/prefillCounter_reg[7]  ( .D(n7798), .CLK(CLK), .Q(
        \U_1/U_0/U_0/prefillCounter[7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[0][6]  ( .D(n10283), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[0][6] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[0][5]  ( .D(n10284), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[0][5] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[0][4]  ( .D(n10285), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[0][4] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[0][3]  ( .D(n7869), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[0][3] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[0][2]  ( .D(n7870), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[0][2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[0][1]  ( .D(n7871), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[0][1] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[0][0]  ( .D(n7872), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[0][0] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[1][7]  ( .D(n10286), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[1][7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[0][7]  ( .D(n10287), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[0][7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[7][0]  ( .D(n10288), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[7][0] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[7][1]  ( .D(n10289), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[7][1] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[7][2]  ( .D(n10290), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[7][2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[7][3]  ( .D(n10291), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[7][3] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[7][4]  ( .D(n10292), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[7][4] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[7][5]  ( .D(n10293), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[7][5] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[7][6]  ( .D(n10294), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[7][6] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[7][7]  ( .D(n10295), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[7][7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[6][0]  ( .D(n10296), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[6][0] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[6][1]  ( .D(n10297), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[6][1] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[6][2]  ( .D(n10298), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[6][2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[6][3]  ( .D(n10299), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[6][3] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[6][4]  ( .D(n10300), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[6][4] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[6][5]  ( .D(n10301), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[6][5] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[6][6]  ( .D(n10302), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[6][6] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[6][7]  ( .D(n10303), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[6][7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[5][0]  ( .D(n10304), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[5][0] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[5][1]  ( .D(n10305), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[5][1] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[5][2]  ( .D(n10306), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[5][2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[5][3]  ( .D(n10307), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[5][3] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[5][4]  ( .D(n10308), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[5][4] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[5][5]  ( .D(n10309), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[5][5] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[5][6]  ( .D(n10310), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[5][6] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[5][7]  ( .D(n10311), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[5][7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[4][0]  ( .D(n10312), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[4][0] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[4][1]  ( .D(n10313), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[4][1] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[4][2]  ( .D(n10314), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[4][2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[4][3]  ( .D(n10315), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[4][3] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[4][4]  ( .D(n10316), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[4][4] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[4][5]  ( .D(n10317), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[4][5] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[4][6]  ( .D(n10318), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[4][6] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[4][7]  ( .D(n10319), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[4][7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[3][0]  ( .D(n10320), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[3][0] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[3][1]  ( .D(n10321), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[3][1] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[3][2]  ( .D(n10322), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[3][2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[3][3]  ( .D(n10323), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[3][3] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[3][4]  ( .D(n10324), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[3][4] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[3][5]  ( .D(n10325), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[3][5] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[3][6]  ( .D(n10326), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[3][6] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[3][7]  ( .D(n10327), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[3][7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[2][0]  ( .D(n10328), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[2][0] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[2][1]  ( .D(n10329), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[2][1] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[2][2]  ( .D(n10330), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[2][2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[2][3]  ( .D(n10331), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[2][3] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[2][4]  ( .D(n10332), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[2][4] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[2][5]  ( .D(n10333), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[2][5] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[2][6]  ( .D(n10334), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[2][6] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[2][7]  ( .D(n10335), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[2][7] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[1][0]  ( .D(n10336), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[1][0] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[1][1]  ( .D(n10337), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[1][1] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[1][2]  ( .D(n10338), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[1][2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[1][3]  ( .D(n10339), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[1][3] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[1][4]  ( .D(n10340), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[1][4] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[1][5]  ( .D(n10341), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[1][5] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyTable_reg[1][6]  ( .D(n10342), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyTable[1][6] ) );
  DFFSR \U_1/U_0/U_0/si_reg[7]  ( .D(n7810), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/si[7] ) );
  DFFSR \U_1/U_0/U_0/si_reg[1]  ( .D(n7816), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/si[1] ) );
  DFFSR \U_1/U_0/U_0/si_reg[2]  ( .D(n7815), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/si[2] ) );
  DFFSR \U_1/U_0/U_0/si_reg[3]  ( .D(n7814), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/si[3] ) );
  DFFSR \U_1/U_0/U_0/si_reg[4]  ( .D(n7813), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/si[4] ) );
  DFFSR \U_1/U_0/U_0/si_reg[5]  ( .D(n7812), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/si[5] ) );
  DFFSR \U_1/U_0/U_0/si_reg[6]  ( .D(n7811), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/si[6] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyi_reg[2]  ( .D(n7809), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyi[2] ) );
  DFFPOSX1 \U_1/U_0/U_0/keyi_reg[1]  ( .D(n7808), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyi[1] ) );
  DFFSR \U_1/U_0/U_0/sj_reg[7]  ( .D(n7825), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/sj[7] ) );
  DFFSR \U_1/U_0/U_0/sj_reg[6]  ( .D(n7824), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/sj[6] ) );
  DFFSR \U_1/U_0/U_0/sj_reg[5]  ( .D(n7823), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/sj[5] ) );
  DFFSR \U_1/U_0/U_0/sj_reg[4]  ( .D(n7822), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/sj[4] ) );
  DFFSR \U_1/U_0/U_0/sj_reg[3]  ( .D(n7821), .CLK(CLK), .R(n9516), .S(1'b1), 
        .Q(\U_1/U_0/U_0/sj[3] ) );
  DFFSR \U_1/U_0/U_0/sj_reg[2]  ( .D(n7820), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/sj[2] ) );
  DFFSR \U_1/U_0/U_0/sj_reg[1]  ( .D(n7819), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/sj[1] ) );
  DFFSR \U_1/U_0/U_0/sj_reg[0]  ( .D(n7818), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/sj[0] ) );
  DFFPOSX1 \U_1/U_0/U_0/inti_reg[7]  ( .D(n7842), .CLK(CLK), .Q(
        \U_1/U_0/U_0/inti[7] ) );
  DFFPOSX1 \U_1/U_0/U_0/inti_reg[0]  ( .D(n7849), .CLK(CLK), .Q(
        \U_1/U_0/U_0/inti[0] ) );
  DFFPOSX1 \U_1/U_0/U_0/inti_reg[1]  ( .D(n7848), .CLK(CLK), .Q(
        \U_1/U_0/U_0/inti[1] ) );
  DFFPOSX1 \U_1/U_0/U_0/inti_reg[2]  ( .D(n7847), .CLK(CLK), .Q(
        \U_1/U_0/U_0/inti[2] ) );
  DFFPOSX1 \U_1/U_0/U_0/inti_reg[3]  ( .D(n7846), .CLK(CLK), .Q(
        \U_1/U_0/U_0/inti[3] ) );
  DFFPOSX1 \U_1/U_0/U_0/inti_reg[4]  ( .D(n7845), .CLK(CLK), .Q(
        \U_1/U_0/U_0/inti[4] ) );
  DFFPOSX1 \U_1/U_0/U_0/inti_reg[5]  ( .D(n7844), .CLK(CLK), .Q(
        \U_1/U_0/U_0/inti[5] ) );
  DFFPOSX1 \U_1/U_0/U_0/inti_reg[6]  ( .D(n7843), .CLK(CLK), .Q(
        \U_1/U_0/U_0/inti[6] ) );
  DFFPOSX1 \U_1/U_0/U_0/delaydata_reg[7]  ( .D(n10538), .CLK(CLK), .Q(
        \U_1/U_0/U_0/delaydata [7]) );
  DFFPOSX1 \U_1/U_0/U_0/delaydata_reg[0]  ( .D(n10537), .CLK(CLK), .Q(
        \U_1/U_0/U_0/delaydata [0]) );
  DFFPOSX1 \U_1/U_0/U_0/delaydata_reg[1]  ( .D(n10536), .CLK(CLK), .Q(
        \U_1/U_0/U_0/delaydata [1]) );
  DFFPOSX1 \U_1/U_0/U_0/delaydata_reg[2]  ( .D(n10535), .CLK(CLK), .Q(
        \U_1/U_0/U_0/delaydata [2]) );
  DFFPOSX1 \U_1/U_0/U_0/delaydata_reg[3]  ( .D(n10534), .CLK(CLK), .Q(
        \U_1/U_0/U_0/delaydata [3]) );
  DFFPOSX1 \U_1/U_0/U_0/delaydata_reg[4]  ( .D(n10533), .CLK(CLK), .Q(
        \U_1/U_0/U_0/delaydata [4]) );
  DFFPOSX1 \U_1/U_0/U_0/delaydata_reg[5]  ( .D(n10532), .CLK(CLK), .Q(
        \U_1/U_0/U_0/delaydata [5]) );
  DFFPOSX1 \U_1/U_0/U_0/delaydata_reg[6]  ( .D(n10531), .CLK(CLK), .Q(
        \U_1/U_0/U_0/delaydata [6]) );
  DFFPOSX1 \U_1/U_0/U_0/intj_reg[0]  ( .D(n7865), .CLK(CLK), .Q(
        \U_1/U_0/U_0/intj[0] ) );
  DFFPOSX1 \U_1/U_0/U_0/intj_reg[1]  ( .D(n7864), .CLK(CLK), .Q(
        \U_1/U_0/U_0/intj[1] ) );
  DFFPOSX1 \U_1/U_0/U_0/intj_reg[2]  ( .D(n7863), .CLK(CLK), .Q(
        \U_1/U_0/U_0/intj[2] ) );
  DFFPOSX1 \U_1/U_0/U_0/intj_reg[3]  ( .D(n7862), .CLK(CLK), .Q(
        \U_1/U_0/U_0/intj[3] ) );
  DFFPOSX1 \U_1/U_0/U_0/intj_reg[4]  ( .D(n7861), .CLK(CLK), .Q(
        \U_1/U_0/U_0/intj[4] ) );
  DFFPOSX1 \U_1/U_0/U_0/intj_reg[5]  ( .D(n7860), .CLK(CLK), .Q(
        \U_1/U_0/U_0/intj[5] ) );
  DFFPOSX1 \U_1/U_0/U_0/intj_reg[6]  ( .D(n7859), .CLK(CLK), .Q(
        \U_1/U_0/U_0/intj[6] ) );
  DFFPOSX1 \U_1/U_0/U_0/intj_reg[7]  ( .D(n7858), .CLK(CLK), .Q(
        \U_1/U_0/U_0/intj[7] ) );
  DFFPOSX1 \U_1/U_0/U_0/extratemp_reg[7]  ( .D(n10528), .CLK(CLK), .Q(
        \U_1/U_0/U_0/extratemp[7] ) );
  DFFPOSX1 \U_1/U_0/U_0/extratemp_reg[6]  ( .D(n10527), .CLK(CLK), .Q(
        \U_1/U_0/U_0/extratemp[6] ) );
  DFFPOSX1 \U_1/U_0/U_0/extratemp_reg[5]  ( .D(n10526), .CLK(CLK), .Q(
        \U_1/U_0/U_0/extratemp[5] ) );
  DFFPOSX1 \U_1/U_0/U_0/extratemp_reg[4]  ( .D(n10525), .CLK(CLK), .Q(
        \U_1/U_0/U_0/extratemp[4] ) );
  DFFPOSX1 \U_1/U_0/U_0/extratemp_reg[3]  ( .D(n10524), .CLK(CLK), .Q(
        \U_1/U_0/U_0/extratemp[3] ) );
  DFFPOSX1 \U_1/U_0/U_0/extratemp_reg[2]  ( .D(n10523), .CLK(CLK), .Q(
        \U_1/U_0/U_0/extratemp[2] ) );
  DFFPOSX1 \U_1/U_0/U_0/extratemp_reg[1]  ( .D(n10522), .CLK(CLK), .Q(
        \U_1/U_0/U_0/extratemp[1] ) );
  DFFPOSX1 \U_1/U_0/U_0/extratemp_reg[0]  ( .D(n10521), .CLK(CLK), .Q(
        \U_1/U_0/U_0/extratemp[0] ) );
  DFFPOSX1 \U_1/U_0/U_0/temp_reg[0]  ( .D(n7833), .CLK(CLK), .Q(
        \U_1/U_0/U_0/temp[0] ) );
  DFFSR \U_1/U_0/U_0/currentProcessedData_reg[0]  ( .D(
        \U_1/U_0/U_0/nextProcessedData[0] ), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/currentProcessedData [0]) );
  DFFPOSX1 \U_1/U_0/U_0/PROCESSED_DATA_reg[0]  ( .D(n10483), .CLK(CLK), .Q(
        \U_1/PROCESSED_DATA [0]) );
  DFFPOSX1 \U_1/U_0/U_0/ADDR_reg[0]  ( .D(n7056), .CLK(CLK), .Q(ADDR_S[0]) );
  DFFPOSX1 \U_1/U_0/U_0/faddr_reg[0]  ( .D(n10484), .CLK(CLK), .Q(
        \U_1/U_0/U_0/faddr [0]) );
  DFFPOSX1 \U_1/U_0/U_0/temp_reg[1]  ( .D(n7832), .CLK(CLK), .Q(
        \U_1/U_0/U_0/temp[1] ) );
  DFFPOSX1 \U_1/U_0/U_0/fdata_reg[1]  ( .D(n10485), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fdata [1]) );
  DFFPOSX1 \U_1/U_0/U_0/DATA_reg[1]  ( .D(n7053), .CLK(CLK), .Q(DATA_S[1]) );
  DFFSR \U_1/U_0/U_0/currentProcessedData_reg[1]  ( .D(
        \U_1/U_0/U_0/nextProcessedData[1] ), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/currentProcessedData [1]) );
  DFFPOSX1 \U_1/U_0/U_0/PROCESSED_DATA_reg[1]  ( .D(n10486), .CLK(CLK), .Q(
        \U_1/PROCESSED_DATA [1]) );
  DFFPOSX1 \U_1/U_0/U_0/ADDR_reg[1]  ( .D(n7050), .CLK(CLK), .Q(ADDR_S[1]) );
  DFFPOSX1 \U_1/U_0/U_0/faddr_reg[1]  ( .D(n10487), .CLK(CLK), .Q(
        \U_1/U_0/U_0/faddr [1]) );
  DFFPOSX1 \U_1/U_0/U_0/temp_reg[2]  ( .D(n7831), .CLK(CLK), .Q(
        \U_1/U_0/U_0/temp[2] ) );
  DFFPOSX1 \U_1/U_0/U_0/fdata_reg[2]  ( .D(n10488), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fdata [2]) );
  DFFPOSX1 \U_1/U_0/U_0/DATA_reg[2]  ( .D(n7047), .CLK(CLK), .Q(DATA_S[2]) );
  DFFSR \U_1/U_0/U_0/currentProcessedData_reg[2]  ( .D(
        \U_1/U_0/U_0/nextProcessedData[2] ), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/currentProcessedData [2]) );
  DFFPOSX1 \U_1/U_0/U_0/PROCESSED_DATA_reg[2]  ( .D(n10489), .CLK(CLK), .Q(
        \U_1/PROCESSED_DATA [2]) );
  DFFPOSX1 \U_1/U_0/U_0/ADDR_reg[2]  ( .D(n7044), .CLK(CLK), .Q(ADDR_S[2]) );
  DFFPOSX1 \U_1/U_0/U_0/faddr_reg[2]  ( .D(n10490), .CLK(CLK), .Q(
        \U_1/U_0/U_0/faddr [2]) );
  DFFPOSX1 \U_1/U_0/U_0/temp_reg[3]  ( .D(n7830), .CLK(CLK), .Q(
        \U_1/U_0/U_0/temp[3] ) );
  DFFPOSX1 \U_1/U_0/U_0/fdata_reg[3]  ( .D(n10491), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fdata [3]) );
  DFFPOSX1 \U_1/U_0/U_0/DATA_reg[3]  ( .D(n7041), .CLK(CLK), .Q(DATA_S[3]) );
  DFFSR \U_1/U_0/U_0/currentProcessedData_reg[3]  ( .D(
        \U_1/U_0/U_0/nextProcessedData[3] ), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/currentProcessedData [3]) );
  DFFPOSX1 \U_1/U_0/U_0/PROCESSED_DATA_reg[3]  ( .D(n10492), .CLK(CLK), .Q(
        \U_1/PROCESSED_DATA [3]) );
  DFFPOSX1 \U_1/U_0/U_0/ADDR_reg[3]  ( .D(n7038), .CLK(CLK), .Q(ADDR_S[3]) );
  DFFPOSX1 \U_1/U_0/U_0/faddr_reg[3]  ( .D(n10493), .CLK(CLK), .Q(
        \U_1/U_0/U_0/faddr [3]) );
  DFFPOSX1 \U_1/U_0/U_0/temp_reg[4]  ( .D(n7829), .CLK(CLK), .Q(
        \U_1/U_0/U_0/temp[4] ) );
  DFFPOSX1 \U_1/U_0/U_0/fdata_reg[4]  ( .D(n10494), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fdata [4]) );
  DFFPOSX1 \U_1/U_0/U_0/DATA_reg[4]  ( .D(n7035), .CLK(CLK), .Q(DATA_S[4]) );
  DFFSR \U_1/U_0/U_0/currentProcessedData_reg[4]  ( .D(
        \U_1/U_0/U_0/nextProcessedData[4] ), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/currentProcessedData [4]) );
  DFFPOSX1 \U_1/U_0/U_0/PROCESSED_DATA_reg[4]  ( .D(n10495), .CLK(CLK), .Q(
        \U_1/PROCESSED_DATA [4]) );
  DFFPOSX1 \U_1/U_0/U_0/ADDR_reg[4]  ( .D(n7032), .CLK(CLK), .Q(ADDR_S[4]) );
  DFFPOSX1 \U_1/U_0/U_0/faddr_reg[4]  ( .D(n10496), .CLK(CLK), .Q(
        \U_1/U_0/U_0/faddr [4]) );
  DFFPOSX1 \U_1/U_0/U_0/temp_reg[5]  ( .D(n7828), .CLK(CLK), .Q(
        \U_1/U_0/U_0/temp[5] ) );
  DFFPOSX1 \U_1/U_0/U_0/fdata_reg[5]  ( .D(n10497), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fdata [5]) );
  DFFPOSX1 \U_1/U_0/U_0/DATA_reg[5]  ( .D(n7029), .CLK(CLK), .Q(DATA_S[5]) );
  DFFSR \U_1/U_0/U_0/currentProcessedData_reg[5]  ( .D(
        \U_1/U_0/U_0/nextProcessedData[5] ), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/currentProcessedData [5]) );
  DFFPOSX1 \U_1/U_0/U_0/PROCESSED_DATA_reg[5]  ( .D(n10498), .CLK(CLK), .Q(
        \U_1/PROCESSED_DATA [5]) );
  DFFPOSX1 \U_1/U_0/U_0/ADDR_reg[5]  ( .D(n7026), .CLK(CLK), .Q(ADDR_S[5]) );
  DFFPOSX1 \U_1/U_0/U_0/faddr_reg[5]  ( .D(n10499), .CLK(CLK), .Q(
        \U_1/U_0/U_0/faddr [5]) );
  DFFPOSX1 \U_1/U_0/U_0/temp_reg[6]  ( .D(n7827), .CLK(CLK), .Q(
        \U_1/U_0/U_0/temp[6] ) );
  DFFPOSX1 \U_1/U_0/U_0/fdata_reg[6]  ( .D(n10500), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fdata [6]) );
  DFFPOSX1 \U_1/U_0/U_0/DATA_reg[6]  ( .D(n7023), .CLK(CLK), .Q(DATA_S[6]) );
  DFFSR \U_1/U_0/U_0/currentProcessedData_reg[6]  ( .D(
        \U_1/U_0/U_0/nextProcessedData[6] ), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/currentProcessedData [6]) );
  DFFPOSX1 \U_1/U_0/U_0/PROCESSED_DATA_reg[6]  ( .D(n10501), .CLK(CLK), .Q(
        \U_1/PROCESSED_DATA [6]) );
  DFFPOSX1 \U_1/U_0/U_0/ADDR_reg[6]  ( .D(n7020), .CLK(CLK), .Q(ADDR_S[6]) );
  DFFPOSX1 \U_1/U_0/U_0/faddr_reg[6]  ( .D(n10502), .CLK(CLK), .Q(
        \U_1/U_0/U_0/faddr [6]) );
  DFFPOSX1 \U_1/U_0/U_0/temp_reg[7]  ( .D(n7826), .CLK(CLK), .Q(
        \U_1/U_0/U_0/temp[7] ) );
  DFFPOSX1 \U_1/U_0/U_0/fdata_reg[7]  ( .D(n10503), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fdata [7]) );
  DFFPOSX1 \U_1/U_0/U_0/DATA_reg[7]  ( .D(n7017), .CLK(CLK), .Q(DATA_S[7]) );
  DFFSR \U_1/U_0/U_0/currentProcessedData_reg[7]  ( .D(
        \U_1/U_0/U_0/nextProcessedData[7] ), .CLK(CLK), .R(n9515), .S(1'b1), 
        .Q(\U_1/U_0/U_0/currentProcessedData [7]) );
  DFFPOSX1 \U_1/U_0/U_0/PROCESSED_DATA_reg[7]  ( .D(n10504), .CLK(CLK), .Q(
        \U_1/PROCESSED_DATA [7]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[0]  ( .D(n7784), .CLK(CLK), .R(n9515), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [0]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[8]  ( .D(n7776), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [8]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[2]  ( .D(n7782), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [2]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[10]  ( .D(n7774), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [10]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[3]  ( .D(n7781), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [3]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[11]  ( .D(n7773), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [11]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[4]  ( .D(n7780), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [4]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[12]  ( .D(n7772), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [12]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[5]  ( .D(n7779), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [5]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[13]  ( .D(n7771), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [13]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[6]  ( .D(n7778), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [6]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[14]  ( .D(n7770), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [14]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[7]  ( .D(n7777), .CLK(CLK), .R(n9514), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [7]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[15]  ( .D(n7769), .CLK(CLK), .R(n9513), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [15]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[1]  ( .D(n7783), .CLK(CLK), .R(n9513), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [1]) );
  DFFSR \U_1/U_3/U_1/current_crc_reg[9]  ( .D(n7775), .CLK(CLK), .R(n9513), 
        .S(1'b1), .Q(\U_1/U_3/TX_CRC [9]) );
  DFFPOSX1 \U_1/U_0/U_0/ADDR_reg[7]  ( .D(n6998), .CLK(CLK), .Q(ADDR_S[7]) );
  DFFPOSX1 \U_1/U_0/U_0/faddr_reg[7]  ( .D(n10505), .CLK(CLK), .Q(
        \U_1/U_0/U_0/faddr [7]) );
  DFFPOSX1 \U_1/U_0/U_0/fdata_reg[0]  ( .D(n10506), .CLK(CLK), .Q(
        \U_1/U_0/U_0/fdata [0]) );
  DFFPOSX1 \U_1/U_0/U_0/DATA_reg[0]  ( .D(n6995), .CLK(CLK), .Q(DATA_S[0]) );
  DFFPOSX1 \U_1/U_0/U_0/keyi_reg[0]  ( .D(n7807), .CLK(CLK), .Q(
        \U_1/U_0/U_0/keyi[0] ) );
  DFFPOSX1 \U_1/U_1/U_0/tempOpcode_reg[1]  ( .D(n6994), .CLK(CLK), .Q(
        \U_1/U_1/U_0/tempOpcode [1]) );
  DFFPOSX1 \U_1/U_3/U_3/flop_data_reg[7]  ( .D(n7751), .CLK(CLK), .Q(
        \U_1/U_3/U_3/flop_data [7]) );
  DFFPOSX1 \U_1/U_3/U_3/flop_data_reg[0]  ( .D(n10517), .CLK(CLK), .Q(
        \U_1/U_3/U_3/flop_data [0]) );
  DFFPOSX1 \U_1/U_3/U_3/flop_data_reg[1]  ( .D(n10516), .CLK(CLK), .Q(
        \U_1/U_3/U_3/flop_data [1]) );
  DFFPOSX1 \U_1/U_3/U_3/flop_data_reg[2]  ( .D(n10515), .CLK(CLK), .Q(
        \U_1/U_3/U_3/flop_data [2]) );
  DFFPOSX1 \U_1/U_3/U_3/flop_data_reg[3]  ( .D(n10514), .CLK(CLK), .Q(
        \U_1/U_3/U_3/flop_data [3]) );
  DFFPOSX1 \U_1/U_3/U_3/flop_data_reg[4]  ( .D(n10513), .CLK(CLK), .Q(
        \U_1/U_3/U_3/flop_data [4]) );
  DFFPOSX1 \U_1/U_3/U_3/flop_data_reg[5]  ( .D(n10512), .CLK(CLK), .Q(
        \U_1/U_3/U_3/flop_data [5]) );
  DFFPOSX1 \U_1/U_3/U_3/flop_data_reg[6]  ( .D(n10511), .CLK(CLK), .Q(
        \U_1/U_3/U_3/flop_data [6]) );
  DFFPOSX1 \U_1/U_3/U_3/current_send_data_reg[6]  ( .D(n6993), .CLK(CLK), .Q(
        \U_1/U_3/U_3/current_send_data [6]) );
  DFFPOSX1 \U_1/U_3/U_3/send_data_reg[6]  ( .D(n6992), .CLK(CLK), .Q(
        \U_1/U_3/send_data [6]) );
  DFFPOSX1 \U_1/U_3/U_3/current_send_data_reg[5]  ( .D(n6991), .CLK(CLK), .Q(
        \U_1/U_3/U_3/current_send_data [5]) );
  DFFPOSX1 \U_1/U_3/U_3/send_data_reg[5]  ( .D(n6990), .CLK(CLK), .Q(
        \U_1/U_3/send_data [5]) );
  DFFPOSX1 \U_1/U_3/U_3/current_send_data_reg[4]  ( .D(n6989), .CLK(CLK), .Q(
        \U_1/U_3/U_3/current_send_data [4]) );
  DFFPOSX1 \U_1/U_3/U_3/send_data_reg[4]  ( .D(n6988), .CLK(CLK), .Q(
        \U_1/U_3/send_data [4]) );
  DFFPOSX1 \U_1/U_3/U_3/current_send_data_reg[3]  ( .D(n6987), .CLK(CLK), .Q(
        \U_1/U_3/U_3/current_send_data [3]) );
  DFFPOSX1 \U_1/U_3/U_3/send_data_reg[3]  ( .D(n6986), .CLK(CLK), .Q(
        \U_1/U_3/send_data [3]) );
  DFFPOSX1 \U_1/U_3/U_3/current_send_data_reg[2]  ( .D(n6985), .CLK(CLK), .Q(
        \U_1/U_3/U_3/current_send_data [2]) );
  DFFPOSX1 \U_1/U_3/U_3/send_data_reg[2]  ( .D(n6984), .CLK(CLK), .Q(
        \U_1/U_3/send_data [2]) );
  DFFPOSX1 \U_1/U_3/U_3/current_send_data_reg[1]  ( .D(n6983), .CLK(CLK), .Q(
        \U_1/U_3/U_3/current_send_data [1]) );
  DFFPOSX1 \U_1/U_3/U_3/send_data_reg[1]  ( .D(n6982), .CLK(CLK), .Q(
        \U_1/U_3/send_data [1]) );
  DFFPOSX1 \U_1/U_3/U_3/current_send_data_reg[0]  ( .D(n6981), .CLK(CLK), .Q(
        \U_1/U_3/U_3/current_send_data [0]) );
  DFFPOSX1 \U_1/U_3/U_3/send_data_reg[0]  ( .D(n6980), .CLK(CLK), .Q(
        \U_1/U_3/send_data [0]) );
  DFFPOSX1 \U_1/U_3/U_3/current_send_data_reg[7]  ( .D(n6979), .CLK(CLK), .Q(
        \U_1/U_3/U_3/current_send_data [7]) );
  DFFPOSX1 \U_1/U_3/U_3/send_data_reg[7]  ( .D(n6978), .CLK(CLK), .Q(
        \U_1/U_3/send_data [7]) );
  DFFSR \U_1/U_3/U_4/state_reg  ( .D(slave_is_sending), .CLK(CLK), .R(n9513), 
        .S(1'b1), .Q(\U_1/U_3/U_4/state ) );
  DFFSR \U_1/U_3/U_4/count_reg[0]  ( .D(\U_1/U_3/U_4/nextcount [0]), .CLK(CLK), 
        .R(n9513), .S(1'b1), .Q(\U_1/U_3/U_4/count[0] ) );
  DFFSR \U_1/U_3/U_4/count_reg[2]  ( .D(\U_1/U_3/U_4/nextcount [2]), .CLK(CLK), 
        .R(n9513), .S(1'b1), .Q(\U_1/U_3/U_4/count[2] ) );
  DFFSR \U_1/U_3/U_4/count_reg[3]  ( .D(\U_1/U_3/U_4/nextcount [3]), .CLK(CLK), 
        .R(n9513), .S(1'b1), .Q(\U_1/U_3/U_4/count[3] ) );
  DFFSR \U_1/U_3/U_4/count_reg[1]  ( .D(\U_1/U_3/U_4/nextcount [1]), .CLK(CLK), 
        .R(n9513), .S(1'b1), .Q(\U_1/U_3/U_4/count[1] ) );
  DFFSR \U_1/U_3/U_2/count_reg[1]  ( .D(n7767), .CLK(CLK), .R(1'b1), .S(n9522), 
        .Q(\U_1/U_3/U_2/count[1] ) );
  DFFSR \U_1/U_3/U_2/count_reg[2]  ( .D(n7766), .CLK(CLK), .R(1'b1), .S(n9522), 
        .Q(\U_1/U_3/U_2/count[2] ) );
  DFFSR \U_1/U_3/U_2/count_reg[0]  ( .D(n11625), .CLK(CLK), .R(1'b1), .S(n9522), .Q(\U_1/U_3/U_2/count[0] ) );
  DFFSR \U_1/U_3/U_2/present_val_reg[7]  ( .D(n11626), .CLK(CLK), .R(n9513), 
        .S(1'b1), .Q(\U_1/U_3/U_2/present_val [7]) );
  DFFSR \U_1/U_3/U_2/present_val_reg[6]  ( .D(n7759), .CLK(CLK), .R(n9513), 
        .S(1'b1), .Q(\U_1/U_3/U_2/present_val [6]) );
  DFFSR \U_1/U_3/U_2/present_val_reg[5]  ( .D(n7760), .CLK(CLK), .R(n9513), 
        .S(1'b1), .Q(\U_1/U_3/U_2/present_val [5]) );
  DFFSR \U_1/U_3/U_2/present_val_reg[4]  ( .D(n7761), .CLK(CLK), .R(n9513), 
        .S(1'b1), .Q(\U_1/U_3/U_2/present_val [4]) );
  DFFSR \U_1/U_3/U_2/present_val_reg[3]  ( .D(n7762), .CLK(CLK), .R(n9500), 
        .S(1'b1), .Q(\U_1/U_3/U_2/present_val [3]) );
  DFFSR \U_1/U_3/U_2/present_val_reg[2]  ( .D(n7763), .CLK(CLK), .R(n9497), 
        .S(1'b1), .Q(\U_1/U_3/U_2/present_val [2]) );
  DFFSR \U_1/U_3/U_2/present_val_reg[1]  ( .D(n7764), .CLK(CLK), .R(n9498), 
        .S(1'b1), .Q(\U_1/U_3/U_2/present_val [1]) );
  DFFSR \U_1/U_3/U_2/present_val_reg[0]  ( .D(n7765), .CLK(CLK), .R(n9499), 
        .S(1'b1), .Q(\U_1/U_3/d_encode ) );
  DFFSR \U_1/U_3/U_0/DE_holdout_BS_reg  ( .D(n7757), .CLK(CLK), .R(n9516), .S(
        1'b1), .Q(\U_1/U_3/U_0/DE_holdout_BS ) );
  DFFSR \U_1/U_3/U_0/dm_tx_out_reg  ( .D(\U_1/U_3/U_0/dm_tx_nxt ), .CLK(CLK), 
        .R(n9517), .S(1'b1), .Q(DMTH) );
  NAND2X1 U1 ( .A(n177), .B(n178), .Y(n6978) );
  AOI22X1 U2 ( .A(\U_1/U_3/U_3/current_send_data [7]), .B(n179), .C(
        \U_1/U_3/send_data [7]), .D(RST), .Y(n177) );
  OAI21X1 U3 ( .A(n180), .B(n12069), .C(n178), .Y(n6979) );
  AOI21X1 U4 ( .A(n182), .B(\U_1/U_3/TX_CRC [15]), .C(n10508), .Y(n178) );
  OAI21X1 U6 ( .A(n185), .B(n186), .C(n9512), .Y(n184) );
  OAI21X1 U7 ( .A(n187), .B(n12035), .C(n189), .Y(n186) );
  OAI21X1 U8 ( .A(\U_1/U_3/TX_CRC [7]), .B(\U_1/U_3/U_3/N188 ), .C(n190), .Y(
        n189) );
  NOR2X1 U9 ( .A(n191), .B(n12054), .Y(n185) );
  NAND2X1 U11 ( .A(n193), .B(n194), .Y(n6980) );
  AOI22X1 U12 ( .A(\U_1/U_3/U_3/current_send_data [0]), .B(n179), .C(
        \U_1/U_3/send_data [0]), .D(RST), .Y(n193) );
  OAI21X1 U13 ( .A(n180), .B(n12067), .C(n194), .Y(n6981) );
  AOI22X1 U15 ( .A(\U_1/U_3/U_3/flop_data [0]), .B(n198), .C(
        \U_1/U_3/TX_CRC [0]), .D(n10507), .Y(n197) );
  AOI22X1 U16 ( .A(\U_1/PROCESSED_DATA [0]), .B(n200), .C(\U_1/U_3/TX_CRC [8]), 
        .D(n182), .Y(n196) );
  NAND2X1 U18 ( .A(n201), .B(n202), .Y(n6982) );
  AOI22X1 U19 ( .A(\U_1/U_3/U_3/current_send_data [1]), .B(n179), .C(
        \U_1/U_3/send_data [1]), .D(RST), .Y(n201) );
  OAI21X1 U20 ( .A(n180), .B(n12065), .C(n202), .Y(n6983) );
  AOI22X1 U22 ( .A(\U_1/U_3/U_3/flop_data [1]), .B(n198), .C(
        \U_1/U_3/TX_CRC [1]), .D(n10507), .Y(n205) );
  AOI22X1 U23 ( .A(\U_1/PROCESSED_DATA [1]), .B(n200), .C(\U_1/U_3/TX_CRC [9]), 
        .D(n182), .Y(n204) );
  NAND2X1 U25 ( .A(n206), .B(n207), .Y(n6984) );
  AOI22X1 U26 ( .A(\U_1/U_3/U_3/current_send_data [2]), .B(n179), .C(
        \U_1/U_3/send_data [2]), .D(RST), .Y(n206) );
  OAI21X1 U27 ( .A(n180), .B(n12063), .C(n207), .Y(n6985) );
  AOI22X1 U29 ( .A(\U_1/U_3/U_3/flop_data [2]), .B(n198), .C(
        \U_1/U_3/TX_CRC [2]), .D(n10507), .Y(n210) );
  AOI22X1 U30 ( .A(\U_1/PROCESSED_DATA [2]), .B(n200), .C(\U_1/U_3/TX_CRC [10]), .D(n182), .Y(n209) );
  NAND2X1 U32 ( .A(n211), .B(n212), .Y(n6986) );
  AOI22X1 U33 ( .A(\U_1/U_3/U_3/current_send_data [3]), .B(n179), .C(
        \U_1/U_3/send_data [3]), .D(RST), .Y(n211) );
  OAI21X1 U34 ( .A(n180), .B(n12061), .C(n212), .Y(n6987) );
  AOI22X1 U36 ( .A(\U_1/U_3/U_3/flop_data [3]), .B(n198), .C(
        \U_1/U_3/TX_CRC [3]), .D(n10507), .Y(n215) );
  AOI22X1 U37 ( .A(\U_1/PROCESSED_DATA [3]), .B(n200), .C(\U_1/U_3/TX_CRC [11]), .D(n182), .Y(n214) );
  NAND2X1 U39 ( .A(n216), .B(n217), .Y(n6988) );
  AOI22X1 U40 ( .A(\U_1/U_3/U_3/current_send_data [4]), .B(n179), .C(
        \U_1/U_3/send_data [4]), .D(RST), .Y(n216) );
  OAI21X1 U41 ( .A(n180), .B(n12059), .C(n217), .Y(n6989) );
  AOI22X1 U43 ( .A(\U_1/U_3/U_3/flop_data [4]), .B(n198), .C(
        \U_1/U_3/TX_CRC [4]), .D(n10507), .Y(n220) );
  AOI22X1 U44 ( .A(\U_1/PROCESSED_DATA [4]), .B(n200), .C(\U_1/U_3/TX_CRC [12]), .D(n182), .Y(n219) );
  NAND2X1 U46 ( .A(n221), .B(n222), .Y(n6990) );
  AOI22X1 U47 ( .A(\U_1/U_3/U_3/current_send_data [5]), .B(n179), .C(
        \U_1/U_3/send_data [5]), .D(RST), .Y(n221) );
  OAI21X1 U49 ( .A(n180), .B(n12057), .C(n222), .Y(n6991) );
  AOI22X1 U52 ( .A(\U_1/U_3/U_3/flop_data [5]), .B(n198), .C(
        \U_1/U_3/TX_CRC [5]), .D(n10507), .Y(n225) );
  AOI22X1 U67 ( .A(\U_1/PROCESSED_DATA [5]), .B(n200), .C(\U_1/U_3/TX_CRC [13]), .D(n182), .Y(n224) );
  NAND2X1 U70 ( .A(n226), .B(n227), .Y(n6992) );
  AOI22X1 U96 ( .A(\U_1/U_3/U_3/current_send_data [6]), .B(n179), .C(
        \U_1/U_3/send_data [6]), .D(RST), .Y(n226) );
  OAI21X1 U98 ( .A(n180), .B(n12055), .C(n227), .Y(n6993) );
  AOI22X1 U100 ( .A(\U_1/U_3/U_3/flop_data [6]), .B(n198), .C(
        \U_1/U_3/TX_CRC [6]), .D(n10507), .Y(n231) );
  NAND3X1 U102 ( .A(n9534), .B(n11644), .C(n190), .Y(n232) );
  NOR2X1 U103 ( .A(n191), .B(RST), .Y(n198) );
  AOI22X1 U104 ( .A(\U_1/PROCESSED_DATA [6]), .B(n200), .C(
        \U_1/U_3/TX_CRC [14]), .D(n182), .Y(n230) );
  NOR2X1 U105 ( .A(n11652), .B(RST), .Y(n182) );
  NOR2X1 U106 ( .A(n187), .B(RST), .Y(n200) );
  NOR2X1 U108 ( .A(n228), .B(RST), .Y(n180) );
  OAI21X1 U109 ( .A(n11656), .B(n236), .C(n237), .Y(n228) );
  OAI22X1 U110 ( .A(n238), .B(n11840), .C(n240), .D(n12053), .Y(n6994) );
  OAI21X1 U112 ( .A(RST), .B(n10559), .C(n243), .Y(n6995) );
  NAND2X1 U113 ( .A(DATA_S[0]), .B(RST), .Y(n243) );
  AOI22X1 U116 ( .A(RST), .B(\U_1/U_0/U_0/fdata [0]), .C(n9523), .D(
        \U_1/U_0/U_0/nfdata[0] ), .Y(n244) );
  AOI22X1 U118 ( .A(RST), .B(\U_1/U_0/U_0/faddr [7]), .C(n9507), .D(
        \U_1/U_0/U_0/nfaddr[7] ), .Y(n245) );
  OAI21X1 U119 ( .A(RST), .B(n11880), .C(n247), .Y(n6998) );
  NAND2X1 U120 ( .A(ADDR_S[7]), .B(RST), .Y(n247) );
  AOI22X1 U123 ( .A(RST), .B(\U_1/PROCESSED_DATA [7]), .C(n9506), .D(
        \U_1/U_0/U_0/nextProcessedData[7] ), .Y(n248) );
  OAI21X1 U124 ( .A(RST), .B(n10552), .C(n250), .Y(n7017) );
  NAND2X1 U125 ( .A(DATA_S[7]), .B(RST), .Y(n250) );
  AOI22X1 U128 ( .A(RST), .B(\U_1/U_0/U_0/fdata [7]), .C(n9505), .D(
        \U_1/U_0/U_0/nfdata[7] ), .Y(n251) );
  AOI22X1 U130 ( .A(RST), .B(\U_1/U_0/U_0/faddr [6]), .C(n9504), .D(
        \U_1/U_0/U_0/nfaddr[6] ), .Y(n252) );
  OAI21X1 U131 ( .A(RST), .B(n11879), .C(n254), .Y(n7020) );
  NAND2X1 U132 ( .A(ADDR_S[6]), .B(RST), .Y(n254) );
  AOI22X1 U135 ( .A(RST), .B(\U_1/PROCESSED_DATA [6]), .C(n9503), .D(
        \U_1/U_0/U_0/nextProcessedData[6] ), .Y(n255) );
  OAI21X1 U136 ( .A(RST), .B(n10553), .C(n257), .Y(n7023) );
  NAND2X1 U137 ( .A(DATA_S[6]), .B(RST), .Y(n257) );
  AOI22X1 U140 ( .A(RST), .B(\U_1/U_0/U_0/fdata [6]), .C(n9502), .D(
        \U_1/U_0/U_0/nfdata[6] ), .Y(n258) );
  AOI22X1 U142 ( .A(RST), .B(\U_1/U_0/U_0/faddr [5]), .C(n9501), .D(
        \U_1/U_0/U_0/nfaddr[5] ), .Y(n259) );
  OAI21X1 U143 ( .A(RST), .B(n11878), .C(n261), .Y(n7026) );
  NAND2X1 U144 ( .A(ADDR_S[5]), .B(RST), .Y(n261) );
  AOI22X1 U147 ( .A(RST), .B(\U_1/PROCESSED_DATA [5]), .C(n9510), .D(
        \U_1/U_0/U_0/nextProcessedData[5] ), .Y(n262) );
  OAI21X1 U148 ( .A(RST), .B(n10554), .C(n264), .Y(n7029) );
  NAND2X1 U149 ( .A(DATA_S[5]), .B(RST), .Y(n264) );
  AOI22X1 U152 ( .A(RST), .B(\U_1/U_0/U_0/fdata [5]), .C(n9509), .D(
        \U_1/U_0/U_0/nfdata[5] ), .Y(n265) );
  AOI22X1 U154 ( .A(RST), .B(\U_1/U_0/U_0/faddr [4]), .C(n9512), .D(
        \U_1/U_0/U_0/nfaddr[4] ), .Y(n266) );
  OAI21X1 U155 ( .A(RST), .B(n11877), .C(n268), .Y(n7032) );
  NAND2X1 U156 ( .A(ADDR_S[4]), .B(RST), .Y(n268) );
  AOI22X1 U159 ( .A(RST), .B(\U_1/PROCESSED_DATA [4]), .C(n9511), .D(
        \U_1/U_0/U_0/nextProcessedData[4] ), .Y(n269) );
  OAI21X1 U160 ( .A(RST), .B(n10555), .C(n271), .Y(n7035) );
  NAND2X1 U161 ( .A(DATA_S[4]), .B(RST), .Y(n271) );
  AOI22X1 U164 ( .A(RST), .B(\U_1/U_0/U_0/fdata [4]), .C(n9527), .D(
        \U_1/U_0/U_0/nfdata[4] ), .Y(n272) );
  AOI22X1 U166 ( .A(RST), .B(\U_1/U_0/U_0/faddr [3]), .C(n9527), .D(
        \U_1/U_0/U_0/nfaddr[3] ), .Y(n273) );
  OAI21X1 U167 ( .A(RST), .B(n11876), .C(n275), .Y(n7038) );
  NAND2X1 U168 ( .A(ADDR_S[3]), .B(RST), .Y(n275) );
  AOI22X1 U171 ( .A(RST), .B(\U_1/PROCESSED_DATA [3]), .C(n9527), .D(
        \U_1/U_0/U_0/nextProcessedData[3] ), .Y(n276) );
  OAI21X1 U172 ( .A(RST), .B(n10556), .C(n278), .Y(n7041) );
  NAND2X1 U173 ( .A(DATA_S[3]), .B(RST), .Y(n278) );
  AOI22X1 U176 ( .A(RST), .B(\U_1/U_0/U_0/fdata [3]), .C(n9527), .D(
        \U_1/U_0/U_0/nfdata[3] ), .Y(n279) );
  AOI22X1 U178 ( .A(RST), .B(\U_1/U_0/U_0/faddr [2]), .C(n9527), .D(
        \U_1/U_0/U_0/nfaddr[2] ), .Y(n280) );
  OAI21X1 U179 ( .A(RST), .B(n11875), .C(n282), .Y(n7044) );
  NAND2X1 U180 ( .A(ADDR_S[2]), .B(RST), .Y(n282) );
  AOI22X1 U183 ( .A(RST), .B(\U_1/PROCESSED_DATA [2]), .C(n9527), .D(
        \U_1/U_0/U_0/nextProcessedData[2] ), .Y(n283) );
  OAI21X1 U184 ( .A(RST), .B(n10557), .C(n285), .Y(n7047) );
  NAND2X1 U185 ( .A(DATA_S[2]), .B(RST), .Y(n285) );
  AOI22X1 U188 ( .A(RST), .B(\U_1/U_0/U_0/fdata [2]), .C(n9527), .D(
        \U_1/U_0/U_0/nfdata[2] ), .Y(n286) );
  AOI22X1 U190 ( .A(RST), .B(\U_1/U_0/U_0/faddr [1]), .C(n9527), .D(
        \U_1/U_0/U_0/nfaddr[1] ), .Y(n287) );
  OAI21X1 U191 ( .A(RST), .B(n11874), .C(n289), .Y(n7050) );
  NAND2X1 U192 ( .A(ADDR_S[1]), .B(RST), .Y(n289) );
  AOI22X1 U195 ( .A(RST), .B(\U_1/PROCESSED_DATA [1]), .C(n9527), .D(
        \U_1/U_0/U_0/nextProcessedData[1] ), .Y(n290) );
  OAI21X1 U196 ( .A(RST), .B(n10558), .C(n292), .Y(n7053) );
  NAND2X1 U197 ( .A(DATA_S[1]), .B(RST), .Y(n292) );
  AOI22X1 U200 ( .A(RST), .B(\U_1/U_0/U_0/fdata [1]), .C(n9527), .D(
        \U_1/U_0/U_0/nfdata[1] ), .Y(n293) );
  AOI22X1 U202 ( .A(RST), .B(\U_1/U_0/U_0/faddr [0]), .C(n9527), .D(
        \U_1/U_0/U_0/nfaddr[0] ), .Y(n294) );
  OAI21X1 U203 ( .A(RST), .B(n11873), .C(n296), .Y(n7056) );
  NAND2X1 U204 ( .A(ADDR_S[0]), .B(RST), .Y(n296) );
  AOI22X1 U207 ( .A(RST), .B(\U_1/PROCESSED_DATA [0]), .C(n9527), .D(
        \U_1/U_0/U_0/nextProcessedData[0] ), .Y(n297) );
  OAI21X1 U208 ( .A(RST), .B(n298), .C(n299), .Y(n7074) );
  NAND2X1 U209 ( .A(W_ENABLE_S), .B(RST), .Y(n299) );
  AOI21X1 U210 ( .A(\U_1/U_0/U_0/fw_enable ), .B(n300), .C(n301), .Y(n298) );
  OAI21X1 U211 ( .A(RST), .B(n11893), .C(n303), .Y(n7075) );
  OAI21X1 U212 ( .A(RST), .B(n300), .C(\U_1/U_0/U_0/fw_enable ), .Y(n303) );
  NAND3X1 U214 ( .A(n304), .B(n9179), .C(n306), .Y(n301) );
  NOR2X1 U215 ( .A(n307), .B(n308), .Y(n306) );
  OAI21X1 U216 ( .A(RST), .B(n309), .C(n310), .Y(n7076) );
  NAND2X1 U217 ( .A(R_ENABLE_S), .B(RST), .Y(n310) );
  AOI21X1 U218 ( .A(\U_1/U_0/U_0/fr_enable ), .B(n311), .C(n312), .Y(n309) );
  OAI21X1 U219 ( .A(RST), .B(n11897), .C(n314), .Y(n7077) );
  OAI21X1 U220 ( .A(RST), .B(n311), .C(\U_1/U_0/U_0/fr_enable ), .Y(n314) );
  NAND3X1 U221 ( .A(n315), .B(n316), .C(n317), .Y(n311) );
  NAND3X1 U225 ( .A(n321), .B(n322), .C(n11912), .Y(n312) );
  OAI21X1 U226 ( .A(n9534), .B(n11865), .C(n325), .Y(n7091) );
  AOI22X1 U227 ( .A(n326), .B(\U_1/U_1/U_0/tempOpcode [1]), .C(
        \U_1/U_1/OUT_OPCODE [1]), .D(n10509), .Y(n325) );
  OAI21X1 U228 ( .A(n9534), .B(n11864), .C(n329), .Y(n7092) );
  AOI22X1 U229 ( .A(\U_1/U_1/U_0/tempData [0]), .B(n326), .C(\U_1/U_1/DATA [0]), .D(n10509), .Y(n329) );
  OAI22X1 U231 ( .A(n238), .B(n11831), .C(n240), .D(n11863), .Y(n7093) );
  OAI21X1 U233 ( .A(n9534), .B(n11862), .C(n333), .Y(n7094) );
  AOI22X1 U234 ( .A(\U_1/U_1/U_0/tempData [1]), .B(n326), .C(\U_1/U_1/DATA [1]), .D(n10509), .Y(n333) );
  OAI22X1 U236 ( .A(n238), .B(n11832), .C(n240), .D(n11861), .Y(n7095) );
  OAI21X1 U238 ( .A(n9534), .B(n11860), .C(n337), .Y(n7096) );
  AOI22X1 U239 ( .A(\U_1/U_1/U_0/tempData [2]), .B(n326), .C(\U_1/U_1/DATA [2]), .D(n10509), .Y(n337) );
  OAI22X1 U241 ( .A(n238), .B(n11833), .C(n240), .D(n11859), .Y(n7097) );
  OAI21X1 U243 ( .A(n9534), .B(n11858), .C(n341), .Y(n7098) );
  AOI22X1 U244 ( .A(\U_1/U_1/U_0/tempData [3]), .B(n326), .C(\U_1/U_1/DATA [3]), .D(n10509), .Y(n341) );
  OAI22X1 U246 ( .A(n238), .B(n11834), .C(n240), .D(n11857), .Y(n7099) );
  OAI21X1 U248 ( .A(n9533), .B(n11856), .C(n345), .Y(n7100) );
  AOI22X1 U249 ( .A(\U_1/U_1/U_0/tempData [4]), .B(n326), .C(\U_1/U_1/DATA [4]), .D(n10509), .Y(n345) );
  OAI22X1 U251 ( .A(n238), .B(n11835), .C(n240), .D(n11855), .Y(n7101) );
  OAI21X1 U253 ( .A(n9534), .B(n11854), .C(n349), .Y(n7102) );
  AOI22X1 U254 ( .A(\U_1/U_1/U_0/tempData [5]), .B(n326), .C(\U_1/U_1/DATA [5]), .D(n10509), .Y(n349) );
  OAI22X1 U256 ( .A(n238), .B(n11836), .C(n240), .D(n11853), .Y(n7103) );
  OAI21X1 U258 ( .A(n9533), .B(n11852), .C(n353), .Y(n7104) );
  AOI22X1 U259 ( .A(\U_1/U_1/U_0/tempData [6]), .B(n326), .C(\U_1/U_1/DATA [6]), .D(n10509), .Y(n353) );
  OAI22X1 U261 ( .A(n238), .B(n11837), .C(n240), .D(n11851), .Y(n7105) );
  OAI21X1 U263 ( .A(n9534), .B(n11850), .C(n357), .Y(n7106) );
  AOI22X1 U264 ( .A(\U_1/U_1/U_0/tempData [7]), .B(n326), .C(\U_1/U_1/DATA [7]), .D(n10509), .Y(n357) );
  OAI22X1 U266 ( .A(n238), .B(n11838), .C(n240), .D(n11849), .Y(n7107) );
  OAI22X1 U268 ( .A(n238), .B(n11839), .C(n240), .D(n11848), .Y(n7108) );
  NOR2X1 U270 ( .A(n362), .B(RST), .Y(n240) );
  OAI21X1 U271 ( .A(n9534), .B(n11847), .C(n364), .Y(n7109) );
  AOI22X1 U272 ( .A(\U_1/U_1/U_0/tempOpcode [0]), .B(n326), .C(
        \U_1/U_1/OUT_OPCODE [0]), .D(n10509), .Y(n364) );
  NAND2X1 U275 ( .A(\U_1/U_1/U_0/state[2] ), .B(n11841), .Y(n362) );
  OAI21X1 U276 ( .A(n9534), .B(n11844), .C(n238), .Y(n7110) );
  NAND3X1 U277 ( .A(n11842), .B(n11843), .C(n369), .Y(n238) );
  NOR2X1 U278 ( .A(RST), .B(n11657), .Y(n369) );
  AOI22X1 U280 ( .A(EMPTY_S), .B(RST), .C(\U_1/U_1/U_1/N349 ), .D(n9522), .Y(
        n371) );
  AOI22X1 U282 ( .A(FULL_S), .B(RST), .C(\U_1/U_1/U_1/N355 ), .D(n9522), .Y(
        n372) );
  OAI21X1 U283 ( .A(n9533), .B(n11660), .C(n374), .Y(n7130) );
  NAND3X1 U284 ( .A(n11843), .B(n11657), .C(n375), .Y(n374) );
  NOR2X1 U285 ( .A(RST), .B(n11842), .Y(n375) );
  OAI22X1 U287 ( .A(n9532), .B(n11632), .C(RST), .D(n11631), .Y(n7140) );
  OAI22X1 U289 ( .A(n9532), .B(n11543), .C(RST), .D(n11542), .Y(n7207) );
  AOI22X1 U292 ( .A(RST), .B(\U_1/U_0/PLAINKEY [62]), .C(n9527), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[62] ), .Y(n380) );
  AOI22X1 U294 ( .A(RST), .B(\U_1/U_0/PLAINKEY [61]), .C(n9527), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[61] ), .Y(n381) );
  AOI22X1 U296 ( .A(RST), .B(\U_1/U_0/PLAINKEY [60]), .C(n9527), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[60] ), .Y(n382) );
  AOI22X1 U298 ( .A(RST), .B(\U_1/U_0/PLAINKEY [59]), .C(n9527), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[59] ), .Y(n383) );
  AOI22X1 U300 ( .A(RST), .B(\U_1/U_0/PLAINKEY [58]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[58] ), .Y(n384) );
  AOI22X1 U302 ( .A(RST), .B(\U_1/U_0/PLAINKEY [57]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[57] ), .Y(n385) );
  AOI22X1 U304 ( .A(RST), .B(\U_1/U_0/PLAINKEY [56]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[56] ), .Y(n386) );
  AOI22X1 U306 ( .A(RST), .B(\U_1/U_0/PLAINKEY [55]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[55] ), .Y(n387) );
  AOI22X1 U308 ( .A(RST), .B(\U_1/U_0/PLAINKEY [54]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[54] ), .Y(n388) );
  AOI22X1 U310 ( .A(RST), .B(\U_1/U_0/PLAINKEY [53]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[53] ), .Y(n389) );
  AOI22X1 U312 ( .A(RST), .B(\U_1/U_0/PLAINKEY [52]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[52] ), .Y(n390) );
  AOI22X1 U314 ( .A(RST), .B(\U_1/U_0/PLAINKEY [51]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[51] ), .Y(n391) );
  AOI22X1 U316 ( .A(RST), .B(\U_1/U_0/PLAINKEY [50]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[50] ), .Y(n392) );
  AOI22X1 U318 ( .A(RST), .B(\U_1/U_0/PLAINKEY [49]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[49] ), .Y(n393) );
  AOI22X1 U320 ( .A(RST), .B(\U_1/U_0/PLAINKEY [48]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[48] ), .Y(n394) );
  AOI22X1 U322 ( .A(RST), .B(\U_1/U_0/PLAINKEY [47]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[47] ), .Y(n395) );
  AOI22X1 U324 ( .A(RST), .B(\U_1/U_0/PLAINKEY [46]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[46] ), .Y(n396) );
  AOI22X1 U326 ( .A(RST), .B(\U_1/U_0/PLAINKEY [45]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[45] ), .Y(n397) );
  AOI22X1 U328 ( .A(RST), .B(\U_1/U_0/PLAINKEY [44]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[44] ), .Y(n398) );
  AOI22X1 U330 ( .A(RST), .B(\U_1/U_0/PLAINKEY [43]), .C(n9526), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[43] ), .Y(n399) );
  AOI22X1 U332 ( .A(RST), .B(\U_1/U_0/PLAINKEY [42]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[42] ), .Y(n400) );
  AOI22X1 U334 ( .A(RST), .B(\U_1/U_0/PLAINKEY [41]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[41] ), .Y(n401) );
  AOI22X1 U336 ( .A(RST), .B(\U_1/U_0/PLAINKEY [40]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[40] ), .Y(n402) );
  AOI22X1 U338 ( .A(RST), .B(\U_1/U_0/PLAINKEY [39]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[39] ), .Y(n403) );
  AOI22X1 U340 ( .A(RST), .B(\U_1/U_0/PLAINKEY [38]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[38] ), .Y(n404) );
  AOI22X1 U342 ( .A(RST), .B(\U_1/U_0/PLAINKEY [37]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[37] ), .Y(n405) );
  AOI22X1 U344 ( .A(RST), .B(\U_1/U_0/PLAINKEY [36]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[36] ), .Y(n406) );
  AOI22X1 U346 ( .A(RST), .B(\U_1/U_0/PLAINKEY [35]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[35] ), .Y(n407) );
  AOI22X1 U348 ( .A(RST), .B(\U_1/U_0/PLAINKEY [34]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[34] ), .Y(n408) );
  AOI22X1 U350 ( .A(RST), .B(\U_1/U_0/PLAINKEY [33]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[33] ), .Y(n409) );
  AOI22X1 U352 ( .A(RST), .B(\U_1/U_0/PLAINKEY [32]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[32] ), .Y(n410) );
  AOI22X1 U354 ( .A(RST), .B(\U_1/U_0/PLAINKEY [31]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[31] ), .Y(n411) );
  AOI22X1 U356 ( .A(RST), .B(\U_1/U_0/PLAINKEY [30]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[30] ), .Y(n412) );
  AOI22X1 U358 ( .A(RST), .B(\U_1/U_0/PLAINKEY [29]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[29] ), .Y(n413) );
  AOI22X1 U360 ( .A(RST), .B(\U_1/U_0/PLAINKEY [28]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[28] ), .Y(n414) );
  AOI22X1 U362 ( .A(RST), .B(\U_1/U_0/PLAINKEY [27]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[27] ), .Y(n415) );
  AOI22X1 U364 ( .A(RST), .B(\U_1/U_0/PLAINKEY [26]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[26] ), .Y(n416) );
  AOI22X1 U366 ( .A(RST), .B(\U_1/U_0/PLAINKEY [25]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[25] ), .Y(n417) );
  AOI22X1 U368 ( .A(RST), .B(\U_1/U_0/PLAINKEY [24]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[24] ), .Y(n418) );
  AOI22X1 U370 ( .A(RST), .B(\U_1/U_0/PLAINKEY [23]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[23] ), .Y(n419) );
  AOI22X1 U372 ( .A(RST), .B(\U_1/U_0/PLAINKEY [22]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[22] ), .Y(n420) );
  AOI22X1 U374 ( .A(RST), .B(\U_1/U_0/PLAINKEY [21]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[21] ), .Y(n421) );
  AOI22X1 U376 ( .A(RST), .B(\U_1/U_0/PLAINKEY [20]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[20] ), .Y(n422) );
  AOI22X1 U378 ( .A(RST), .B(\U_1/U_0/PLAINKEY [19]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[19] ), .Y(n423) );
  AOI22X1 U380 ( .A(RST), .B(\U_1/U_0/PLAINKEY [18]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[18] ), .Y(n424) );
  AOI22X1 U382 ( .A(RST), .B(\U_1/U_0/PLAINKEY [17]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[17] ), .Y(n425) );
  AOI22X1 U384 ( .A(RST), .B(\U_1/U_0/PLAINKEY [16]), .C(n9525), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[16] ), .Y(n426) );
  AOI22X1 U386 ( .A(RST), .B(\U_1/U_0/PLAINKEY [15]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[15] ), .Y(n427) );
  AOI22X1 U388 ( .A(RST), .B(\U_1/U_0/PLAINKEY [14]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[14] ), .Y(n428) );
  AOI22X1 U390 ( .A(RST), .B(\U_1/U_0/PLAINKEY [13]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[13] ), .Y(n429) );
  AOI22X1 U392 ( .A(RST), .B(\U_1/U_0/PLAINKEY [12]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[12] ), .Y(n430) );
  AOI22X1 U394 ( .A(RST), .B(\U_1/U_0/PLAINKEY [11]), .C(n9524), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[11] ), .Y(n431) );
  AOI22X1 U396 ( .A(RST), .B(\U_1/U_0/PLAINKEY [10]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[10] ), .Y(n432) );
  AOI22X1 U398 ( .A(RST), .B(\U_1/U_0/PLAINKEY [9]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[9] ), .Y(n433) );
  AOI22X1 U400 ( .A(RST), .B(\U_1/U_0/PLAINKEY [8]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[8] ), .Y(n434) );
  AOI22X1 U402 ( .A(RST), .B(\U_1/U_0/PLAINKEY [7]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[7] ), .Y(n435) );
  AOI22X1 U404 ( .A(RST), .B(\U_1/U_0/PLAINKEY [6]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[6] ), .Y(n436) );
  AOI22X1 U406 ( .A(RST), .B(\U_1/U_0/PLAINKEY [5]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[5] ), .Y(n437) );
  AOI22X1 U408 ( .A(RST), .B(\U_1/U_0/PLAINKEY [4]), .C(n9523), .D(
        \U_1/U_0/U_1/U_8/currentPlainKey[4] ), .Y(n438) );
  OAI22X1 U409 ( .A(n9532), .B(n11541), .C(RST), .D(n11540), .Y(n7267) );
  OAI22X1 U410 ( .A(n9533), .B(n11539), .C(RST), .D(n11538), .Y(n7268) );
  OAI22X1 U411 ( .A(n9532), .B(n11537), .C(RST), .D(n11536), .Y(n7269) );
  OAI22X1 U412 ( .A(n9532), .B(n11535), .C(RST), .D(n11534), .Y(n7270) );
  OAI22X1 U413 ( .A(\U_1/U_0/U_1/RBUF_LOAD ), .B(n9480), .C(n11524), .D(n9319), 
        .Y(n7274) );
  OAI22X1 U414 ( .A(\U_1/U_0/U_1/RBUF_LOAD ), .B(n9398), .C(n9319), .D(n11522), 
        .Y(n7277) );
  OAI22X1 U415 ( .A(\U_1/U_0/U_1/RBUF_LOAD ), .B(n9475), .C(n9319), .D(n11521), 
        .Y(n7280) );
  OAI22X1 U416 ( .A(\U_1/U_0/U_1/RBUF_LOAD ), .B(n9393), .C(n9319), .D(n11519), 
        .Y(n7283) );
  OAI22X1 U417 ( .A(\U_1/U_0/U_1/RBUF_LOAD ), .B(n11518), .C(n9319), .D(n11517), .Y(n7286) );
  OAI22X1 U418 ( .A(\U_1/U_0/U_1/RBUF_LOAD ), .B(n11516), .C(n9319), .D(n11515), .Y(n7289) );
  AOI22X1 U420 ( .A(n9319), .B(\U_1/U_0/U_1/RCV_DATA [6]), .C(
        \U_1/U_0/U_1/RBUF_LOAD ), .D(\U_1/U_0/U_1/LOAD_DATA [6]), .Y(n460) );
  OAI22X1 U421 ( .A(\U_1/U_0/U_1/RBUF_LOAD ), .B(n11513), .C(n9319), .D(n11512), .Y(n7295) );
  NAND2X1 U424 ( .A(n463), .B(n464), .Y(n7370) );
  AOI22X1 U425 ( .A(\U_0/U_3/U_3/current_send_data [7]), .B(n465), .C(
        \U_0/U_3/send_data [7]), .D(RST), .Y(n463) );
  OAI21X1 U426 ( .A(n466), .B(n11303), .C(n464), .Y(n7371) );
  AOI21X1 U427 ( .A(n468), .B(\U_0/U_3/TX_CRC [15]), .C(n10421), .Y(n464) );
  OAI21X1 U429 ( .A(n471), .B(n472), .C(n9511), .Y(n470) );
  OAI21X1 U430 ( .A(n473), .B(n11207), .C(n475), .Y(n472) );
  OAI21X1 U431 ( .A(\U_0/U_3/TX_CRC [7]), .B(\U_0/U_3/U_3/N188 ), .C(n10897), 
        .Y(n475) );
  NOR2X1 U432 ( .A(n477), .B(n11288), .Y(n471) );
  NAND2X1 U434 ( .A(n479), .B(n480), .Y(n7372) );
  AOI22X1 U435 ( .A(\U_0/U_3/U_3/current_send_data [0]), .B(n465), .C(
        \U_0/U_3/send_data [0]), .D(RST), .Y(n479) );
  OAI21X1 U436 ( .A(n466), .B(n11301), .C(n480), .Y(n7373) );
  AOI22X1 U438 ( .A(\U_0/U_3/U_3/flop_data [0]), .B(n484), .C(
        \U_0/U_3/TX_CRC [0]), .D(n485), .Y(n483) );
  AOI22X1 U439 ( .A(\U_0/PROCESSED_DATA [0]), .B(n486), .C(\U_0/U_3/TX_CRC [8]), .D(n468), .Y(n482) );
  NAND2X1 U441 ( .A(n487), .B(n488), .Y(n7374) );
  AOI22X1 U442 ( .A(\U_0/U_3/U_3/current_send_data [1]), .B(n465), .C(
        \U_0/U_3/send_data [1]), .D(RST), .Y(n487) );
  OAI21X1 U443 ( .A(n466), .B(n11299), .C(n488), .Y(n7375) );
  AOI22X1 U445 ( .A(\U_0/U_3/U_3/flop_data [1]), .B(n484), .C(
        \U_0/U_3/TX_CRC [1]), .D(n485), .Y(n491) );
  AOI22X1 U446 ( .A(\U_0/PROCESSED_DATA [1]), .B(n486), .C(\U_0/U_3/TX_CRC [9]), .D(n468), .Y(n490) );
  NAND2X1 U448 ( .A(n492), .B(n493), .Y(n7376) );
  AOI22X1 U449 ( .A(\U_0/U_3/U_3/current_send_data [2]), .B(n465), .C(
        \U_0/U_3/send_data [2]), .D(RST), .Y(n492) );
  OAI21X1 U450 ( .A(n466), .B(n11297), .C(n493), .Y(n7377) );
  AOI22X1 U452 ( .A(\U_0/U_3/U_3/flop_data [2]), .B(n484), .C(
        \U_0/U_3/TX_CRC [2]), .D(n485), .Y(n496) );
  AOI22X1 U453 ( .A(\U_0/PROCESSED_DATA [2]), .B(n486), .C(
        \U_0/U_3/TX_CRC [10]), .D(n468), .Y(n495) );
  NAND2X1 U455 ( .A(n497), .B(n498), .Y(n7378) );
  AOI22X1 U456 ( .A(\U_0/U_3/U_3/current_send_data [3]), .B(n465), .C(
        \U_0/U_3/send_data [3]), .D(RST), .Y(n497) );
  OAI21X1 U457 ( .A(n466), .B(n11295), .C(n498), .Y(n7379) );
  AOI22X1 U459 ( .A(\U_0/U_3/U_3/flop_data [3]), .B(n484), .C(
        \U_0/U_3/TX_CRC [3]), .D(n485), .Y(n501) );
  AOI22X1 U460 ( .A(\U_0/PROCESSED_DATA [3]), .B(n486), .C(
        \U_0/U_3/TX_CRC [11]), .D(n468), .Y(n500) );
  NAND2X1 U462 ( .A(n502), .B(n503), .Y(n7380) );
  AOI22X1 U463 ( .A(\U_0/U_3/U_3/current_send_data [4]), .B(n465), .C(
        \U_0/U_3/send_data [4]), .D(RST), .Y(n502) );
  OAI21X1 U464 ( .A(n466), .B(n11293), .C(n503), .Y(n7381) );
  AOI22X1 U466 ( .A(\U_0/U_3/U_3/flop_data [4]), .B(n484), .C(
        \U_0/U_3/TX_CRC [4]), .D(n485), .Y(n506) );
  AOI22X1 U467 ( .A(\U_0/PROCESSED_DATA [4]), .B(n486), .C(
        \U_0/U_3/TX_CRC [12]), .D(n468), .Y(n505) );
  NAND2X1 U469 ( .A(n507), .B(n508), .Y(n7382) );
  AOI22X1 U470 ( .A(\U_0/U_3/U_3/current_send_data [5]), .B(n465), .C(
        \U_0/U_3/send_data [5]), .D(RST), .Y(n507) );
  OAI21X1 U471 ( .A(n466), .B(n11291), .C(n508), .Y(n7383) );
  AOI22X1 U473 ( .A(\U_0/U_3/U_3/flop_data [5]), .B(n484), .C(
        \U_0/U_3/TX_CRC [5]), .D(n485), .Y(n511) );
  AOI22X1 U474 ( .A(\U_0/PROCESSED_DATA [5]), .B(n486), .C(
        \U_0/U_3/TX_CRC [13]), .D(n468), .Y(n510) );
  NAND2X1 U476 ( .A(n512), .B(n513), .Y(n7384) );
  AOI22X1 U477 ( .A(\U_0/U_3/U_3/current_send_data [6]), .B(n465), .C(
        \U_0/U_3/send_data [6]), .D(RST), .Y(n512) );
  OAI21X1 U479 ( .A(n466), .B(n11289), .C(n513), .Y(n7385) );
  AOI22X1 U481 ( .A(\U_0/U_3/U_3/flop_data [6]), .B(n484), .C(
        \U_0/U_3/TX_CRC [6]), .D(n485), .Y(n517) );
  NOR3X1 U482 ( .A(RST), .B(\U_0/U_3/U_3/N188 ), .C(n518), .Y(n485) );
  NOR2X1 U483 ( .A(n477), .B(RST), .Y(n484) );
  AOI22X1 U484 ( .A(\U_0/PROCESSED_DATA [6]), .B(n486), .C(
        \U_0/U_3/TX_CRC [14]), .D(n468), .Y(n516) );
  NOR2X1 U485 ( .A(n519), .B(RST), .Y(n468) );
  NOR2X1 U486 ( .A(n473), .B(RST), .Y(n486) );
  NOR2X1 U488 ( .A(n514), .B(RST), .Y(n466) );
  OAI21X1 U489 ( .A(n10904), .B(n10900), .C(n522), .Y(n514) );
  OAI22X1 U490 ( .A(n523), .B(n11088), .C(n525), .D(n11287), .Y(n7386) );
  OAI21X1 U492 ( .A(RST), .B(n10544), .C(n528), .Y(n7387) );
  NAND2X1 U493 ( .A(DATA_H[7]), .B(RST), .Y(n528) );
  OAI22X1 U494 ( .A(n9532), .B(n11254), .C(RST), .D(n10544), .Y(n7388) );
  AOI22X1 U497 ( .A(RST), .B(\U_0/U_0/U_0/faddr [7]), .C(n9523), .D(
        \U_0/U_0/U_0/nfaddr[7] ), .Y(n530) );
  OAI21X1 U498 ( .A(RST), .B(n11128), .C(n532), .Y(n7390) );
  NAND2X1 U499 ( .A(ADDR_H[7]), .B(RST), .Y(n532) );
  AOI22X1 U502 ( .A(RST), .B(\U_0/U_0/U_0/faddr [6]), .C(n9523), .D(
        \U_0/U_0/U_0/nfaddr[6] ), .Y(n533) );
  OAI21X1 U503 ( .A(RST), .B(n11127), .C(n535), .Y(n7392) );
  NAND2X1 U504 ( .A(ADDR_H[6]), .B(RST), .Y(n535) );
  AOI22X1 U507 ( .A(RST), .B(\U_0/U_0/U_0/faddr [5]), .C(n9523), .D(
        \U_0/U_0/U_0/nfaddr[5] ), .Y(n536) );
  OAI21X1 U508 ( .A(RST), .B(n11126), .C(n538), .Y(n7394) );
  NAND2X1 U509 ( .A(ADDR_H[5]), .B(RST), .Y(n538) );
  AOI22X1 U512 ( .A(RST), .B(\U_0/U_0/U_0/faddr [4]), .C(n9523), .D(
        \U_0/U_0/U_0/nfaddr[4] ), .Y(n539) );
  OAI21X1 U513 ( .A(RST), .B(n11125), .C(n541), .Y(n7396) );
  NAND2X1 U514 ( .A(ADDR_H[4]), .B(RST), .Y(n541) );
  AOI22X1 U517 ( .A(RST), .B(\U_0/U_0/U_0/faddr [3]), .C(n9523), .D(
        \U_0/U_0/U_0/nfaddr[3] ), .Y(n542) );
  OAI21X1 U518 ( .A(RST), .B(n11124), .C(n544), .Y(n7398) );
  NAND2X1 U519 ( .A(ADDR_H[3]), .B(RST), .Y(n544) );
  AOI22X1 U522 ( .A(RST), .B(\U_0/U_0/U_0/faddr [2]), .C(n9524), .D(
        \U_0/U_0/U_0/nfaddr[2] ), .Y(n545) );
  OAI21X1 U523 ( .A(RST), .B(n11123), .C(n547), .Y(n7400) );
  NAND2X1 U524 ( .A(ADDR_H[2]), .B(RST), .Y(n547) );
  AOI22X1 U527 ( .A(RST), .B(\U_0/U_0/U_0/faddr [1]), .C(n9523), .D(
        \U_0/U_0/U_0/nfaddr[1] ), .Y(n548) );
  OAI21X1 U528 ( .A(RST), .B(n11122), .C(n550), .Y(n7402) );
  NAND2X1 U529 ( .A(ADDR_H[1]), .B(RST), .Y(n550) );
  AOI22X1 U532 ( .A(RST), .B(\U_0/U_0/U_0/faddr [0]), .C(n9522), .D(
        \U_0/U_0/U_0/nfaddr[0] ), .Y(n551) );
  OAI21X1 U533 ( .A(RST), .B(n11121), .C(n553), .Y(n7404) );
  NAND2X1 U534 ( .A(ADDR_H[0]), .B(RST), .Y(n553) );
  OAI21X1 U536 ( .A(RST), .B(n554), .C(n555), .Y(n7413) );
  NAND2X1 U537 ( .A(R_ENABLE_H), .B(RST), .Y(n555) );
  AOI21X1 U538 ( .A(\U_0/U_0/U_0/fr_enable ), .B(n556), .C(n557), .Y(n554) );
  OAI21X1 U539 ( .A(RST), .B(n11135), .C(n559), .Y(n7414) );
  OAI21X1 U540 ( .A(RST), .B(n556), .C(\U_0/U_0/U_0/fr_enable ), .Y(n559) );
  NAND3X1 U542 ( .A(n562), .B(n11153), .C(n11141), .Y(n561) );
  NAND3X1 U543 ( .A(n11155), .B(n566), .C(n567), .Y(n560) );
  NAND2X1 U545 ( .A(n568), .B(n569), .Y(n557) );
  OAI21X1 U546 ( .A(RST), .B(n10551), .C(n571), .Y(n7415) );
  NAND2X1 U547 ( .A(DATA_H[0]), .B(RST), .Y(n571) );
  OAI22X1 U548 ( .A(n9532), .B(n11240), .C(RST), .D(n10551), .Y(n7416) );
  OAI21X1 U550 ( .A(RST), .B(n10550), .C(n574), .Y(n7417) );
  NAND2X1 U551 ( .A(DATA_H[1]), .B(RST), .Y(n574) );
  OAI22X1 U552 ( .A(n9532), .B(n11239), .C(RST), .D(n10550), .Y(n7418) );
  OAI21X1 U554 ( .A(RST), .B(n10549), .C(n577), .Y(n7419) );
  NAND2X1 U555 ( .A(DATA_H[2]), .B(RST), .Y(n577) );
  OAI22X1 U556 ( .A(n9533), .B(n11238), .C(RST), .D(n10549), .Y(n7420) );
  OAI21X1 U558 ( .A(RST), .B(n10548), .C(n580), .Y(n7421) );
  NAND2X1 U559 ( .A(DATA_H[3]), .B(RST), .Y(n580) );
  OAI22X1 U560 ( .A(n9533), .B(n11237), .C(RST), .D(n10548), .Y(n7422) );
  OAI21X1 U562 ( .A(RST), .B(n10547), .C(n583), .Y(n7423) );
  NAND2X1 U563 ( .A(DATA_H[4]), .B(RST), .Y(n583) );
  OAI22X1 U564 ( .A(n9533), .B(n11236), .C(RST), .D(n10547), .Y(n7424) );
  OAI21X1 U566 ( .A(RST), .B(n10546), .C(n586), .Y(n7425) );
  NAND2X1 U567 ( .A(DATA_H[5]), .B(RST), .Y(n586) );
  OAI22X1 U568 ( .A(n9533), .B(n11235), .C(RST), .D(n10546), .Y(n7426) );
  OAI21X1 U570 ( .A(RST), .B(n10545), .C(n589), .Y(n7427) );
  NAND2X1 U571 ( .A(DATA_H[6]), .B(RST), .Y(n589) );
  OAI22X1 U572 ( .A(n9532), .B(n11234), .C(RST), .D(n10545), .Y(n7428) );
  AOI22X1 U575 ( .A(RST), .B(\U_0/PROCESSED_DATA [0]), .C(n9525), .D(
        \U_0/U_0/U_0/nextProcessedData[0] ), .Y(n591) );
  AOI22X1 U577 ( .A(RST), .B(\U_0/PROCESSED_DATA [1]), .C(n9529), .D(
        \U_0/U_0/U_0/nextProcessedData[1] ), .Y(n592) );
  AOI22X1 U579 ( .A(RST), .B(\U_0/PROCESSED_DATA [2]), .C(n9530), .D(
        \U_0/U_0/U_0/nextProcessedData[2] ), .Y(n593) );
  AOI22X1 U581 ( .A(RST), .B(\U_0/PROCESSED_DATA [3]), .C(n9528), .D(
        \U_0/U_0/U_0/nextProcessedData[3] ), .Y(n594) );
  AOI22X1 U583 ( .A(RST), .B(\U_0/PROCESSED_DATA [4]), .C(n9528), .D(
        \U_0/U_0/U_0/nextProcessedData[4] ), .Y(n595) );
  AOI22X1 U585 ( .A(RST), .B(\U_0/PROCESSED_DATA [5]), .C(n9528), .D(
        \U_0/U_0/U_0/nextProcessedData[5] ), .Y(n596) );
  AOI22X1 U587 ( .A(RST), .B(\U_0/PROCESSED_DATA [6]), .C(n9528), .D(
        \U_0/U_0/U_0/nextProcessedData[6] ), .Y(n597) );
  AOI22X1 U589 ( .A(RST), .B(\U_0/PROCESSED_DATA [7]), .C(n9528), .D(
        \U_0/U_0/U_0/nextProcessedData[7] ), .Y(n598) );
  OAI21X1 U590 ( .A(RST), .B(n599), .C(n600), .Y(n7461) );
  NAND2X1 U591 ( .A(W_ENABLE_H), .B(RST), .Y(n600) );
  AOI21X1 U592 ( .A(\U_0/U_0/U_0/fw_enable ), .B(n601), .C(n602), .Y(n599) );
  OAI21X1 U593 ( .A(RST), .B(n11140), .C(n604), .Y(n7462) );
  OAI21X1 U594 ( .A(RST), .B(n601), .C(\U_0/U_0/U_0/fw_enable ), .Y(n604) );
  NAND2X1 U595 ( .A(n11130), .B(n562), .Y(n601) );
  NAND3X1 U597 ( .A(n11160), .B(n567), .C(n607), .Y(n602) );
  OAI21X1 U598 ( .A(n9534), .B(n11113), .C(n609), .Y(n7483) );
  AOI22X1 U599 ( .A(n610), .B(\U_0/U_1/U_0/tempOpcode [1]), .C(
        \U_0/U_1/OUT_OPCODE [1]), .D(n10510), .Y(n609) );
  OAI21X1 U600 ( .A(n9534), .B(n11112), .C(n613), .Y(n7484) );
  AOI22X1 U601 ( .A(\U_0/U_1/U_0/tempData [0]), .B(n610), .C(\U_0/U_1/DATA [0]), .D(n10510), .Y(n613) );
  OAI22X1 U603 ( .A(n523), .B(n11079), .C(n525), .D(n11111), .Y(n7485) );
  OAI21X1 U605 ( .A(n9534), .B(n11110), .C(n617), .Y(n7486) );
  AOI22X1 U606 ( .A(\U_0/U_1/U_0/tempData [1]), .B(n610), .C(\U_0/U_1/DATA [1]), .D(n10510), .Y(n617) );
  OAI22X1 U608 ( .A(n523), .B(n11080), .C(n525), .D(n11109), .Y(n7487) );
  OAI21X1 U610 ( .A(n9533), .B(n11108), .C(n621), .Y(n7488) );
  AOI22X1 U611 ( .A(\U_0/U_1/U_0/tempData [2]), .B(n610), .C(\U_0/U_1/DATA [2]), .D(n10510), .Y(n621) );
  OAI22X1 U613 ( .A(n523), .B(n11081), .C(n525), .D(n11107), .Y(n7489) );
  OAI21X1 U615 ( .A(n9533), .B(n11106), .C(n625), .Y(n7490) );
  AOI22X1 U616 ( .A(\U_0/U_1/U_0/tempData [3]), .B(n610), .C(\U_0/U_1/DATA [3]), .D(n10510), .Y(n625) );
  OAI22X1 U618 ( .A(n523), .B(n11082), .C(n525), .D(n11105), .Y(n7491) );
  OAI21X1 U620 ( .A(n9533), .B(n11104), .C(n629), .Y(n7492) );
  AOI22X1 U621 ( .A(\U_0/U_1/U_0/tempData [4]), .B(n610), .C(\U_0/U_1/DATA [4]), .D(n10510), .Y(n629) );
  OAI22X1 U623 ( .A(n523), .B(n11083), .C(n525), .D(n11103), .Y(n7493) );
  OAI21X1 U625 ( .A(n9533), .B(n11102), .C(n633), .Y(n7494) );
  AOI22X1 U626 ( .A(\U_0/U_1/U_0/tempData [5]), .B(n610), .C(\U_0/U_1/DATA [5]), .D(n10510), .Y(n633) );
  OAI22X1 U628 ( .A(n523), .B(n11084), .C(n525), .D(n11101), .Y(n7495) );
  OAI21X1 U630 ( .A(n9534), .B(n11100), .C(n637), .Y(n7496) );
  AOI22X1 U631 ( .A(\U_0/U_1/U_0/tempData [6]), .B(n610), .C(\U_0/U_1/DATA [6]), .D(n10510), .Y(n637) );
  OAI22X1 U633 ( .A(n523), .B(n11085), .C(n525), .D(n11099), .Y(n7497) );
  OAI21X1 U635 ( .A(n9533), .B(n11098), .C(n641), .Y(n7498) );
  AOI22X1 U636 ( .A(\U_0/U_1/U_0/tempData [7]), .B(n610), .C(\U_0/U_1/DATA [7]), .D(n10510), .Y(n641) );
  OAI22X1 U638 ( .A(n523), .B(n11086), .C(n525), .D(n11097), .Y(n7499) );
  OAI22X1 U640 ( .A(n523), .B(n11087), .C(n525), .D(n11096), .Y(n7500) );
  NOR2X1 U642 ( .A(n646), .B(RST), .Y(n525) );
  OAI21X1 U643 ( .A(n9533), .B(n11095), .C(n648), .Y(n7501) );
  AOI22X1 U644 ( .A(\U_0/U_1/U_0/tempOpcode [0]), .B(n610), .C(
        \U_0/U_1/OUT_OPCODE [0]), .D(n10510), .Y(n648) );
  NAND2X1 U647 ( .A(\U_0/U_1/U_0/state[2] ), .B(n11089), .Y(n646) );
  OAI21X1 U648 ( .A(n9533), .B(n11092), .C(n523), .Y(n7502) );
  NAND3X1 U649 ( .A(n11090), .B(n11091), .C(n653), .Y(n523) );
  NOR2X1 U650 ( .A(RST), .B(n10905), .Y(n653) );
  AOI22X1 U652 ( .A(EMPTY_H), .B(RST), .C(\U_0/U_1/U_1/N349 ), .D(n9522), .Y(
        n655) );
  AOI22X1 U654 ( .A(FULL_H), .B(RST), .C(\U_0/U_1/U_1/N355 ), .D(n9522), .Y(
        n656) );
  OAI21X1 U655 ( .A(n9533), .B(n10908), .C(n658), .Y(n7522) );
  NAND3X1 U656 ( .A(n11091), .B(n10905), .C(n659), .Y(n658) );
  NOR2X1 U657 ( .A(RST), .B(n11090), .Y(n659) );
  OAI22X1 U659 ( .A(n9532), .B(n10880), .C(RST), .D(n10879), .Y(n7532) );
  OAI22X1 U661 ( .A(n9532), .B(n10791), .C(RST), .D(n10790), .Y(n7599) );
  AOI22X1 U664 ( .A(RST), .B(\U_0/U_0/PLAINKEY [62]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[62] ), .Y(n664) );
  AOI22X1 U666 ( .A(RST), .B(\U_0/U_0/PLAINKEY [61]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[61] ), .Y(n665) );
  AOI22X1 U668 ( .A(RST), .B(\U_0/U_0/PLAINKEY [60]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[60] ), .Y(n666) );
  AOI22X1 U670 ( .A(RST), .B(\U_0/U_0/PLAINKEY [59]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[59] ), .Y(n667) );
  AOI22X1 U672 ( .A(RST), .B(\U_0/U_0/PLAINKEY [58]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[58] ), .Y(n668) );
  AOI22X1 U674 ( .A(RST), .B(\U_0/U_0/PLAINKEY [57]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[57] ), .Y(n669) );
  AOI22X1 U676 ( .A(RST), .B(\U_0/U_0/PLAINKEY [56]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[56] ), .Y(n670) );
  AOI22X1 U678 ( .A(RST), .B(\U_0/U_0/PLAINKEY [55]), .C(n9525), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[55] ), .Y(n671) );
  AOI22X1 U680 ( .A(RST), .B(\U_0/U_0/PLAINKEY [54]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[54] ), .Y(n672) );
  AOI22X1 U682 ( .A(RST), .B(\U_0/U_0/PLAINKEY [53]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[53] ), .Y(n673) );
  AOI22X1 U684 ( .A(RST), .B(\U_0/U_0/PLAINKEY [52]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[52] ), .Y(n674) );
  AOI22X1 U686 ( .A(RST), .B(\U_0/U_0/PLAINKEY [51]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[51] ), .Y(n675) );
  AOI22X1 U688 ( .A(RST), .B(\U_0/U_0/PLAINKEY [50]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[50] ), .Y(n676) );
  AOI22X1 U690 ( .A(RST), .B(\U_0/U_0/PLAINKEY [49]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[49] ), .Y(n677) );
  AOI22X1 U692 ( .A(RST), .B(\U_0/U_0/PLAINKEY [48]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[48] ), .Y(n678) );
  AOI22X1 U694 ( .A(RST), .B(\U_0/U_0/PLAINKEY [47]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[47] ), .Y(n679) );
  AOI22X1 U696 ( .A(RST), .B(\U_0/U_0/PLAINKEY [46]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[46] ), .Y(n680) );
  AOI22X1 U698 ( .A(RST), .B(\U_0/U_0/PLAINKEY [45]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[45] ), .Y(n681) );
  AOI22X1 U700 ( .A(RST), .B(\U_0/U_0/PLAINKEY [44]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[44] ), .Y(n682) );
  AOI22X1 U702 ( .A(RST), .B(\U_0/U_0/PLAINKEY [43]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[43] ), .Y(n683) );
  AOI22X1 U704 ( .A(RST), .B(\U_0/U_0/PLAINKEY [42]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[42] ), .Y(n684) );
  AOI22X1 U706 ( .A(RST), .B(\U_0/U_0/PLAINKEY [41]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[41] ), .Y(n685) );
  AOI22X1 U708 ( .A(RST), .B(\U_0/U_0/PLAINKEY [40]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[40] ), .Y(n686) );
  AOI22X1 U710 ( .A(RST), .B(\U_0/U_0/PLAINKEY [39]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[39] ), .Y(n687) );
  AOI22X1 U712 ( .A(RST), .B(\U_0/U_0/PLAINKEY [38]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[38] ), .Y(n688) );
  AOI22X1 U714 ( .A(RST), .B(\U_0/U_0/PLAINKEY [37]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[37] ), .Y(n689) );
  AOI22X1 U716 ( .A(RST), .B(\U_0/U_0/PLAINKEY [36]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[36] ), .Y(n690) );
  AOI22X1 U718 ( .A(RST), .B(\U_0/U_0/PLAINKEY [35]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[35] ), .Y(n691) );
  AOI22X1 U720 ( .A(RST), .B(\U_0/U_0/PLAINKEY [34]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[34] ), .Y(n692) );
  AOI22X1 U722 ( .A(RST), .B(\U_0/U_0/PLAINKEY [33]), .C(n9530), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[33] ), .Y(n693) );
  AOI22X1 U724 ( .A(RST), .B(\U_0/U_0/PLAINKEY [32]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[32] ), .Y(n694) );
  AOI22X1 U726 ( .A(RST), .B(\U_0/U_0/PLAINKEY [31]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[31] ), .Y(n695) );
  AOI22X1 U728 ( .A(RST), .B(\U_0/U_0/PLAINKEY [30]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[30] ), .Y(n696) );
  AOI22X1 U730 ( .A(RST), .B(\U_0/U_0/PLAINKEY [29]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[29] ), .Y(n697) );
  AOI22X1 U732 ( .A(RST), .B(\U_0/U_0/PLAINKEY [28]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[28] ), .Y(n698) );
  AOI22X1 U734 ( .A(RST), .B(\U_0/U_0/PLAINKEY [27]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[27] ), .Y(n699) );
  AOI22X1 U736 ( .A(RST), .B(\U_0/U_0/PLAINKEY [26]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[26] ), .Y(n700) );
  AOI22X1 U738 ( .A(RST), .B(\U_0/U_0/PLAINKEY [25]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[25] ), .Y(n701) );
  AOI22X1 U740 ( .A(RST), .B(\U_0/U_0/PLAINKEY [24]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[24] ), .Y(n702) );
  AOI22X1 U742 ( .A(RST), .B(\U_0/U_0/PLAINKEY [23]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[23] ), .Y(n703) );
  AOI22X1 U744 ( .A(RST), .B(\U_0/U_0/PLAINKEY [22]), .C(n9531), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[22] ), .Y(n704) );
  AOI22X1 U746 ( .A(RST), .B(\U_0/U_0/PLAINKEY [21]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[21] ), .Y(n705) );
  AOI22X1 U748 ( .A(RST), .B(\U_0/U_0/PLAINKEY [20]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[20] ), .Y(n706) );
  AOI22X1 U750 ( .A(RST), .B(\U_0/U_0/PLAINKEY [19]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[19] ), .Y(n707) );
  AOI22X1 U752 ( .A(RST), .B(\U_0/U_0/PLAINKEY [18]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[18] ), .Y(n708) );
  AOI22X1 U754 ( .A(RST), .B(\U_0/U_0/PLAINKEY [17]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[17] ), .Y(n709) );
  AOI22X1 U756 ( .A(RST), .B(\U_0/U_0/PLAINKEY [16]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[16] ), .Y(n710) );
  AOI22X1 U758 ( .A(RST), .B(\U_0/U_0/PLAINKEY [15]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[15] ), .Y(n711) );
  AOI22X1 U760 ( .A(RST), .B(\U_0/U_0/PLAINKEY [14]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[14] ), .Y(n712) );
  AOI22X1 U762 ( .A(RST), .B(\U_0/U_0/PLAINKEY [13]), .C(n9529), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[13] ), .Y(n713) );
  AOI22X1 U764 ( .A(RST), .B(\U_0/U_0/PLAINKEY [12]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[12] ), .Y(n714) );
  AOI22X1 U766 ( .A(RST), .B(\U_0/U_0/PLAINKEY [11]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[11] ), .Y(n715) );
  AOI22X1 U768 ( .A(RST), .B(\U_0/U_0/PLAINKEY [10]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[10] ), .Y(n716) );
  AOI22X1 U770 ( .A(RST), .B(\U_0/U_0/PLAINKEY [9]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[9] ), .Y(n717) );
  AOI22X1 U772 ( .A(RST), .B(\U_0/U_0/PLAINKEY [8]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[8] ), .Y(n718) );
  AOI22X1 U774 ( .A(RST), .B(\U_0/U_0/PLAINKEY [7]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[7] ), .Y(n719) );
  AOI22X1 U776 ( .A(RST), .B(\U_0/U_0/PLAINKEY [6]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[6] ), .Y(n720) );
  AOI22X1 U778 ( .A(RST), .B(\U_0/U_0/PLAINKEY [5]), .C(n9528), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[5] ), .Y(n721) );
  AOI22X1 U780 ( .A(RST), .B(\U_0/U_0/PLAINKEY [4]), .C(n9508), .D(
        \U_0/U_0/U_1/U_8/currentPlainKey[4] ), .Y(n722) );
  OAI22X1 U781 ( .A(n9532), .B(n10789), .C(RST), .D(n10788), .Y(n7659) );
  OAI22X1 U782 ( .A(n9532), .B(n10787), .C(RST), .D(n10786), .Y(n7660) );
  OAI22X1 U783 ( .A(n9532), .B(n10785), .C(RST), .D(n10784), .Y(n7661) );
  OAI22X1 U784 ( .A(n9532), .B(n10783), .C(RST), .D(n10782), .Y(n7662) );
  OAI22X1 U785 ( .A(\U_0/U_0/U_1/RBUF_LOAD ), .B(n9487), .C(n10772), .D(n9354), 
        .Y(n7666) );
  OAI22X1 U786 ( .A(\U_0/U_0/U_1/RBUF_LOAD ), .B(n9388), .C(n9354), .D(n10770), 
        .Y(n7669) );
  OAI22X1 U787 ( .A(\U_0/U_0/U_1/RBUF_LOAD ), .B(n9482), .C(n9354), .D(n10769), 
        .Y(n7672) );
  OAI22X1 U788 ( .A(\U_0/U_0/U_1/RBUF_LOAD ), .B(n9383), .C(n9354), .D(n10767), 
        .Y(n7675) );
  OAI22X1 U789 ( .A(\U_0/U_0/U_1/RBUF_LOAD ), .B(n10766), .C(n9354), .D(n10765), .Y(n7678) );
  OAI22X1 U790 ( .A(\U_0/U_0/U_1/RBUF_LOAD ), .B(n10764), .C(n9354), .D(n10763), .Y(n7681) );
  AOI22X1 U792 ( .A(n9354), .B(\U_0/U_0/U_1/RCV_DATA [6]), .C(
        \U_0/U_0/U_1/RBUF_LOAD ), .D(\U_0/U_0/U_1/LOAD_DATA [6]), .Y(n744) );
  OAI22X1 U793 ( .A(\U_0/U_0/U_1/RBUF_LOAD ), .B(n10761), .C(n9354), .D(n10760), .Y(n7687) );
  OAI21X1 U798 ( .A(n749), .B(n750), .C(n9690), .Y(n748) );
  OAI21X1 U799 ( .A(n9710), .B(n753), .C(n754), .Y(n750) );
  OAI21X1 U800 ( .A(n9705), .B(n756), .C(n757), .Y(n749) );
  NAND3X1 U801 ( .A(\U_0/U_2/U_1/state[1] ), .B(n758), .C(n10810), .Y(n757) );
  OAI21X1 U805 ( .A(n763), .B(n764), .C(n9698), .Y(n762) );
  OAI21X1 U806 ( .A(n9716), .B(n767), .C(n768), .Y(n764) );
  OAI21X1 U807 ( .A(n9708), .B(n770), .C(n771), .Y(n763) );
  NAND3X1 U808 ( .A(\U_1/U_2/U_1/state[1] ), .B(n772), .C(n11562), .Y(n771) );
  OAI22X1 U810 ( .A(n11207), .B(n10051), .C(n9239), .D(n11288), .Y(n7750) );
  OAI22X1 U813 ( .A(n12035), .B(n777), .C(n9281), .D(n12054), .Y(n7751) );
  OAI22X1 U816 ( .A(n11620), .B(n12077), .C(n11631), .D(n781), .Y(n7757) );
  NAND3X1 U818 ( .A(\U_1/U_3/U_0/N59 ), .B(n11627), .C(n783), .Y(n781) );
  NOR2X1 U819 ( .A(n784), .B(n785), .Y(n783) );
  AOI22X1 U821 ( .A(\U_1/U_3/send_data [7]), .B(n11641), .C(n788), .D(
        \U_1/U_3/U_2/present_val [7]), .Y(n786) );
  OAI21X1 U822 ( .A(n12056), .B(n790), .C(n791), .Y(n7759) );
  AOI22X1 U823 ( .A(n9285), .B(\U_1/U_3/U_2/present_val [7]), .C(
        \U_1/U_3/U_2/present_val [6]), .D(n788), .Y(n791) );
  OAI21X1 U825 ( .A(n12058), .B(n790), .C(n794), .Y(n7760) );
  AOI22X1 U826 ( .A(\U_1/U_3/U_2/present_val [6]), .B(n9285), .C(
        \U_1/U_3/U_2/present_val [5]), .D(n788), .Y(n794) );
  OAI21X1 U828 ( .A(n12060), .B(n790), .C(n796), .Y(n7761) );
  AOI22X1 U829 ( .A(\U_1/U_3/U_2/present_val [5]), .B(n9285), .C(
        \U_1/U_3/U_2/present_val [4]), .D(n788), .Y(n796) );
  OAI21X1 U831 ( .A(n12062), .B(n790), .C(n798), .Y(n7762) );
  AOI22X1 U832 ( .A(\U_1/U_3/U_2/present_val [4]), .B(n9285), .C(
        \U_1/U_3/U_2/present_val [3]), .D(n788), .Y(n798) );
  OAI21X1 U834 ( .A(n12064), .B(n790), .C(n800), .Y(n7763) );
  AOI22X1 U835 ( .A(\U_1/U_3/U_2/present_val [3]), .B(n9285), .C(
        \U_1/U_3/U_2/present_val [2]), .D(n788), .Y(n800) );
  OAI21X1 U837 ( .A(n12066), .B(n790), .C(n802), .Y(n7764) );
  AOI22X1 U838 ( .A(\U_1/U_3/U_2/present_val [2]), .B(n9285), .C(
        \U_1/U_3/U_2/present_val [1]), .D(n788), .Y(n802) );
  OAI21X1 U840 ( .A(n12068), .B(n790), .C(n804), .Y(n7765) );
  AOI22X1 U841 ( .A(\U_1/U_3/U_2/present_val [1]), .B(n9285), .C(
        \U_1/U_3/d_encode ), .D(n788), .Y(n804) );
  OAI21X1 U843 ( .A(n11641), .B(n12074), .C(n806), .Y(n7766) );
  NAND3X1 U844 ( .A(\U_1/U_3/U_2/count[1] ), .B(\U_1/U_3/U_2/count[0] ), .C(
        n9285), .Y(n806) );
  OAI21X1 U845 ( .A(n11624), .B(n808), .C(n809), .Y(n7767) );
  OAI21X1 U846 ( .A(n788), .B(n12075), .C(\U_1/U_3/U_2/count[1] ), .Y(n809) );
  NAND2X1 U847 ( .A(\U_1/U_3/U_2/count[0] ), .B(n12073), .Y(n808) );
  AOI22X1 U850 ( .A(\U_1/U_3/U_2/count[0] ), .B(n788), .C(n12075), .D(n9285), 
        .Y(n812) );
  NOR2X1 U851 ( .A(n11641), .B(n788), .Y(n792) );
  AOI21X1 U853 ( .A(\U_1/U_3/U_0/N59 ), .B(n7756), .C(n11641), .Y(n788) );
  NAND3X1 U855 ( .A(\U_1/U_3/U_2/count[0] ), .B(n7756), .C(n813), .Y(n790) );
  NOR2X1 U856 ( .A(n12073), .B(n12074), .Y(n813) );
  NOR2X1 U859 ( .A(n814), .B(n815), .Y(n7756) );
  NAND3X1 U860 ( .A(\U_1/U_3/U_4/count[3] ), .B(slave_is_sending), .C(
        \U_1/U_3/U_4/state ), .Y(n815) );
  OAI22X1 U861 ( .A(n12049), .B(n9284), .C(n818), .D(n9283), .Y(n7769) );
  XNOR2X1 U862 ( .A(n820), .B(n12048), .Y(n818) );
  OAI22X1 U864 ( .A(n12046), .B(n9283), .C(n12047), .D(n9284), .Y(n7770) );
  OAI22X1 U866 ( .A(n12044), .B(n9283), .C(n12045), .D(n9284), .Y(n7771) );
  OAI22X1 U868 ( .A(n12042), .B(n9283), .C(n12043), .D(n9284), .Y(n7772) );
  OAI22X1 U870 ( .A(n12040), .B(n9283), .C(n12041), .D(n9284), .Y(n7773) );
  OAI22X1 U871 ( .A(n12038), .B(n9283), .C(n12039), .D(n9284), .Y(n7774) );
  OAI22X1 U873 ( .A(n12051), .B(n9284), .C(n833), .D(n9283), .Y(n7775) );
  XNOR2X1 U874 ( .A(\U_1/U_3/TX_CRC [1]), .B(n834), .Y(n833) );
  OAI22X1 U876 ( .A(n12037), .B(n9284), .C(n836), .D(n9283), .Y(n7776) );
  XOR2X1 U877 ( .A(n837), .B(n838), .Y(n836) );
  XNOR2X1 U878 ( .A(\U_1/U_3/TX_CRC [0]), .B(n834), .Y(n837) );
  OAI22X1 U879 ( .A(n12048), .B(n9284), .C(n839), .D(n9283), .Y(n7777) );
  OAI22X1 U881 ( .A(n12046), .B(n9284), .C(n840), .D(n819), .Y(n7778) );
  XNOR2X1 U882 ( .A(n841), .B(n842), .Y(n840) );
  OAI22X1 U884 ( .A(n12044), .B(n9284), .C(n843), .D(n819), .Y(n7779) );
  OAI22X1 U886 ( .A(n12042), .B(n9284), .C(n844), .D(n819), .Y(n7780) );
  XNOR2X1 U887 ( .A(n845), .B(n846), .Y(n844) );
  OAI22X1 U889 ( .A(n12040), .B(n9284), .C(n847), .D(n819), .Y(n7781) );
  OAI22X1 U891 ( .A(n12038), .B(n9284), .C(n848), .D(n819), .Y(n7782) );
  XOR2X1 U892 ( .A(n849), .B(n850), .Y(n848) );
  OAI22X1 U894 ( .A(n12050), .B(n9284), .C(n852), .D(n819), .Y(n7783) );
  XNOR2X1 U895 ( .A(n853), .B(n839), .Y(n852) );
  XNOR2X1 U896 ( .A(n834), .B(n854), .Y(n853) );
  OAI22X1 U898 ( .A(n12036), .B(n9284), .C(n820), .D(n819), .Y(n7784) );
  XOR2X1 U899 ( .A(n856), .B(n857), .Y(n820) );
  XOR2X1 U900 ( .A(n834), .B(n850), .Y(n857) );
  XNOR2X1 U901 ( .A(n12037), .B(\U_1/PROCESSED_DATA [0]), .Y(n850) );
  XOR2X1 U903 ( .A(\U_1/U_3/TX_CRC [15]), .B(\U_1/PROCESSED_DATA [7]), .Y(n834) );
  XNOR2X1 U904 ( .A(n12029), .B(n854), .Y(n856) );
  XOR2X1 U905 ( .A(n847), .B(n843), .Y(n854) );
  XNOR2X1 U906 ( .A(n842), .B(n846), .Y(n843) );
  XNOR2X1 U907 ( .A(n12041), .B(\U_1/PROCESSED_DATA [3]), .Y(n846) );
  XNOR2X1 U909 ( .A(\U_1/U_3/TX_CRC [12]), .B(n12026), .Y(n842) );
  XOR2X1 U911 ( .A(n849), .B(n845), .Y(n847) );
  XOR2X1 U912 ( .A(\U_1/U_3/TX_CRC [10]), .B(\U_1/PROCESSED_DATA [2]), .Y(n845) );
  XNOR2X1 U913 ( .A(\U_1/U_3/TX_CRC [9]), .B(\U_1/PROCESSED_DATA [1]), .Y(n849) );
  XNOR2X1 U915 ( .A(n838), .B(n841), .Y(n839) );
  XOR2X1 U916 ( .A(\U_1/U_3/TX_CRC [13]), .B(\U_1/PROCESSED_DATA [5]), .Y(n841) );
  XNOR2X1 U917 ( .A(\U_1/U_3/TX_CRC [14]), .B(n12032), .Y(n838) );
  NAND3X1 U920 ( .A(n862), .B(n11866), .C(n864), .Y(n819) );
  NOR2X1 U921 ( .A(n865), .B(n11846), .Y(n864) );
  AOI22X1 U924 ( .A(\U_1/PROCESSED_DATA [6]), .B(n9281), .C(n777), .D(
        \U_1/U_3/U_3/flop_data [6]), .Y(n867) );
  AOI22X1 U926 ( .A(\U_1/PROCESSED_DATA [5]), .B(n9281), .C(n777), .D(
        \U_1/U_3/U_3/flop_data [5]), .Y(n868) );
  AOI22X1 U928 ( .A(\U_1/PROCESSED_DATA [4]), .B(n9281), .C(n777), .D(
        \U_1/U_3/U_3/flop_data [4]), .Y(n869) );
  AOI22X1 U930 ( .A(\U_1/PROCESSED_DATA [3]), .B(n9281), .C(n777), .D(
        \U_1/U_3/U_3/flop_data [3]), .Y(n870) );
  AOI22X1 U932 ( .A(\U_1/PROCESSED_DATA [2]), .B(n9281), .C(n777), .D(
        \U_1/U_3/U_3/flop_data [2]), .Y(n871) );
  AOI22X1 U934 ( .A(\U_1/PROCESSED_DATA [1]), .B(n9281), .C(n777), .D(
        \U_1/U_3/U_3/flop_data [1]), .Y(n872) );
  AOI22X1 U936 ( .A(\U_1/PROCESSED_DATA [0]), .B(n9281), .C(n777), .D(
        \U_1/U_3/U_3/flop_data [0]), .Y(n873) );
  NAND3X1 U938 ( .A(n874), .B(n236), .C(n875), .Y(n777) );
  NOR2X1 U940 ( .A(RST), .B(n877), .Y(n874) );
  OAI21X1 U941 ( .A(n11644), .B(n879), .C(n880), .Y(n7792) );
  AOI22X1 U942 ( .A(\U_1/U_3/U_3/N90 ), .B(n881), .C(\U_1/U_3/U_3/N65 ), .D(
        n882), .Y(n880) );
  OAI21X1 U943 ( .A(n11867), .B(n879), .C(n884), .Y(n7793) );
  AOI22X1 U944 ( .A(\U_1/U_3/U_3/N89 ), .B(n881), .C(\U_1/U_3/U_3/N64 ), .D(
        n882), .Y(n884) );
  OAI21X1 U945 ( .A(n11872), .B(n879), .C(n886), .Y(n7794) );
  AOI22X1 U946 ( .A(\U_1/U_3/U_3/N88 ), .B(n881), .C(\U_1/U_3/U_3/N63 ), .D(
        n882), .Y(n886) );
  OAI21X1 U947 ( .A(n11871), .B(n879), .C(n888), .Y(n7795) );
  AOI22X1 U948 ( .A(\U_1/U_3/U_3/N87 ), .B(n881), .C(\U_1/U_3/U_3/N62 ), .D(
        n882), .Y(n888) );
  OAI21X1 U949 ( .A(n11870), .B(n879), .C(n890), .Y(n7796) );
  AOI22X1 U950 ( .A(\U_1/U_3/U_3/N86 ), .B(n881), .C(\U_1/U_3/U_3/N61 ), .D(
        n882), .Y(n890) );
  OAI21X1 U951 ( .A(n11869), .B(n879), .C(n892), .Y(n7797) );
  AOI22X1 U952 ( .A(\U_1/U_3/U_3/N85 ), .B(n881), .C(\U_1/U_3/U_3/N60 ), .D(
        n882), .Y(n892) );
  OAI21X1 U953 ( .A(n9276), .B(n11941), .C(n895), .Y(n7798) );
  NAND2X1 U954 ( .A(\U_1/U_0/U_0/N414 ), .B(n896), .Y(n895) );
  OAI21X1 U956 ( .A(n9276), .B(n11940), .C(n898), .Y(n7799) );
  NAND2X1 U957 ( .A(\U_1/U_0/U_0/N413 ), .B(n896), .Y(n898) );
  OAI21X1 U959 ( .A(n9276), .B(n11939), .C(n900), .Y(n7800) );
  NAND2X1 U960 ( .A(\U_1/U_0/U_0/N412 ), .B(n896), .Y(n900) );
  OAI21X1 U961 ( .A(n9276), .B(n11938), .C(n902), .Y(n7801) );
  NAND2X1 U962 ( .A(\U_1/U_0/U_0/N411 ), .B(n896), .Y(n902) );
  OAI21X1 U964 ( .A(n9276), .B(n11937), .C(n904), .Y(n7802) );
  NAND2X1 U965 ( .A(\U_1/U_0/U_0/N410 ), .B(n896), .Y(n904) );
  OAI21X1 U967 ( .A(n9276), .B(n11936), .C(n906), .Y(n7803) );
  NAND2X1 U968 ( .A(\U_1/U_0/U_0/N409 ), .B(n896), .Y(n906) );
  OAI21X1 U970 ( .A(n9276), .B(n11935), .C(n908), .Y(n7804) );
  NAND2X1 U971 ( .A(\U_1/U_0/U_0/N408 ), .B(n896), .Y(n908) );
  OAI21X1 U973 ( .A(n9276), .B(n11934), .C(n910), .Y(n7805) );
  NAND2X1 U974 ( .A(\U_1/U_0/U_0/N407 ), .B(n896), .Y(n910) );
  OAI21X1 U976 ( .A(n912), .B(n913), .C(n914), .Y(n7806) );
  OAI21X1 U977 ( .A(n9186), .B(n916), .C(\U_1/U_0/U_0/permuteComplete ), .Y(
        n914) );
  NAND2X1 U980 ( .A(n919), .B(n10518), .Y(n913) );
  NAND3X1 U982 ( .A(n921), .B(n322), .C(n10520), .Y(n917) );
  OAI22X1 U983 ( .A(n10343), .B(n12052), .C(n11923), .D(n926), .Y(n7807) );
  OAI22X1 U984 ( .A(n10343), .B(n11984), .C(n9554), .D(n926), .Y(n7808) );
  OAI22X1 U985 ( .A(n10343), .B(n11979), .C(n11975), .D(n926), .Y(n7809) );
  NAND3X1 U987 ( .A(n931), .B(n9534), .C(n11883), .Y(n926) );
  OAI21X1 U988 ( .A(n11883), .B(n11974), .C(n934), .Y(n7810) );
  NAND2X1 U989 ( .A(\U_1/U_0/U_0/N431 ), .B(n935), .Y(n934) );
  OAI21X1 U991 ( .A(n11883), .B(n11978), .C(n937), .Y(n7811) );
  NAND2X1 U992 ( .A(\U_1/U_0/U_0/N430 ), .B(n935), .Y(n937) );
  OAI21X1 U994 ( .A(n11883), .B(n11977), .C(n939), .Y(n7812) );
  NAND2X1 U995 ( .A(\U_1/U_0/U_0/N429 ), .B(n935), .Y(n939) );
  OAI21X1 U996 ( .A(n11883), .B(n11976), .C(n941), .Y(n7813) );
  NAND2X1 U997 ( .A(\U_1/U_0/U_0/N428 ), .B(n935), .Y(n941) );
  OAI21X1 U998 ( .A(n11883), .B(n9553), .C(n943), .Y(n7814) );
  NAND2X1 U999 ( .A(\U_1/U_0/U_0/N427 ), .B(n935), .Y(n943) );
  OAI21X1 U1001 ( .A(n11883), .B(n11975), .C(n944), .Y(n7815) );
  NAND2X1 U1002 ( .A(\U_1/U_0/U_0/N426 ), .B(n935), .Y(n944) );
  OAI21X1 U1004 ( .A(n11883), .B(n9554), .C(n945), .Y(n7816) );
  NAND2X1 U1005 ( .A(\U_1/U_0/U_0/N425 ), .B(n935), .Y(n945) );
  OAI21X1 U1006 ( .A(n11883), .B(n11923), .C(n946), .Y(n7817) );
  NAND2X1 U1007 ( .A(\U_1/U_0/U_0/N424 ), .B(n935), .Y(n946) );
  NOR2X1 U1008 ( .A(n912), .B(n919), .Y(n935) );
  NOR2X1 U1009 ( .A(n947), .B(n948), .Y(n919) );
  NAND3X1 U1010 ( .A(\U_1/U_0/U_0/si[7] ), .B(\U_1/U_0/U_0/si[6] ), .C(n949), 
        .Y(n948) );
  NOR2X1 U1011 ( .A(n11976), .B(n11977), .Y(n949) );
  NAND3X1 U1014 ( .A(\U_1/U_0/U_0/si[3] ), .B(\U_1/U_0/U_0/si[2] ), .C(n950), 
        .Y(n947) );
  NOR2X1 U1015 ( .A(n11923), .B(n9554), .Y(n950) );
  NAND3X1 U1019 ( .A(n11885), .B(n11889), .C(n954), .Y(n951) );
  NOR2X1 U1020 ( .A(n11899), .B(n956), .Y(n954) );
  OAI21X1 U1021 ( .A(n11884), .B(n11992), .C(n959), .Y(n7818) );
  NAND2X1 U1022 ( .A(\U_1/U_0/U_0/N480 ), .B(n11896), .Y(n959) );
  OAI21X1 U1024 ( .A(n11884), .B(n11991), .C(n962), .Y(n7819) );
  NAND2X1 U1025 ( .A(\U_1/U_0/U_0/N481 ), .B(n11896), .Y(n962) );
  OAI21X1 U1027 ( .A(n11884), .B(n11990), .C(n964), .Y(n7820) );
  NAND2X1 U1028 ( .A(\U_1/U_0/U_0/N482 ), .B(n11896), .Y(n964) );
  OAI21X1 U1030 ( .A(n11884), .B(n11989), .C(n966), .Y(n7821) );
  NAND2X1 U1031 ( .A(\U_1/U_0/U_0/N483 ), .B(n11896), .Y(n966) );
  OAI21X1 U1033 ( .A(n11884), .B(n11988), .C(n968), .Y(n7822) );
  NAND2X1 U1034 ( .A(\U_1/U_0/U_0/N484 ), .B(n11896), .Y(n968) );
  OAI21X1 U1036 ( .A(n11884), .B(n11987), .C(n970), .Y(n7823) );
  NAND2X1 U1037 ( .A(\U_1/U_0/U_0/N485 ), .B(n11896), .Y(n970) );
  OAI21X1 U1039 ( .A(n11884), .B(n11986), .C(n972), .Y(n7824) );
  NAND2X1 U1040 ( .A(\U_1/U_0/U_0/N486 ), .B(n11896), .Y(n972) );
  OAI21X1 U1042 ( .A(n11884), .B(n11985), .C(n974), .Y(n7825) );
  NAND2X1 U1043 ( .A(\U_1/U_0/U_0/N487 ), .B(n11896), .Y(n974) );
  NAND3X1 U1046 ( .A(n11885), .B(n11891), .C(n977), .Y(n975) );
  NOR2X1 U1047 ( .A(n11900), .B(n979), .Y(n977) );
  NAND2X1 U1048 ( .A(n912), .B(n980), .Y(n979) );
  OAI21X1 U1050 ( .A(n9280), .B(n12033), .C(n984), .Y(n7826) );
  AOI22X1 U1051 ( .A(DATA_IN_S[7]), .B(n10519), .C(\U_1/U_0/U_0/N527 ), .D(
        n986), .Y(n984) );
  OAI21X1 U1052 ( .A(n9280), .B(n12030), .C(n988), .Y(n7827) );
  AOI22X1 U1053 ( .A(DATA_IN_S[6]), .B(n10519), .C(\U_1/U_0/U_0/N526 ), .D(
        n986), .Y(n988) );
  OAI21X1 U1054 ( .A(n9280), .B(n12027), .C(n990), .Y(n7828) );
  AOI22X1 U1055 ( .A(DATA_IN_S[5]), .B(n10519), .C(\U_1/U_0/U_0/N525 ), .D(
        n986), .Y(n990) );
  OAI21X1 U1056 ( .A(n9280), .B(n12024), .C(n992), .Y(n7829) );
  AOI22X1 U1057 ( .A(DATA_IN_S[4]), .B(n10519), .C(\U_1/U_0/U_0/N524 ), .D(
        n986), .Y(n992) );
  OAI21X1 U1058 ( .A(n9280), .B(n12022), .C(n994), .Y(n7830) );
  AOI22X1 U1059 ( .A(DATA_IN_S[3]), .B(n10519), .C(\U_1/U_0/U_0/N523 ), .D(
        n986), .Y(n994) );
  OAI21X1 U1060 ( .A(n9280), .B(n12020), .C(n996), .Y(n7831) );
  AOI22X1 U1061 ( .A(DATA_IN_S[2]), .B(n10519), .C(\U_1/U_0/U_0/N522 ), .D(
        n986), .Y(n996) );
  OAI21X1 U1062 ( .A(n9280), .B(n12018), .C(n998), .Y(n7832) );
  AOI22X1 U1063 ( .A(DATA_IN_S[1]), .B(n10519), .C(\U_1/U_0/U_0/N521 ), .D(
        n986), .Y(n998) );
  OAI21X1 U1064 ( .A(n9280), .B(n12016), .C(n1000), .Y(n7833) );
  AOI22X1 U1065 ( .A(DATA_IN_S[0]), .B(n10519), .C(\U_1/U_0/U_0/N520 ), .D(
        n986), .Y(n1000) );
  NOR2X1 U1066 ( .A(n1001), .B(n9167), .Y(n986) );
  OAI21X1 U1069 ( .A(n11896), .B(n1004), .C(n9280), .Y(n1003) );
  NAND3X1 U1071 ( .A(n1007), .B(n1008), .C(n1009), .Y(n1006) );
  NAND3X1 U1074 ( .A(n1011), .B(n9198), .C(n1013), .Y(n1010) );
  NOR2X1 U1075 ( .A(n11914), .B(n981), .Y(n1013) );
  NAND3X1 U1076 ( .A(n11892), .B(n1016), .C(n1017), .Y(n981) );
  NOR2X1 U1077 ( .A(RST), .B(n9197), .Y(n1011) );
  NAND3X1 U1078 ( .A(n1018), .B(n322), .C(n1019), .Y(n1005) );
  AOI22X1 U1081 ( .A(n1022), .B(\U_1/U_0/U_0/extratemp[0] ), .C(DATA_IN_S[0]), 
        .D(n10529), .Y(n1021) );
  AOI22X1 U1083 ( .A(n1022), .B(\U_1/U_0/U_0/extratemp[1] ), .C(DATA_IN_S[1]), 
        .D(n10529), .Y(n1024) );
  AOI22X1 U1085 ( .A(n1022), .B(\U_1/U_0/U_0/extratemp[2] ), .C(DATA_IN_S[2]), 
        .D(n10529), .Y(n1025) );
  AOI22X1 U1087 ( .A(n1022), .B(\U_1/U_0/U_0/extratemp[3] ), .C(DATA_IN_S[3]), 
        .D(n10529), .Y(n1026) );
  AOI22X1 U1089 ( .A(n1022), .B(\U_1/U_0/U_0/extratemp[4] ), .C(DATA_IN_S[4]), 
        .D(n10529), .Y(n1027) );
  AOI22X1 U1091 ( .A(n1022), .B(\U_1/U_0/U_0/extratemp[5] ), .C(DATA_IN_S[5]), 
        .D(n10529), .Y(n1028) );
  AOI22X1 U1093 ( .A(n1022), .B(\U_1/U_0/U_0/extratemp[6] ), .C(DATA_IN_S[6]), 
        .D(n10529), .Y(n1029) );
  AOI22X1 U1095 ( .A(n1022), .B(\U_1/U_0/U_0/extratemp[7] ), .C(DATA_IN_S[7]), 
        .D(n10529), .Y(n1030) );
  NAND3X1 U1097 ( .A(n1017), .B(n931), .C(n10530), .Y(n1022) );
  OAI22X1 U1100 ( .A(n9279), .B(n11994), .C(n1036), .D(n11993), .Y(n7842) );
  OAI22X1 U1103 ( .A(n9279), .B(n12007), .C(n1036), .D(n11995), .Y(n7843) );
  OAI22X1 U1106 ( .A(n9279), .B(n12006), .C(n1036), .D(n11996), .Y(n7844) );
  OAI22X1 U1109 ( .A(n9279), .B(n12005), .C(n1036), .D(n11997), .Y(n7845) );
  OAI22X1 U1112 ( .A(n9279), .B(n12004), .C(n1036), .D(n11998), .Y(n7846) );
  OAI22X1 U1115 ( .A(n9279), .B(n12003), .C(n1036), .D(n11999), .Y(n7847) );
  OAI22X1 U1118 ( .A(n9279), .B(n12002), .C(n1036), .D(n12000), .Y(n7848) );
  OAI22X1 U1121 ( .A(n9279), .B(n12001), .C(n1036), .D(\U_1/U_0/U_0/inti[0] ), 
        .Y(n7849) );
  NAND2X1 U1123 ( .A(n11899), .B(n9279), .Y(n1036) );
  NOR2X1 U1125 ( .A(n1032), .B(n956), .Y(n1034) );
  NAND3X1 U1126 ( .A(n11885), .B(n11889), .C(n1052), .Y(n1032) );
  NOR2X1 U1127 ( .A(RST), .B(n11915), .Y(n1052) );
  AOI22X1 U1130 ( .A(n1056), .B(\U_1/U_0/U_0/delaydata [6]), .C(
        \U_1/PRGA_IN [6]), .D(n9278), .Y(n1055) );
  AOI22X1 U1132 ( .A(n1056), .B(\U_1/U_0/U_0/delaydata [5]), .C(
        \U_1/PRGA_IN [5]), .D(n9278), .Y(n1058) );
  AOI22X1 U1134 ( .A(n1056), .B(\U_1/U_0/U_0/delaydata [4]), .C(
        \U_1/PRGA_IN [4]), .D(n9278), .Y(n1059) );
  AOI22X1 U1136 ( .A(n1056), .B(\U_1/U_0/U_0/delaydata [3]), .C(
        \U_1/PRGA_IN [3]), .D(n9278), .Y(n1060) );
  AOI22X1 U1138 ( .A(n1056), .B(\U_1/U_0/U_0/delaydata [2]), .C(
        \U_1/PRGA_IN [2]), .D(n9278), .Y(n1061) );
  AOI22X1 U1140 ( .A(n1056), .B(\U_1/U_0/U_0/delaydata [1]), .C(
        \U_1/PRGA_IN [1]), .D(n9278), .Y(n1062) );
  AOI22X1 U1142 ( .A(n1056), .B(\U_1/U_0/U_0/delaydata [0]), .C(
        \U_1/PRGA_IN [0]), .D(n9278), .Y(n1063) );
  AOI22X1 U1144 ( .A(n1056), .B(\U_1/U_0/U_0/delaydata [7]), .C(
        \U_1/PRGA_IN [7]), .D(n9278), .Y(n1064) );
  NAND2X1 U1146 ( .A(n9277), .B(n931), .Y(n1056) );
  OAI21X1 U1147 ( .A(n9277), .B(n12015), .C(n1067), .Y(n7858) );
  NAND2X1 U1148 ( .A(\U_1/U_0/U_0/N519 ), .B(n1068), .Y(n1067) );
  OAI21X1 U1150 ( .A(n9277), .B(n12014), .C(n1070), .Y(n7859) );
  NAND2X1 U1151 ( .A(\U_1/U_0/U_0/N518 ), .B(n1068), .Y(n1070) );
  OAI21X1 U1153 ( .A(n9277), .B(n12013), .C(n1072), .Y(n7860) );
  NAND2X1 U1154 ( .A(\U_1/U_0/U_0/N517 ), .B(n1068), .Y(n1072) );
  OAI21X1 U1156 ( .A(n9277), .B(n12012), .C(n1074), .Y(n7861) );
  NAND2X1 U1157 ( .A(\U_1/U_0/U_0/N516 ), .B(n1068), .Y(n1074) );
  OAI21X1 U1159 ( .A(n9277), .B(n12011), .C(n1076), .Y(n7862) );
  NAND2X1 U1160 ( .A(\U_1/U_0/U_0/N515 ), .B(n1068), .Y(n1076) );
  OAI21X1 U1162 ( .A(n9277), .B(n12010), .C(n1078), .Y(n7863) );
  NAND2X1 U1163 ( .A(\U_1/U_0/U_0/N514 ), .B(n1068), .Y(n1078) );
  OAI21X1 U1165 ( .A(n9277), .B(n12009), .C(n1080), .Y(n7864) );
  NAND2X1 U1166 ( .A(\U_1/U_0/U_0/N513 ), .B(n1068), .Y(n1080) );
  OAI21X1 U1168 ( .A(n9277), .B(n12008), .C(n1082), .Y(n7865) );
  NAND2X1 U1169 ( .A(\U_1/U_0/U_0/N512 ), .B(n1068), .Y(n1082) );
  NOR2X1 U1172 ( .A(n1084), .B(n1085), .Y(n1065) );
  NAND3X1 U1173 ( .A(n11885), .B(n9200), .C(n1087), .Y(n1085) );
  NOR2X1 U1174 ( .A(n9199), .B(n11900), .Y(n1087) );
  NAND3X1 U1177 ( .A(n1091), .B(n1092), .C(n1093), .Y(n1090) );
  NOR2X1 U1178 ( .A(n1094), .B(n1095), .Y(n1093) );
  NAND2X1 U1179 ( .A(n1018), .B(n1096), .Y(n1095) );
  NAND3X1 U1180 ( .A(n322), .B(n1097), .C(n1001), .Y(n1094) );
  NOR2X1 U1182 ( .A(n11922), .B(n11914), .Y(n1091) );
  NAND3X1 U1183 ( .A(n912), .B(n321), .C(n1101), .Y(n1084) );
  NOR2X1 U1184 ( .A(RST), .B(n11896), .Y(n1101) );
  AOI22X1 U1186 ( .A(\U_1/U_0/PLAINKEY [6]), .B(n9468), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[0][6] ), .Y(n1102) );
  AOI22X1 U1188 ( .A(\U_1/U_0/PLAINKEY [5]), .B(n9461), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[0][5] ), .Y(n1105) );
  AOI22X1 U1190 ( .A(\U_1/U_0/PLAINKEY [4]), .B(n9461), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[0][4] ), .Y(n1106) );
  OAI22X1 U1191 ( .A(n11541), .B(n9459), .C(n9473), .D(n11945), .Y(n7869) );
  OAI22X1 U1193 ( .A(n11539), .B(n9460), .C(n9473), .D(n11946), .Y(n7870) );
  OAI22X1 U1195 ( .A(n11537), .B(n9460), .C(n9473), .D(n11947), .Y(n7871) );
  OAI22X1 U1197 ( .A(n11535), .B(n9459), .C(n9473), .D(n11948), .Y(n7872) );
  AOI22X1 U1200 ( .A(\U_1/U_0/PLAINKEY [15]), .B(n9462), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[1][7] ), .Y(n1111) );
  AOI22X1 U1202 ( .A(\U_1/U_0/PLAINKEY [7]), .B(n9462), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[0][7] ), .Y(n1112) );
  AOI22X1 U1204 ( .A(\U_1/U_0/PLAINKEY [56]), .B(n9462), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[7][0] ), .Y(n1113) );
  AOI22X1 U1206 ( .A(\U_1/U_0/PLAINKEY [57]), .B(n9463), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[7][1] ), .Y(n1114) );
  AOI22X1 U1208 ( .A(\U_1/U_0/PLAINKEY [58]), .B(n9463), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[7][2] ), .Y(n1115) );
  AOI22X1 U1210 ( .A(\U_1/U_0/PLAINKEY [59]), .B(n9463), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[7][3] ), .Y(n1116) );
  AOI22X1 U1212 ( .A(\U_1/U_0/PLAINKEY [60]), .B(n9464), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[7][4] ), .Y(n1117) );
  AOI22X1 U1214 ( .A(\U_1/U_0/PLAINKEY [61]), .B(n9464), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[7][5] ), .Y(n1118) );
  AOI22X1 U1216 ( .A(\U_1/U_0/PLAINKEY [62]), .B(n9464), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[7][6] ), .Y(n1119) );
  AOI22X1 U1218 ( .A(\U_1/U_0/PLAINKEY [63]), .B(n9465), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[7][7] ), .Y(n1120) );
  AOI22X1 U1220 ( .A(\U_1/U_0/PLAINKEY [48]), .B(n9465), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[6][0] ), .Y(n1121) );
  AOI22X1 U1222 ( .A(\U_1/U_0/PLAINKEY [49]), .B(n9465), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[6][1] ), .Y(n1122) );
  AOI22X1 U1224 ( .A(\U_1/U_0/PLAINKEY [50]), .B(n9466), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[6][2] ), .Y(n1123) );
  AOI22X1 U1226 ( .A(\U_1/U_0/PLAINKEY [51]), .B(n9466), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[6][3] ), .Y(n1124) );
  AOI22X1 U1228 ( .A(\U_1/U_0/PLAINKEY [52]), .B(n9466), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[6][4] ), .Y(n1125) );
  AOI22X1 U1230 ( .A(\U_1/U_0/PLAINKEY [53]), .B(n9467), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[6][5] ), .Y(n1126) );
  AOI22X1 U1232 ( .A(\U_1/U_0/PLAINKEY [54]), .B(n9467), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[6][6] ), .Y(n1127) );
  AOI22X1 U1234 ( .A(\U_1/U_0/PLAINKEY [55]), .B(n9467), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[6][7] ), .Y(n1128) );
  AOI22X1 U1236 ( .A(\U_1/U_0/PLAINKEY [40]), .B(n9467), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[5][0] ), .Y(n1129) );
  AOI22X1 U1238 ( .A(\U_1/U_0/PLAINKEY [41]), .B(n9467), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[5][1] ), .Y(n1130) );
  AOI22X1 U1240 ( .A(\U_1/U_0/PLAINKEY [42]), .B(n9467), .C(n9457), .D(
        \U_1/U_0/U_0/keyTable[5][2] ), .Y(n1131) );
  AOI22X1 U1242 ( .A(\U_1/U_0/PLAINKEY [43]), .B(n9467), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[5][3] ), .Y(n1132) );
  AOI22X1 U1244 ( .A(\U_1/U_0/PLAINKEY [44]), .B(n9468), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[5][4] ), .Y(n1133) );
  AOI22X1 U1246 ( .A(\U_1/U_0/PLAINKEY [45]), .B(n9468), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[5][5] ), .Y(n1134) );
  AOI22X1 U1248 ( .A(\U_1/U_0/PLAINKEY [46]), .B(n9468), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[5][6] ), .Y(n1135) );
  AOI22X1 U1250 ( .A(\U_1/U_0/PLAINKEY [47]), .B(n9468), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[5][7] ), .Y(n1136) );
  AOI22X1 U1252 ( .A(\U_1/U_0/PLAINKEY [32]), .B(n9468), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[4][0] ), .Y(n1137) );
  AOI22X1 U1254 ( .A(\U_1/U_0/PLAINKEY [33]), .B(n9468), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[4][1] ), .Y(n1138) );
  AOI22X1 U1256 ( .A(\U_1/U_0/PLAINKEY [34]), .B(n9469), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[4][2] ), .Y(n1139) );
  AOI22X1 U1258 ( .A(\U_1/U_0/PLAINKEY [35]), .B(n9469), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[4][3] ), .Y(n1140) );
  AOI22X1 U1260 ( .A(\U_1/U_0/PLAINKEY [36]), .B(n9469), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[4][4] ), .Y(n1141) );
  AOI22X1 U1262 ( .A(\U_1/U_0/PLAINKEY [37]), .B(n9469), .C(n9458), .D(
        \U_1/U_0/U_0/keyTable[4][5] ), .Y(n1142) );
  AOI22X1 U1264 ( .A(\U_1/U_0/PLAINKEY [38]), .B(n9469), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[4][6] ), .Y(n1143) );
  AOI22X1 U1266 ( .A(\U_1/U_0/PLAINKEY [39]), .B(n9469), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[4][7] ), .Y(n1144) );
  AOI22X1 U1268 ( .A(\U_1/U_0/PLAINKEY [24]), .B(n9469), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[3][0] ), .Y(n1145) );
  AOI22X1 U1270 ( .A(\U_1/U_0/PLAINKEY [25]), .B(n9470), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[3][1] ), .Y(n1146) );
  AOI22X1 U1272 ( .A(\U_1/U_0/PLAINKEY [26]), .B(n9470), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[3][2] ), .Y(n1147) );
  AOI22X1 U1274 ( .A(\U_1/U_0/PLAINKEY [27]), .B(n9470), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[3][3] ), .Y(n1148) );
  AOI22X1 U1276 ( .A(\U_1/U_0/PLAINKEY [28]), .B(n9470), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[3][4] ), .Y(n1149) );
  AOI22X1 U1278 ( .A(\U_1/U_0/PLAINKEY [29]), .B(n9470), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[3][5] ), .Y(n1150) );
  AOI22X1 U1280 ( .A(\U_1/U_0/PLAINKEY [30]), .B(n9470), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[3][6] ), .Y(n1151) );
  AOI22X1 U1282 ( .A(\U_1/U_0/PLAINKEY [31]), .B(n9470), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[3][7] ), .Y(n1152) );
  AOI22X1 U1284 ( .A(\U_1/U_0/PLAINKEY [16]), .B(n9471), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[2][0] ), .Y(n1153) );
  AOI22X1 U1286 ( .A(\U_1/U_0/PLAINKEY [17]), .B(n9471), .C(n9459), .D(
        \U_1/U_0/U_0/keyTable[2][1] ), .Y(n1154) );
  AOI22X1 U1288 ( .A(\U_1/U_0/PLAINKEY [18]), .B(n9471), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[2][2] ), .Y(n1155) );
  AOI22X1 U1290 ( .A(\U_1/U_0/PLAINKEY [19]), .B(n9471), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[2][3] ), .Y(n1156) );
  AOI22X1 U1292 ( .A(\U_1/U_0/PLAINKEY [20]), .B(n9471), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[2][4] ), .Y(n1157) );
  AOI22X1 U1294 ( .A(\U_1/U_0/PLAINKEY [21]), .B(n9471), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[2][5] ), .Y(n1158) );
  AOI22X1 U1296 ( .A(\U_1/U_0/PLAINKEY [22]), .B(n9471), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[2][6] ), .Y(n1159) );
  AOI22X1 U1298 ( .A(\U_1/U_0/PLAINKEY [23]), .B(n9472), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[2][7] ), .Y(n1160) );
  AOI22X1 U1300 ( .A(\U_1/U_0/PLAINKEY [8]), .B(n9472), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[1][0] ), .Y(n1161) );
  AOI22X1 U1302 ( .A(\U_1/U_0/PLAINKEY [9]), .B(n9472), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[1][1] ), .Y(n1162) );
  AOI22X1 U1304 ( .A(\U_1/U_0/PLAINKEY [10]), .B(n9472), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[1][2] ), .Y(n1163) );
  AOI22X1 U1306 ( .A(\U_1/U_0/PLAINKEY [11]), .B(n9472), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[1][3] ), .Y(n1164) );
  AOI22X1 U1308 ( .A(\U_1/U_0/PLAINKEY [12]), .B(n9472), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[1][4] ), .Y(n1165) );
  AOI22X1 U1310 ( .A(\U_1/U_0/PLAINKEY [13]), .B(n9472), .C(n9460), .D(
        \U_1/U_0/U_0/keyTable[1][5] ), .Y(n1166) );
  AOI22X1 U1312 ( .A(\U_1/U_0/PLAINKEY [14]), .B(n9461), .C(n9456), .D(
        \U_1/U_0/U_0/keyTable[1][6] ), .Y(n1167) );
  NOR2X1 U1315 ( .A(n1168), .B(n1169), .Y(n893) );
  NAND3X1 U1316 ( .A(n318), .B(n11881), .C(n11898), .Y(n1169) );
  NAND3X1 U1317 ( .A(n11921), .B(n9516), .C(n11892), .Y(n1168) );
  OAI21X1 U1318 ( .A(n10282), .B(n11840), .C(n1173), .Y(n7930) );
  OAI21X1 U1319 ( .A(n1174), .B(n1175), .C(n10282), .Y(n1173) );
  NAND3X1 U1321 ( .A(n1178), .B(n1179), .C(n1180), .Y(n1177) );
  NOR2X1 U1322 ( .A(n1181), .B(n1182), .Y(n1180) );
  OAI22X1 U1323 ( .A(n1183), .B(n11771), .C(n1185), .D(n11781), .Y(n1182) );
  OAI22X1 U1324 ( .A(n1187), .B(n11751), .C(n1189), .D(n11761), .Y(n1181) );
  AOI22X1 U1325 ( .A(\U_1/U_1/U_1/opcode[26][1] ), .B(n1191), .C(
        \U_1/U_1/U_1/opcode[27][1] ), .D(n1192), .Y(n1179) );
  AOI22X1 U1326 ( .A(\U_1/U_1/U_1/opcode[24][1] ), .B(n1193), .C(
        \U_1/U_1/U_1/opcode[25][1] ), .D(n1194), .Y(n1178) );
  NAND3X1 U1327 ( .A(n1195), .B(n1196), .C(n1197), .Y(n1176) );
  NOR2X1 U1328 ( .A(n1198), .B(n1199), .Y(n1197) );
  OAI22X1 U1329 ( .A(n1200), .B(n11811), .C(n1202), .D(n11821), .Y(n1199) );
  OAI22X1 U1330 ( .A(n1204), .B(n11791), .C(n1206), .D(n11801), .Y(n1198) );
  AOI22X1 U1331 ( .A(\U_1/U_1/U_1/opcode[22][1] ), .B(n1208), .C(
        \U_1/U_1/U_1/opcode[23][1] ), .D(n1209), .Y(n1196) );
  AOI22X1 U1332 ( .A(\U_1/U_1/U_1/opcode[20][1] ), .B(n1210), .C(
        \U_1/U_1/U_1/opcode[21][1] ), .D(n1211), .Y(n1195) );
  NAND3X1 U1334 ( .A(n1214), .B(n1215), .C(n1216), .Y(n1213) );
  NOR2X1 U1335 ( .A(n1217), .B(n1218), .Y(n1216) );
  OAI22X1 U1336 ( .A(n1219), .B(n11741), .C(n1221), .D(n11706), .Y(n1218) );
  OAI22X1 U1337 ( .A(n1223), .B(n11721), .C(n1225), .D(n11731), .Y(n1217) );
  AOI22X1 U1338 ( .A(\U_1/U_1/U_1/opcode[14][1] ), .B(n1227), .C(
        \U_1/U_1/U_1/opcode[15][1] ), .D(n1228), .Y(n1215) );
  AOI22X1 U1339 ( .A(\U_1/U_1/U_1/opcode[12][1] ), .B(n1229), .C(
        \U_1/U_1/U_1/opcode[13][1] ), .D(n1230), .Y(n1214) );
  NAND3X1 U1340 ( .A(n1231), .B(n1232), .C(n1233), .Y(n1212) );
  NOR2X1 U1341 ( .A(n1234), .B(n1235), .Y(n1233) );
  OAI22X1 U1342 ( .A(n1236), .B(n11681), .C(n1238), .D(n11671), .Y(n1235) );
  OAI22X1 U1343 ( .A(n1240), .B(n11711), .C(n1242), .D(n11709), .Y(n1234) );
  AOI22X1 U1344 ( .A(\U_1/U_1/U_1/opcode[1][1] ), .B(n1244), .C(
        \U_1/U_1/U_1/opcode[0][1] ), .D(n1245), .Y(n1232) );
  AOI22X1 U1345 ( .A(\U_1/U_1/U_1/opcode[3][1] ), .B(n1246), .C(
        \U_1/U_1/U_1/opcode[2][1] ), .D(n1247), .Y(n1231) );
  OAI21X1 U1347 ( .A(n10282), .B(n11839), .C(n1248), .Y(n7931) );
  OAI21X1 U1348 ( .A(n1249), .B(n1250), .C(n10282), .Y(n1248) );
  NAND3X1 U1350 ( .A(n1253), .B(n1254), .C(n1255), .Y(n1252) );
  NOR2X1 U1351 ( .A(n1256), .B(n1257), .Y(n1255) );
  OAI22X1 U1352 ( .A(n1183), .B(n11770), .C(n1185), .D(n11780), .Y(n1257) );
  OAI22X1 U1353 ( .A(n1187), .B(n11750), .C(n1189), .D(n11760), .Y(n1256) );
  AOI22X1 U1354 ( .A(\U_1/U_1/U_1/opcode[26][0] ), .B(n1191), .C(
        \U_1/U_1/U_1/opcode[27][0] ), .D(n1192), .Y(n1254) );
  AOI22X1 U1355 ( .A(\U_1/U_1/U_1/opcode[24][0] ), .B(n1193), .C(
        \U_1/U_1/U_1/opcode[25][0] ), .D(n1194), .Y(n1253) );
  NAND3X1 U1356 ( .A(n1262), .B(n1263), .C(n1264), .Y(n1251) );
  NOR2X1 U1357 ( .A(n1265), .B(n1266), .Y(n1264) );
  OAI22X1 U1358 ( .A(n1200), .B(n11810), .C(n1202), .D(n11820), .Y(n1266) );
  OAI22X1 U1359 ( .A(n1204), .B(n11790), .C(n1206), .D(n11800), .Y(n1265) );
  AOI22X1 U1360 ( .A(\U_1/U_1/U_1/opcode[22][0] ), .B(n1208), .C(
        \U_1/U_1/U_1/opcode[23][0] ), .D(n1209), .Y(n1263) );
  AOI22X1 U1361 ( .A(\U_1/U_1/U_1/opcode[20][0] ), .B(n1210), .C(
        \U_1/U_1/U_1/opcode[21][0] ), .D(n1211), .Y(n1262) );
  NAND3X1 U1363 ( .A(n1273), .B(n1274), .C(n1275), .Y(n1272) );
  NOR2X1 U1364 ( .A(n1276), .B(n1277), .Y(n1275) );
  OAI22X1 U1365 ( .A(n1219), .B(n11740), .C(n1221), .D(n11707), .Y(n1277) );
  OAI22X1 U1366 ( .A(n1223), .B(n11720), .C(n1225), .D(n11730), .Y(n1276) );
  AOI22X1 U1367 ( .A(\U_1/U_1/U_1/opcode[14][0] ), .B(n1227), .C(
        \U_1/U_1/U_1/opcode[15][0] ), .D(n1228), .Y(n1274) );
  AOI22X1 U1368 ( .A(\U_1/U_1/U_1/opcode[12][0] ), .B(n1229), .C(
        \U_1/U_1/U_1/opcode[13][0] ), .D(n1230), .Y(n1273) );
  NAND3X1 U1369 ( .A(n1282), .B(n1283), .C(n1284), .Y(n1271) );
  NOR2X1 U1370 ( .A(n1285), .B(n1286), .Y(n1284) );
  OAI22X1 U1371 ( .A(n1236), .B(n11680), .C(n1238), .D(n11670), .Y(n1286) );
  OAI22X1 U1372 ( .A(n1240), .B(n11710), .C(n1242), .D(n11708), .Y(n1285) );
  AOI22X1 U1373 ( .A(\U_1/U_1/U_1/opcode[1][0] ), .B(n1244), .C(
        \U_1/U_1/U_1/opcode[0][0] ), .D(n1245), .Y(n1283) );
  AOI22X1 U1374 ( .A(\U_1/U_1/U_1/opcode[3][0] ), .B(n1246), .C(
        \U_1/U_1/U_1/opcode[2][0] ), .D(n1247), .Y(n1282) );
  OAI21X1 U1376 ( .A(n10282), .B(n11838), .C(n1291), .Y(n7932) );
  OAI21X1 U1377 ( .A(n1292), .B(n1293), .C(n10282), .Y(n1291) );
  NAND3X1 U1379 ( .A(n1296), .B(n1297), .C(n1298), .Y(n1295) );
  NOR2X1 U1380 ( .A(n1299), .B(n1300), .Y(n1298) );
  OAI22X1 U1381 ( .A(n1183), .B(n11779), .C(n1185), .D(n11789), .Y(n1300) );
  OAI22X1 U1382 ( .A(n1187), .B(n11759), .C(n1189), .D(n11769), .Y(n1299) );
  AOI22X1 U1383 ( .A(\U_1/U_1/U_1/memory[26][7] ), .B(n1191), .C(
        \U_1/U_1/U_1/memory[27][7] ), .D(n1192), .Y(n1297) );
  AOI22X1 U1384 ( .A(\U_1/U_1/U_1/memory[24][7] ), .B(n1193), .C(
        \U_1/U_1/U_1/memory[25][7] ), .D(n1194), .Y(n1296) );
  NAND3X1 U1385 ( .A(n1305), .B(n1306), .C(n1307), .Y(n1294) );
  NOR2X1 U1386 ( .A(n1308), .B(n1309), .Y(n1307) );
  OAI22X1 U1387 ( .A(n1200), .B(n11819), .C(n1202), .D(n11826), .Y(n1309) );
  OAI22X1 U1388 ( .A(n1204), .B(n11799), .C(n1206), .D(n11809), .Y(n1308) );
  AOI22X1 U1389 ( .A(\U_1/U_1/U_1/memory[22][7] ), .B(n1208), .C(
        \U_1/U_1/U_1/memory[23][7] ), .D(n1209), .Y(n1306) );
  AOI22X1 U1390 ( .A(\U_1/U_1/U_1/memory[20][7] ), .B(n1210), .C(
        \U_1/U_1/U_1/memory[21][7] ), .D(n1211), .Y(n1305) );
  NAND3X1 U1392 ( .A(n1316), .B(n1317), .C(n1318), .Y(n1315) );
  NOR2X1 U1393 ( .A(n1319), .B(n1320), .Y(n1318) );
  OAI22X1 U1394 ( .A(n1219), .B(n11749), .C(n1221), .D(n11719), .Y(n1320) );
  OAI22X1 U1395 ( .A(n1223), .B(n11729), .C(n1225), .D(n11739), .Y(n1319) );
  AOI22X1 U1396 ( .A(\U_1/U_1/U_1/memory[14][7] ), .B(n1227), .C(
        \U_1/U_1/U_1/memory[15][7] ), .D(n1228), .Y(n1317) );
  AOI22X1 U1397 ( .A(\U_1/U_1/U_1/memory[12][7] ), .B(n1229), .C(
        \U_1/U_1/U_1/memory[13][7] ), .D(n1230), .Y(n1316) );
  NAND3X1 U1398 ( .A(n1325), .B(n1326), .C(n1327), .Y(n1314) );
  NOR2X1 U1399 ( .A(n1328), .B(n1329), .Y(n1327) );
  OAI22X1 U1400 ( .A(n1236), .B(n11689), .C(n1238), .D(n11679), .Y(n1329) );
  OAI22X1 U1401 ( .A(n1240), .B(n11699), .C(n1242), .D(n11697), .Y(n1328) );
  AOI22X1 U1402 ( .A(\U_1/U_1/U_1/memory[1][7] ), .B(n1244), .C(
        \U_1/U_1/U_1/memory[0][7] ), .D(n1245), .Y(n1326) );
  AOI22X1 U1403 ( .A(\U_1/U_1/U_1/memory[3][7] ), .B(n1246), .C(
        \U_1/U_1/U_1/memory[2][7] ), .D(n1247), .Y(n1325) );
  OAI21X1 U1405 ( .A(n10282), .B(n11837), .C(n1334), .Y(n7933) );
  OAI21X1 U1406 ( .A(n1335), .B(n1336), .C(n10282), .Y(n1334) );
  NAND3X1 U1408 ( .A(n1339), .B(n1340), .C(n1341), .Y(n1338) );
  NOR2X1 U1409 ( .A(n1342), .B(n1343), .Y(n1341) );
  OAI22X1 U1410 ( .A(n1183), .B(n11778), .C(n1185), .D(n11788), .Y(n1343) );
  OAI22X1 U1411 ( .A(n1187), .B(n11758), .C(n1189), .D(n11768), .Y(n1342) );
  AOI22X1 U1412 ( .A(\U_1/U_1/U_1/memory[26][6] ), .B(n1191), .C(
        \U_1/U_1/U_1/memory[27][6] ), .D(n1192), .Y(n1340) );
  AOI22X1 U1413 ( .A(\U_1/U_1/U_1/memory[24][6] ), .B(n1193), .C(
        \U_1/U_1/U_1/memory[25][6] ), .D(n1194), .Y(n1339) );
  NAND3X1 U1414 ( .A(n1348), .B(n1349), .C(n1350), .Y(n1337) );
  NOR2X1 U1415 ( .A(n1351), .B(n1352), .Y(n1350) );
  OAI22X1 U1416 ( .A(n1200), .B(n11818), .C(n1202), .D(n11825), .Y(n1352) );
  OAI22X1 U1417 ( .A(n1204), .B(n11798), .C(n1206), .D(n11808), .Y(n1351) );
  AOI22X1 U1418 ( .A(\U_1/U_1/U_1/memory[22][6] ), .B(n1208), .C(
        \U_1/U_1/U_1/memory[23][6] ), .D(n1209), .Y(n1349) );
  AOI22X1 U1419 ( .A(\U_1/U_1/U_1/memory[20][6] ), .B(n1210), .C(
        \U_1/U_1/U_1/memory[21][6] ), .D(n1211), .Y(n1348) );
  NAND3X1 U1421 ( .A(n1359), .B(n1360), .C(n1361), .Y(n1358) );
  NOR2X1 U1422 ( .A(n1362), .B(n1363), .Y(n1361) );
  OAI22X1 U1423 ( .A(n1219), .B(n11748), .C(n1221), .D(n11718), .Y(n1363) );
  OAI22X1 U1424 ( .A(n1223), .B(n11728), .C(n1225), .D(n11738), .Y(n1362) );
  AOI22X1 U1425 ( .A(\U_1/U_1/U_1/memory[14][6] ), .B(n1227), .C(
        \U_1/U_1/U_1/memory[15][6] ), .D(n1228), .Y(n1360) );
  AOI22X1 U1426 ( .A(\U_1/U_1/U_1/memory[12][6] ), .B(n1229), .C(
        \U_1/U_1/U_1/memory[13][6] ), .D(n1230), .Y(n1359) );
  NAND3X1 U1427 ( .A(n1368), .B(n1369), .C(n1370), .Y(n1357) );
  NOR2X1 U1428 ( .A(n1371), .B(n1372), .Y(n1370) );
  OAI22X1 U1429 ( .A(n1236), .B(n11688), .C(n1238), .D(n11678), .Y(n1372) );
  OAI22X1 U1430 ( .A(n1240), .B(n11698), .C(n1242), .D(n11696), .Y(n1371) );
  AOI22X1 U1431 ( .A(\U_1/U_1/U_1/memory[1][6] ), .B(n1244), .C(
        \U_1/U_1/U_1/memory[0][6] ), .D(n1245), .Y(n1369) );
  AOI22X1 U1432 ( .A(\U_1/U_1/U_1/memory[3][6] ), .B(n1246), .C(
        \U_1/U_1/U_1/memory[2][6] ), .D(n1247), .Y(n1368) );
  OAI21X1 U1434 ( .A(n10282), .B(n11836), .C(n1377), .Y(n7934) );
  OAI21X1 U1435 ( .A(n1378), .B(n1379), .C(n10282), .Y(n1377) );
  NAND3X1 U1437 ( .A(n1382), .B(n1383), .C(n1384), .Y(n1381) );
  NOR2X1 U1438 ( .A(n1385), .B(n1386), .Y(n1384) );
  OAI22X1 U1439 ( .A(n1183), .B(n11777), .C(n1185), .D(n11787), .Y(n1386) );
  OAI22X1 U1440 ( .A(n1187), .B(n11757), .C(n1189), .D(n11767), .Y(n1385) );
  AOI22X1 U1441 ( .A(\U_1/U_1/U_1/memory[26][5] ), .B(n1191), .C(
        \U_1/U_1/U_1/memory[27][5] ), .D(n1192), .Y(n1383) );
  AOI22X1 U1442 ( .A(\U_1/U_1/U_1/memory[24][5] ), .B(n1193), .C(
        \U_1/U_1/U_1/memory[25][5] ), .D(n1194), .Y(n1382) );
  NAND3X1 U1443 ( .A(n1391), .B(n1392), .C(n1393), .Y(n1380) );
  NOR2X1 U1444 ( .A(n1394), .B(n1395), .Y(n1393) );
  OAI22X1 U1445 ( .A(n1200), .B(n11817), .C(n1202), .D(n11824), .Y(n1395) );
  OAI22X1 U1446 ( .A(n1204), .B(n11797), .C(n1206), .D(n11807), .Y(n1394) );
  AOI22X1 U1447 ( .A(\U_1/U_1/U_1/memory[22][5] ), .B(n1208), .C(
        \U_1/U_1/U_1/memory[23][5] ), .D(n1209), .Y(n1392) );
  AOI22X1 U1448 ( .A(\U_1/U_1/U_1/memory[20][5] ), .B(n1210), .C(
        \U_1/U_1/U_1/memory[21][5] ), .D(n1211), .Y(n1391) );
  NAND3X1 U1450 ( .A(n1402), .B(n1403), .C(n1404), .Y(n1401) );
  NOR2X1 U1451 ( .A(n1405), .B(n1406), .Y(n1404) );
  OAI22X1 U1452 ( .A(n1219), .B(n11747), .C(n1221), .D(n11717), .Y(n1406) );
  OAI22X1 U1453 ( .A(n1223), .B(n11727), .C(n1225), .D(n11737), .Y(n1405) );
  AOI22X1 U1454 ( .A(\U_1/U_1/U_1/memory[14][5] ), .B(n1227), .C(
        \U_1/U_1/U_1/memory[15][5] ), .D(n1228), .Y(n1403) );
  AOI22X1 U1455 ( .A(\U_1/U_1/U_1/memory[12][5] ), .B(n1229), .C(
        \U_1/U_1/U_1/memory[13][5] ), .D(n1230), .Y(n1402) );
  NAND3X1 U1456 ( .A(n1411), .B(n1412), .C(n1413), .Y(n1400) );
  NOR2X1 U1457 ( .A(n1414), .B(n1415), .Y(n1413) );
  OAI22X1 U1458 ( .A(n1236), .B(n11687), .C(n1238), .D(n11677), .Y(n1415) );
  OAI22X1 U1459 ( .A(n1240), .B(n11705), .C(n1242), .D(n11695), .Y(n1414) );
  AOI22X1 U1460 ( .A(\U_1/U_1/U_1/memory[1][5] ), .B(n1244), .C(
        \U_1/U_1/U_1/memory[0][5] ), .D(n1245), .Y(n1412) );
  AOI22X1 U1461 ( .A(\U_1/U_1/U_1/memory[3][5] ), .B(n1246), .C(
        \U_1/U_1/U_1/memory[2][5] ), .D(n1247), .Y(n1411) );
  OAI21X1 U1463 ( .A(n10282), .B(n11835), .C(n1420), .Y(n7935) );
  OAI21X1 U1464 ( .A(n1421), .B(n1422), .C(n10282), .Y(n1420) );
  NAND3X1 U1466 ( .A(n1425), .B(n1426), .C(n1427), .Y(n1424) );
  NOR2X1 U1467 ( .A(n1428), .B(n1429), .Y(n1427) );
  OAI22X1 U1468 ( .A(n1183), .B(n11776), .C(n1185), .D(n11786), .Y(n1429) );
  OAI22X1 U1469 ( .A(n1187), .B(n11756), .C(n1189), .D(n11766), .Y(n1428) );
  AOI22X1 U1470 ( .A(\U_1/U_1/U_1/memory[26][4] ), .B(n1191), .C(
        \U_1/U_1/U_1/memory[27][4] ), .D(n1192), .Y(n1426) );
  AOI22X1 U1471 ( .A(\U_1/U_1/U_1/memory[24][4] ), .B(n1193), .C(
        \U_1/U_1/U_1/memory[25][4] ), .D(n1194), .Y(n1425) );
  NAND3X1 U1472 ( .A(n1434), .B(n1435), .C(n1436), .Y(n1423) );
  NOR2X1 U1473 ( .A(n1437), .B(n1438), .Y(n1436) );
  OAI22X1 U1474 ( .A(n1200), .B(n11816), .C(n1202), .D(n11823), .Y(n1438) );
  OAI22X1 U1475 ( .A(n1204), .B(n11796), .C(n1206), .D(n11806), .Y(n1437) );
  AOI22X1 U1476 ( .A(\U_1/U_1/U_1/memory[22][4] ), .B(n1208), .C(
        \U_1/U_1/U_1/memory[23][4] ), .D(n1209), .Y(n1435) );
  AOI22X1 U1477 ( .A(\U_1/U_1/U_1/memory[20][4] ), .B(n1210), .C(
        \U_1/U_1/U_1/memory[21][4] ), .D(n1211), .Y(n1434) );
  NAND3X1 U1479 ( .A(n1445), .B(n1446), .C(n1447), .Y(n1444) );
  NOR2X1 U1480 ( .A(n1448), .B(n1449), .Y(n1447) );
  OAI22X1 U1481 ( .A(n1219), .B(n11746), .C(n1221), .D(n11716), .Y(n1449) );
  OAI22X1 U1482 ( .A(n1223), .B(n11726), .C(n1225), .D(n11736), .Y(n1448) );
  AOI22X1 U1483 ( .A(\U_1/U_1/U_1/memory[14][4] ), .B(n1227), .C(
        \U_1/U_1/U_1/memory[15][4] ), .D(n1228), .Y(n1446) );
  AOI22X1 U1484 ( .A(\U_1/U_1/U_1/memory[12][4] ), .B(n1229), .C(
        \U_1/U_1/U_1/memory[13][4] ), .D(n1230), .Y(n1445) );
  NAND3X1 U1485 ( .A(n1454), .B(n1455), .C(n1456), .Y(n1443) );
  NOR2X1 U1486 ( .A(n1457), .B(n1458), .Y(n1456) );
  OAI22X1 U1487 ( .A(n1236), .B(n11686), .C(n1238), .D(n11676), .Y(n1458) );
  OAI22X1 U1488 ( .A(n1240), .B(n11704), .C(n1242), .D(n11694), .Y(n1457) );
  AOI22X1 U1489 ( .A(\U_1/U_1/U_1/memory[1][4] ), .B(n1244), .C(
        \U_1/U_1/U_1/memory[0][4] ), .D(n1245), .Y(n1455) );
  AOI22X1 U1490 ( .A(\U_1/U_1/U_1/memory[3][4] ), .B(n1246), .C(
        \U_1/U_1/U_1/memory[2][4] ), .D(n1247), .Y(n1454) );
  OAI21X1 U1492 ( .A(n10282), .B(n11834), .C(n1463), .Y(n7936) );
  OAI21X1 U1493 ( .A(n1464), .B(n1465), .C(n10282), .Y(n1463) );
  NAND3X1 U1495 ( .A(n1468), .B(n1469), .C(n1470), .Y(n1467) );
  NOR2X1 U1496 ( .A(n1471), .B(n1472), .Y(n1470) );
  OAI22X1 U1497 ( .A(n1183), .B(n11775), .C(n1185), .D(n11785), .Y(n1472) );
  OAI22X1 U1498 ( .A(n1187), .B(n11755), .C(n1189), .D(n11765), .Y(n1471) );
  AOI22X1 U1499 ( .A(\U_1/U_1/U_1/memory[26][3] ), .B(n1191), .C(
        \U_1/U_1/U_1/memory[27][3] ), .D(n1192), .Y(n1469) );
  AOI22X1 U1500 ( .A(\U_1/U_1/U_1/memory[24][3] ), .B(n1193), .C(
        \U_1/U_1/U_1/memory[25][3] ), .D(n1194), .Y(n1468) );
  NAND3X1 U1501 ( .A(n1477), .B(n1478), .C(n1479), .Y(n1466) );
  NOR2X1 U1502 ( .A(n1480), .B(n1481), .Y(n1479) );
  OAI22X1 U1503 ( .A(n1200), .B(n11815), .C(n1202), .D(n11822), .Y(n1481) );
  OAI22X1 U1504 ( .A(n1204), .B(n11795), .C(n1206), .D(n11805), .Y(n1480) );
  AOI22X1 U1505 ( .A(\U_1/U_1/U_1/memory[22][3] ), .B(n1208), .C(
        \U_1/U_1/U_1/memory[23][3] ), .D(n1209), .Y(n1478) );
  AOI22X1 U1506 ( .A(\U_1/U_1/U_1/memory[20][3] ), .B(n1210), .C(
        \U_1/U_1/U_1/memory[21][3] ), .D(n1211), .Y(n1477) );
  NAND3X1 U1508 ( .A(n1488), .B(n1489), .C(n1490), .Y(n1487) );
  NOR2X1 U1509 ( .A(n1491), .B(n1492), .Y(n1490) );
  OAI22X1 U1510 ( .A(n1219), .B(n11745), .C(n1221), .D(n11715), .Y(n1492) );
  OAI22X1 U1511 ( .A(n1223), .B(n11725), .C(n1225), .D(n11735), .Y(n1491) );
  AOI22X1 U1512 ( .A(\U_1/U_1/U_1/memory[14][3] ), .B(n1227), .C(
        \U_1/U_1/U_1/memory[15][3] ), .D(n1228), .Y(n1489) );
  AOI22X1 U1513 ( .A(\U_1/U_1/U_1/memory[12][3] ), .B(n1229), .C(
        \U_1/U_1/U_1/memory[13][3] ), .D(n1230), .Y(n1488) );
  NAND3X1 U1514 ( .A(n1497), .B(n1498), .C(n1499), .Y(n1486) );
  NOR2X1 U1515 ( .A(n1500), .B(n1501), .Y(n1499) );
  OAI22X1 U1516 ( .A(n1236), .B(n11685), .C(n1238), .D(n11675), .Y(n1501) );
  OAI22X1 U1517 ( .A(n1240), .B(n11703), .C(n1242), .D(n11693), .Y(n1500) );
  AOI22X1 U1518 ( .A(\U_1/U_1/U_1/memory[1][3] ), .B(n1244), .C(
        \U_1/U_1/U_1/memory[0][3] ), .D(n1245), .Y(n1498) );
  AOI22X1 U1519 ( .A(\U_1/U_1/U_1/memory[3][3] ), .B(n1246), .C(
        \U_1/U_1/U_1/memory[2][3] ), .D(n1247), .Y(n1497) );
  OAI21X1 U1521 ( .A(n10282), .B(n11833), .C(n1506), .Y(n7937) );
  OAI21X1 U1522 ( .A(n1507), .B(n1508), .C(n10282), .Y(n1506) );
  NAND3X1 U1524 ( .A(n1511), .B(n1512), .C(n1513), .Y(n1510) );
  NOR2X1 U1525 ( .A(n1514), .B(n1515), .Y(n1513) );
  OAI22X1 U1526 ( .A(n1183), .B(n11774), .C(n1185), .D(n11784), .Y(n1515) );
  OAI22X1 U1527 ( .A(n1187), .B(n11754), .C(n1189), .D(n11764), .Y(n1514) );
  AOI22X1 U1528 ( .A(\U_1/U_1/U_1/memory[26][2] ), .B(n1191), .C(
        \U_1/U_1/U_1/memory[27][2] ), .D(n1192), .Y(n1512) );
  AOI22X1 U1529 ( .A(\U_1/U_1/U_1/memory[24][2] ), .B(n1193), .C(
        \U_1/U_1/U_1/memory[25][2] ), .D(n1194), .Y(n1511) );
  NAND3X1 U1530 ( .A(n1520), .B(n1521), .C(n1522), .Y(n1509) );
  NOR2X1 U1531 ( .A(n1523), .B(n1524), .Y(n1522) );
  OAI22X1 U1532 ( .A(n1200), .B(n11814), .C(n1202), .D(n11829), .Y(n1524) );
  OAI22X1 U1533 ( .A(n1204), .B(n11794), .C(n1206), .D(n11804), .Y(n1523) );
  AOI22X1 U1534 ( .A(\U_1/U_1/U_1/memory[22][2] ), .B(n1208), .C(
        \U_1/U_1/U_1/memory[23][2] ), .D(n1209), .Y(n1521) );
  AOI22X1 U1535 ( .A(\U_1/U_1/U_1/memory[20][2] ), .B(n1210), .C(
        \U_1/U_1/U_1/memory[21][2] ), .D(n1211), .Y(n1520) );
  NAND3X1 U1537 ( .A(n1531), .B(n1532), .C(n1533), .Y(n1530) );
  NOR2X1 U1538 ( .A(n1534), .B(n1535), .Y(n1533) );
  OAI22X1 U1539 ( .A(n1219), .B(n11744), .C(n1221), .D(n11714), .Y(n1535) );
  OAI22X1 U1540 ( .A(n1223), .B(n11724), .C(n1225), .D(n11734), .Y(n1534) );
  AOI22X1 U1541 ( .A(\U_1/U_1/U_1/memory[14][2] ), .B(n1227), .C(
        \U_1/U_1/U_1/memory[15][2] ), .D(n1228), .Y(n1532) );
  AOI22X1 U1542 ( .A(\U_1/U_1/U_1/memory[12][2] ), .B(n1229), .C(
        \U_1/U_1/U_1/memory[13][2] ), .D(n1230), .Y(n1531) );
  NAND3X1 U1543 ( .A(n1540), .B(n1541), .C(n1542), .Y(n1529) );
  NOR2X1 U1544 ( .A(n1543), .B(n1544), .Y(n1542) );
  OAI22X1 U1545 ( .A(n1236), .B(n11684), .C(n1238), .D(n11674), .Y(n1544) );
  OAI22X1 U1546 ( .A(n1240), .B(n11702), .C(n1242), .D(n11692), .Y(n1543) );
  AOI22X1 U1547 ( .A(\U_1/U_1/U_1/memory[1][2] ), .B(n1244), .C(
        \U_1/U_1/U_1/memory[0][2] ), .D(n1245), .Y(n1541) );
  AOI22X1 U1548 ( .A(\U_1/U_1/U_1/memory[3][2] ), .B(n1246), .C(
        \U_1/U_1/U_1/memory[2][2] ), .D(n1247), .Y(n1540) );
  OAI21X1 U1550 ( .A(n10282), .B(n11832), .C(n1549), .Y(n7938) );
  OAI21X1 U1551 ( .A(n1550), .B(n1551), .C(n10282), .Y(n1549) );
  NAND3X1 U1553 ( .A(n1554), .B(n1555), .C(n1556), .Y(n1553) );
  NOR2X1 U1554 ( .A(n1557), .B(n1558), .Y(n1556) );
  OAI22X1 U1555 ( .A(n1183), .B(n11773), .C(n1185), .D(n11783), .Y(n1558) );
  OAI22X1 U1556 ( .A(n1187), .B(n11753), .C(n1189), .D(n11763), .Y(n1557) );
  AOI22X1 U1557 ( .A(\U_1/U_1/U_1/memory[26][1] ), .B(n1191), .C(
        \U_1/U_1/U_1/memory[27][1] ), .D(n1192), .Y(n1555) );
  AOI22X1 U1558 ( .A(\U_1/U_1/U_1/memory[24][1] ), .B(n1193), .C(
        \U_1/U_1/U_1/memory[25][1] ), .D(n1194), .Y(n1554) );
  NAND3X1 U1559 ( .A(n1563), .B(n1564), .C(n1565), .Y(n1552) );
  NOR2X1 U1560 ( .A(n1566), .B(n1567), .Y(n1565) );
  OAI22X1 U1561 ( .A(n1200), .B(n11813), .C(n1202), .D(n11828), .Y(n1567) );
  OAI22X1 U1562 ( .A(n1204), .B(n11793), .C(n1206), .D(n11803), .Y(n1566) );
  AOI22X1 U1563 ( .A(\U_1/U_1/U_1/memory[22][1] ), .B(n1208), .C(
        \U_1/U_1/U_1/memory[23][1] ), .D(n1209), .Y(n1564) );
  AOI22X1 U1564 ( .A(\U_1/U_1/U_1/memory[20][1] ), .B(n1210), .C(
        \U_1/U_1/U_1/memory[21][1] ), .D(n1211), .Y(n1563) );
  NAND3X1 U1566 ( .A(n1574), .B(n1575), .C(n1576), .Y(n1573) );
  NOR2X1 U1567 ( .A(n1577), .B(n1578), .Y(n1576) );
  OAI22X1 U1568 ( .A(n1219), .B(n11743), .C(n1221), .D(n11713), .Y(n1578) );
  OAI22X1 U1569 ( .A(n1223), .B(n11723), .C(n1225), .D(n11733), .Y(n1577) );
  AOI22X1 U1570 ( .A(\U_1/U_1/U_1/memory[14][1] ), .B(n1227), .C(
        \U_1/U_1/U_1/memory[15][1] ), .D(n1228), .Y(n1575) );
  AOI22X1 U1571 ( .A(\U_1/U_1/U_1/memory[12][1] ), .B(n1229), .C(
        \U_1/U_1/U_1/memory[13][1] ), .D(n1230), .Y(n1574) );
  NAND3X1 U1572 ( .A(n1583), .B(n1584), .C(n1585), .Y(n1572) );
  NOR2X1 U1573 ( .A(n1586), .B(n1587), .Y(n1585) );
  OAI22X1 U1574 ( .A(n1236), .B(n11683), .C(n1238), .D(n11673), .Y(n1587) );
  OAI22X1 U1575 ( .A(n1240), .B(n11701), .C(n1242), .D(n11691), .Y(n1586) );
  AOI22X1 U1576 ( .A(\U_1/U_1/U_1/memory[1][1] ), .B(n1244), .C(
        \U_1/U_1/U_1/memory[0][1] ), .D(n1245), .Y(n1584) );
  AOI22X1 U1577 ( .A(\U_1/U_1/U_1/memory[3][1] ), .B(n1246), .C(
        \U_1/U_1/U_1/memory[2][1] ), .D(n1247), .Y(n1583) );
  OAI21X1 U1579 ( .A(n10282), .B(n11831), .C(n1592), .Y(n7939) );
  OAI21X1 U1580 ( .A(n1593), .B(n1594), .C(n10282), .Y(n1592) );
  NAND3X1 U1582 ( .A(n1597), .B(n1598), .C(n1599), .Y(n1596) );
  NOR2X1 U1583 ( .A(n1600), .B(n1601), .Y(n1599) );
  OAI22X1 U1584 ( .A(n1183), .B(n11772), .C(n1185), .D(n11782), .Y(n1601) );
  NAND2X1 U1585 ( .A(n11665), .B(n1605), .Y(n1185) );
  NAND2X1 U1586 ( .A(n11661), .B(n1605), .Y(n1183) );
  OAI22X1 U1587 ( .A(n1187), .B(n11752), .C(n1189), .D(n11762), .Y(n1600) );
  NAND2X1 U1588 ( .A(n11665), .B(n1609), .Y(n1189) );
  NAND2X1 U1589 ( .A(n11661), .B(n1609), .Y(n1187) );
  AOI22X1 U1590 ( .A(\U_1/U_1/U_1/memory[26][0] ), .B(n1191), .C(
        \U_1/U_1/U_1/memory[27][0] ), .D(n1192), .Y(n1598) );
  AOI22X1 U1593 ( .A(\U_1/U_1/U_1/memory[24][0] ), .B(n1193), .C(
        \U_1/U_1/U_1/memory[25][0] ), .D(n1194), .Y(n1597) );
  NAND3X1 U1596 ( .A(n9297), .B(\U_1/U_1/U_1/readptr[0] ), .C(
        \U_1/U_1/U_1/readptr[4] ), .Y(n1612) );
  NAND3X1 U1599 ( .A(n9297), .B(n9300), .C(\U_1/U_1/U_1/readptr[4] ), .Y(n1613) );
  NAND3X1 U1600 ( .A(n1615), .B(n1616), .C(n1617), .Y(n1595) );
  NOR2X1 U1601 ( .A(n1618), .B(n1619), .Y(n1617) );
  OAI22X1 U1602 ( .A(n1200), .B(n11812), .C(n1202), .D(n11827), .Y(n1619) );
  NAND2X1 U1603 ( .A(n11666), .B(n1610), .Y(n1202) );
  NAND2X1 U1604 ( .A(n11662), .B(n1610), .Y(n1200) );
  OAI22X1 U1605 ( .A(n1204), .B(n11792), .C(n1206), .D(n11802), .Y(n1618) );
  NAND2X1 U1606 ( .A(n11666), .B(n1611), .Y(n1206) );
  NAND2X1 U1607 ( .A(n11662), .B(n1611), .Y(n1204) );
  AOI22X1 U1608 ( .A(\U_1/U_1/U_1/memory[22][0] ), .B(n1208), .C(
        \U_1/U_1/U_1/memory[23][0] ), .D(n1209), .Y(n1616) );
  AOI22X1 U1611 ( .A(\U_1/U_1/U_1/memory[20][0] ), .B(n1210), .C(
        \U_1/U_1/U_1/memory[21][0] ), .D(n1211), .Y(n1615) );
  NAND3X1 U1614 ( .A(\U_1/U_1/U_1/readptr[0] ), .B(n9296), .C(
        \U_1/U_1/U_1/readptr[4] ), .Y(n1626) );
  NAND3X1 U1617 ( .A(n9300), .B(n9296), .C(\U_1/U_1/U_1/readptr[4] ), .Y(n1628) );
  NAND3X1 U1619 ( .A(n1631), .B(n1632), .C(n1633), .Y(n1630) );
  NOR2X1 U1620 ( .A(n1634), .B(n1635), .Y(n1633) );
  OAI22X1 U1621 ( .A(n1219), .B(n11742), .C(n1221), .D(n11712), .Y(n1635) );
  NAND2X1 U1622 ( .A(n11667), .B(n1610), .Y(n1221) );
  NAND2X1 U1623 ( .A(n11663), .B(n1610), .Y(n1219) );
  OAI22X1 U1624 ( .A(n1223), .B(n11722), .C(n1225), .D(n11732), .Y(n1634) );
  NAND2X1 U1625 ( .A(n11667), .B(n1611), .Y(n1225) );
  NAND2X1 U1626 ( .A(n11663), .B(n1611), .Y(n1223) );
  AOI22X1 U1627 ( .A(\U_1/U_1/U_1/memory[14][0] ), .B(n1227), .C(
        \U_1/U_1/U_1/memory[15][0] ), .D(n1228), .Y(n1632) );
  AOI22X1 U1630 ( .A(\U_1/U_1/U_1/memory[12][0] ), .B(n1229), .C(
        \U_1/U_1/U_1/memory[13][0] ), .D(n1230), .Y(n1631) );
  NAND3X1 U1633 ( .A(\U_1/U_1/U_1/readptr[0] ), .B(n9295), .C(n9297), .Y(n1642) );
  NAND3X1 U1636 ( .A(n9300), .B(n9295), .C(n9297), .Y(n1644) );
  NAND3X1 U1637 ( .A(n1645), .B(n1646), .C(n1647), .Y(n1629) );
  NOR2X1 U1638 ( .A(n1648), .B(n1649), .Y(n1647) );
  OAI22X1 U1639 ( .A(n1236), .B(n11682), .C(n1238), .D(n11672), .Y(n1649) );
  NAND2X1 U1640 ( .A(n1609), .B(n11664), .Y(n1238) );
  NAND2X1 U1641 ( .A(n1609), .B(n11668), .Y(n1236) );
  OAI22X1 U1643 ( .A(n1240), .B(n11700), .C(n1242), .D(n11690), .Y(n1648) );
  NAND2X1 U1644 ( .A(n1605), .B(n11664), .Y(n1242) );
  NAND2X1 U1645 ( .A(n1605), .B(n11668), .Y(n1240) );
  AOI22X1 U1647 ( .A(\U_1/U_1/U_1/memory[1][0] ), .B(n1244), .C(
        \U_1/U_1/U_1/memory[0][0] ), .D(n1245), .Y(n1646) );
  NOR2X1 U1650 ( .A(\U_1/U_1/U_1/readptr[1] ), .B(\U_1/U_1/U_1/readptr[2] ), 
        .Y(n1611) );
  AOI22X1 U1651 ( .A(\U_1/U_1/U_1/memory[3][0] ), .B(n1246), .C(
        \U_1/U_1/U_1/memory[2][0] ), .D(n1247), .Y(n1645) );
  NAND3X1 U1654 ( .A(n9296), .B(n9295), .C(n9300), .Y(n1657) );
  NAND3X1 U1658 ( .A(n9296), .B(n9295), .C(\U_1/U_1/U_1/readptr[0] ), .Y(n1658) );
  NOR2X1 U1661 ( .A(n9299), .B(\U_1/U_1/U_1/readptr[2] ), .Y(n1610) );
  NAND3X1 U1665 ( .A(\U_1/U_1/U_1/N195 ), .B(n9534), .C(n9318), .Y(n1659) );
  AOI22X1 U1667 ( .A(n10280), .B(\U_1/U_1/U_1/memory[0][7] ), .C(n9317), .D(
        n1662), .Y(n1660) );
  AOI22X1 U1669 ( .A(n10280), .B(\U_1/U_1/U_1/memory[0][6] ), .C(n1662), .D(
        \U_1/RCV_DATA [6]), .Y(n1663) );
  AOI22X1 U1671 ( .A(n10280), .B(\U_1/U_1/U_1/memory[0][5] ), .C(n1662), .D(
        n9313), .Y(n1664) );
  AOI22X1 U1673 ( .A(n10280), .B(\U_1/U_1/U_1/memory[0][4] ), .C(n1662), .D(
        n9311), .Y(n1665) );
  AOI22X1 U1675 ( .A(n10280), .B(\U_1/U_1/U_1/memory[0][3] ), .C(n1662), .D(
        n9309), .Y(n1666) );
  AOI22X1 U1677 ( .A(n10280), .B(\U_1/U_1/U_1/memory[0][2] ), .C(n1662), .D(
        n9307), .Y(n1667) );
  AOI22X1 U1679 ( .A(n10280), .B(\U_1/U_1/U_1/memory[0][1] ), .C(n1662), .D(
        n9305), .Y(n1668) );
  AOI22X1 U1681 ( .A(n10280), .B(\U_1/U_1/U_1/memory[0][0] ), .C(n1662), .D(
        n9303), .Y(n1669) );
  AOI22X1 U1683 ( .A(n10271), .B(\U_1/U_1/U_1/memory[1][7] ), .C(
        \U_1/RCV_DATA [7]), .D(n1672), .Y(n1670) );
  AOI22X1 U1685 ( .A(n10271), .B(\U_1/U_1/U_1/memory[1][6] ), .C(
        \U_1/RCV_DATA [6]), .D(n1672), .Y(n1673) );
  AOI22X1 U1687 ( .A(n10271), .B(\U_1/U_1/U_1/memory[1][5] ), .C(
        \U_1/RCV_DATA [5]), .D(n1672), .Y(n1674) );
  AOI22X1 U1689 ( .A(n10271), .B(\U_1/U_1/U_1/memory[1][4] ), .C(n9311), .D(
        n1672), .Y(n1675) );
  AOI22X1 U1691 ( .A(n10271), .B(\U_1/U_1/U_1/memory[1][3] ), .C(n9309), .D(
        n1672), .Y(n1676) );
  AOI22X1 U1693 ( .A(n10271), .B(\U_1/U_1/U_1/memory[1][2] ), .C(
        \U_1/RCV_DATA [2]), .D(n1672), .Y(n1677) );
  AOI22X1 U1695 ( .A(n10271), .B(\U_1/U_1/U_1/memory[1][1] ), .C(
        \U_1/RCV_DATA [1]), .D(n1672), .Y(n1678) );
  AOI22X1 U1697 ( .A(n10271), .B(\U_1/U_1/U_1/memory[1][0] ), .C(n9303), .D(
        n1672), .Y(n1679) );
  AOI22X1 U1699 ( .A(n10262), .B(\U_1/U_1/U_1/memory[2][7] ), .C(n9317), .D(
        n1682), .Y(n1680) );
  AOI22X1 U1701 ( .A(n10262), .B(\U_1/U_1/U_1/memory[2][6] ), .C(
        \U_1/RCV_DATA [6]), .D(n1682), .Y(n1683) );
  AOI22X1 U1703 ( .A(n10262), .B(\U_1/U_1/U_1/memory[2][5] ), .C(n9313), .D(
        n1682), .Y(n1684) );
  AOI22X1 U1705 ( .A(n10262), .B(\U_1/U_1/U_1/memory[2][4] ), .C(n9311), .D(
        n1682), .Y(n1685) );
  AOI22X1 U1707 ( .A(n10262), .B(\U_1/U_1/U_1/memory[2][3] ), .C(n9309), .D(
        n1682), .Y(n1686) );
  AOI22X1 U1709 ( .A(n10262), .B(\U_1/U_1/U_1/memory[2][2] ), .C(n9307), .D(
        n1682), .Y(n1687) );
  AOI22X1 U1711 ( .A(n10262), .B(\U_1/U_1/U_1/memory[2][1] ), .C(n9305), .D(
        n1682), .Y(n1688) );
  AOI22X1 U1713 ( .A(n10262), .B(\U_1/U_1/U_1/memory[2][0] ), .C(n9303), .D(
        n1682), .Y(n1689) );
  AOI22X1 U1715 ( .A(n10253), .B(\U_1/U_1/U_1/memory[3][7] ), .C(
        \U_1/RCV_DATA [7]), .D(n1692), .Y(n1690) );
  AOI22X1 U1717 ( .A(n10253), .B(\U_1/U_1/U_1/memory[3][6] ), .C(
        \U_1/RCV_DATA [6]), .D(n1692), .Y(n1693) );
  AOI22X1 U1719 ( .A(n10253), .B(\U_1/U_1/U_1/memory[3][5] ), .C(
        \U_1/RCV_DATA [5]), .D(n1692), .Y(n1694) );
  AOI22X1 U1721 ( .A(n10253), .B(\U_1/U_1/U_1/memory[3][4] ), .C(n9311), .D(
        n1692), .Y(n1695) );
  AOI22X1 U1723 ( .A(n10253), .B(\U_1/U_1/U_1/memory[3][3] ), .C(n9309), .D(
        n1692), .Y(n1696) );
  AOI22X1 U1725 ( .A(n10253), .B(\U_1/U_1/U_1/memory[3][2] ), .C(
        \U_1/RCV_DATA [2]), .D(n1692), .Y(n1697) );
  AOI22X1 U1727 ( .A(n10253), .B(\U_1/U_1/U_1/memory[3][1] ), .C(
        \U_1/RCV_DATA [1]), .D(n1692), .Y(n1698) );
  AOI22X1 U1729 ( .A(n10253), .B(\U_1/U_1/U_1/memory[3][0] ), .C(n9303), .D(
        n1692), .Y(n1699) );
  OAI22X1 U1730 ( .A(n1700), .B(n11679), .C(n9316), .D(n10244), .Y(n7972) );
  OAI22X1 U1732 ( .A(n1700), .B(n11678), .C(n9314), .D(n10244), .Y(n7973) );
  OAI22X1 U1734 ( .A(n1700), .B(n11677), .C(n9312), .D(n10244), .Y(n7974) );
  OAI22X1 U1736 ( .A(n1700), .B(n11676), .C(n9310), .D(n10244), .Y(n7975) );
  OAI22X1 U1738 ( .A(n1700), .B(n11675), .C(n9308), .D(n10244), .Y(n7976) );
  OAI22X1 U1740 ( .A(n1700), .B(n11674), .C(n9306), .D(n10244), .Y(n7977) );
  OAI22X1 U1742 ( .A(n1700), .B(n11673), .C(n9304), .D(n10244), .Y(n7978) );
  OAI22X1 U1744 ( .A(n1700), .B(n11672), .C(n9302), .D(n10244), .Y(n7979) );
  OAI22X1 U1746 ( .A(n1710), .B(n11689), .C(n9316), .D(n10243), .Y(n7980) );
  OAI22X1 U1748 ( .A(n1710), .B(n11688), .C(n9314), .D(n10243), .Y(n7981) );
  OAI22X1 U1750 ( .A(n1710), .B(n11687), .C(n9312), .D(n10243), .Y(n7982) );
  OAI22X1 U1752 ( .A(n1710), .B(n11686), .C(n9310), .D(n10243), .Y(n7983) );
  OAI22X1 U1754 ( .A(n1710), .B(n11685), .C(n9308), .D(n10243), .Y(n7984) );
  OAI22X1 U1756 ( .A(n1710), .B(n11684), .C(n9306), .D(n10243), .Y(n7985) );
  OAI22X1 U1758 ( .A(n1710), .B(n11683), .C(n9304), .D(n10243), .Y(n7986) );
  OAI22X1 U1760 ( .A(n1710), .B(n11682), .C(n9302), .D(n10243), .Y(n7987) );
  OAI22X1 U1762 ( .A(n1712), .B(n11697), .C(n9316), .D(n10242), .Y(n7988) );
  OAI22X1 U1764 ( .A(n1712), .B(n11696), .C(n9314), .D(n10242), .Y(n7989) );
  OAI22X1 U1766 ( .A(n1712), .B(n11695), .C(n9312), .D(n10242), .Y(n7990) );
  OAI22X1 U1768 ( .A(n1712), .B(n11694), .C(n9310), .D(n10242), .Y(n7991) );
  OAI22X1 U1770 ( .A(n1712), .B(n11693), .C(n9308), .D(n10242), .Y(n7992) );
  OAI22X1 U1772 ( .A(n1712), .B(n11692), .C(n9306), .D(n10242), .Y(n7993) );
  OAI22X1 U1774 ( .A(n1712), .B(n11691), .C(n9304), .D(n10242), .Y(n7994) );
  OAI22X1 U1776 ( .A(n1712), .B(n11690), .C(n9302), .D(n10242), .Y(n7995) );
  OAI22X1 U1778 ( .A(n1714), .B(n11705), .C(n9312), .D(n10241), .Y(n7996) );
  OAI22X1 U1780 ( .A(n1714), .B(n11704), .C(n9310), .D(n10241), .Y(n7997) );
  OAI22X1 U1782 ( .A(n1714), .B(n11703), .C(n9308), .D(n10241), .Y(n7998) );
  OAI22X1 U1784 ( .A(n1714), .B(n11702), .C(n9306), .D(n10241), .Y(n7999) );
  OAI22X1 U1786 ( .A(n1714), .B(n11701), .C(n9304), .D(n10241), .Y(n8000) );
  OAI22X1 U1788 ( .A(n1714), .B(n11700), .C(n9302), .D(n10241), .Y(n8001) );
  OAI22X1 U1790 ( .A(n1714), .B(n11699), .C(n9316), .D(n10241), .Y(n8002) );
  OAI22X1 U1792 ( .A(n1714), .B(n11698), .C(n9314), .D(n10241), .Y(n8003) );
  OAI22X1 U1794 ( .A(n9274), .B(n11729), .C(n9316), .D(n10239), .Y(n8004) );
  OAI22X1 U1796 ( .A(n9274), .B(n11728), .C(n9314), .D(n10239), .Y(n8005) );
  OAI22X1 U1798 ( .A(n9274), .B(n11727), .C(n9312), .D(n10239), .Y(n8006) );
  OAI22X1 U1800 ( .A(n9274), .B(n11726), .C(n9310), .D(n10239), .Y(n8007) );
  OAI22X1 U1802 ( .A(n9274), .B(n11725), .C(n9308), .D(n10239), .Y(n8008) );
  OAI22X1 U1804 ( .A(n9274), .B(n11724), .C(n9306), .D(n10239), .Y(n8009) );
  OAI22X1 U1806 ( .A(n9274), .B(n11723), .C(n9304), .D(n10239), .Y(n8010) );
  OAI22X1 U1808 ( .A(n9274), .B(n11722), .C(n9302), .D(n10239), .Y(n8011) );
  OAI22X1 U1810 ( .A(n9273), .B(n11739), .C(n9316), .D(n10238), .Y(n8012) );
  OAI22X1 U1812 ( .A(n9273), .B(n11738), .C(n9314), .D(n10238), .Y(n8013) );
  OAI22X1 U1814 ( .A(n9273), .B(n11737), .C(n9312), .D(n10238), .Y(n8014) );
  OAI22X1 U1816 ( .A(n9273), .B(n11736), .C(n9310), .D(n10238), .Y(n8015) );
  OAI22X1 U1818 ( .A(n9273), .B(n11735), .C(n9308), .D(n10238), .Y(n8016) );
  OAI22X1 U1820 ( .A(n9273), .B(n11734), .C(n9306), .D(n10238), .Y(n8017) );
  OAI22X1 U1822 ( .A(n9273), .B(n11733), .C(n9304), .D(n10238), .Y(n8018) );
  OAI22X1 U1824 ( .A(n9273), .B(n11732), .C(n9302), .D(n10238), .Y(n8019) );
  OAI22X1 U1826 ( .A(n9272), .B(n11749), .C(n9316), .D(n10237), .Y(n8020) );
  OAI22X1 U1828 ( .A(n9272), .B(n11748), .C(n9314), .D(n10237), .Y(n8021) );
  OAI22X1 U1830 ( .A(n9272), .B(n11747), .C(n9312), .D(n10237), .Y(n8022) );
  OAI22X1 U1832 ( .A(n9272), .B(n11746), .C(n9310), .D(n10237), .Y(n8023) );
  OAI22X1 U1834 ( .A(n9272), .B(n11745), .C(n9308), .D(n10237), .Y(n8024) );
  OAI22X1 U1836 ( .A(n9272), .B(n11744), .C(n9306), .D(n10237), .Y(n8025) );
  OAI22X1 U1838 ( .A(n9272), .B(n11743), .C(n9304), .D(n10237), .Y(n8026) );
  OAI22X1 U1840 ( .A(n9272), .B(n11742), .C(n9302), .D(n10237), .Y(n8027) );
  OAI22X1 U1842 ( .A(n9275), .B(n11719), .C(n9316), .D(n10240), .Y(n8028) );
  OAI22X1 U1844 ( .A(n9275), .B(n11718), .C(n9314), .D(n10240), .Y(n8029) );
  OAI22X1 U1846 ( .A(n9275), .B(n11717), .C(n9312), .D(n10240), .Y(n8030) );
  OAI22X1 U1848 ( .A(n9275), .B(n11716), .C(n9310), .D(n10240), .Y(n8031) );
  OAI22X1 U1850 ( .A(n9275), .B(n11715), .C(n9308), .D(n10240), .Y(n8032) );
  OAI22X1 U1852 ( .A(n9275), .B(n11714), .C(n9306), .D(n10240), .Y(n8033) );
  OAI22X1 U1854 ( .A(n9275), .B(n11713), .C(n9304), .D(n10240), .Y(n8034) );
  OAI22X1 U1856 ( .A(n9275), .B(n11712), .C(n9302), .D(n10240), .Y(n8035) );
  NOR2X1 U1859 ( .A(n1724), .B(n1725), .Y(n1722) );
  AOI22X1 U1861 ( .A(n10236), .B(\U_1/U_1/U_1/memory[12][7] ), .C(n9317), .D(
        n9271), .Y(n1726) );
  AOI22X1 U1863 ( .A(n10236), .B(\U_1/U_1/U_1/memory[12][6] ), .C(
        \U_1/RCV_DATA [6]), .D(n9271), .Y(n1729) );
  AOI22X1 U1865 ( .A(n10236), .B(\U_1/U_1/U_1/memory[12][5] ), .C(n9313), .D(
        n9271), .Y(n1730) );
  AOI22X1 U1867 ( .A(n10236), .B(\U_1/U_1/U_1/memory[12][4] ), .C(n9311), .D(
        n9271), .Y(n1731) );
  AOI22X1 U1869 ( .A(n10236), .B(\U_1/U_1/U_1/memory[12][3] ), .C(n9309), .D(
        n9271), .Y(n1732) );
  AOI22X1 U1871 ( .A(n10236), .B(\U_1/U_1/U_1/memory[12][2] ), .C(n9307), .D(
        n9271), .Y(n1733) );
  AOI22X1 U1873 ( .A(n10236), .B(\U_1/U_1/U_1/memory[12][1] ), .C(n9305), .D(
        n9271), .Y(n1734) );
  AOI22X1 U1875 ( .A(n10236), .B(\U_1/U_1/U_1/memory[12][0] ), .C(n9303), .D(
        n9271), .Y(n1735) );
  AOI22X1 U1877 ( .A(n10227), .B(\U_1/U_1/U_1/memory[13][7] ), .C(
        \U_1/RCV_DATA [7]), .D(n9270), .Y(n1736) );
  AOI22X1 U1879 ( .A(n10227), .B(\U_1/U_1/U_1/memory[13][6] ), .C(
        \U_1/RCV_DATA [6]), .D(n9270), .Y(n1739) );
  AOI22X1 U1881 ( .A(n10227), .B(\U_1/U_1/U_1/memory[13][5] ), .C(
        \U_1/RCV_DATA [5]), .D(n9270), .Y(n1740) );
  AOI22X1 U1883 ( .A(n10227), .B(\U_1/U_1/U_1/memory[13][4] ), .C(n9311), .D(
        n9270), .Y(n1741) );
  AOI22X1 U1885 ( .A(n10227), .B(\U_1/U_1/U_1/memory[13][3] ), .C(n9309), .D(
        n9270), .Y(n1742) );
  AOI22X1 U1887 ( .A(n10227), .B(\U_1/U_1/U_1/memory[13][2] ), .C(
        \U_1/RCV_DATA [2]), .D(n9270), .Y(n1743) );
  AOI22X1 U1889 ( .A(n10227), .B(\U_1/U_1/U_1/memory[13][1] ), .C(
        \U_1/RCV_DATA [1]), .D(n9270), .Y(n1744) );
  AOI22X1 U1891 ( .A(n10227), .B(\U_1/U_1/U_1/memory[13][0] ), .C(n9303), .D(
        n9270), .Y(n1745) );
  AOI22X1 U1893 ( .A(n10218), .B(\U_1/U_1/U_1/memory[14][7] ), .C(n9317), .D(
        n9269), .Y(n1746) );
  AOI22X1 U1895 ( .A(n10218), .B(\U_1/U_1/U_1/memory[14][6] ), .C(
        \U_1/RCV_DATA [6]), .D(n9269), .Y(n1749) );
  AOI22X1 U1897 ( .A(n10218), .B(\U_1/U_1/U_1/memory[14][5] ), .C(n9313), .D(
        n9269), .Y(n1750) );
  AOI22X1 U1899 ( .A(n10218), .B(\U_1/U_1/U_1/memory[14][4] ), .C(n9311), .D(
        n9269), .Y(n1751) );
  AOI22X1 U1901 ( .A(n10218), .B(\U_1/U_1/U_1/memory[14][3] ), .C(n9309), .D(
        n9269), .Y(n1752) );
  AOI22X1 U1903 ( .A(n10218), .B(\U_1/U_1/U_1/memory[14][2] ), .C(n9307), .D(
        n9269), .Y(n1753) );
  AOI22X1 U1905 ( .A(n10218), .B(\U_1/U_1/U_1/memory[14][1] ), .C(n9305), .D(
        n9269), .Y(n1754) );
  AOI22X1 U1907 ( .A(n10218), .B(\U_1/U_1/U_1/memory[14][0] ), .C(n9303), .D(
        n9269), .Y(n1755) );
  AOI22X1 U1909 ( .A(n10209), .B(\U_1/U_1/U_1/memory[15][7] ), .C(
        \U_1/RCV_DATA [7]), .D(n9268), .Y(n1756) );
  AOI22X1 U1911 ( .A(n10209), .B(\U_1/U_1/U_1/memory[15][6] ), .C(n9315), .D(
        n9268), .Y(n1759) );
  AOI22X1 U1913 ( .A(n10209), .B(\U_1/U_1/U_1/memory[15][5] ), .C(
        \U_1/RCV_DATA [5]), .D(n9268), .Y(n1760) );
  AOI22X1 U1915 ( .A(n10209), .B(\U_1/U_1/U_1/memory[15][4] ), .C(
        \U_1/RCV_DATA [4]), .D(n9268), .Y(n1761) );
  AOI22X1 U1917 ( .A(n10209), .B(\U_1/U_1/U_1/memory[15][3] ), .C(
        \U_1/RCV_DATA [3]), .D(n9268), .Y(n1762) );
  AOI22X1 U1919 ( .A(n10209), .B(\U_1/U_1/U_1/memory[15][2] ), .C(
        \U_1/RCV_DATA [2]), .D(n9268), .Y(n1763) );
  AOI22X1 U1921 ( .A(n10209), .B(\U_1/U_1/U_1/memory[15][1] ), .C(
        \U_1/RCV_DATA [1]), .D(n9268), .Y(n1764) );
  AOI22X1 U1923 ( .A(n10209), .B(\U_1/U_1/U_1/memory[15][0] ), .C(
        \U_1/RCV_DATA [0]), .D(n9268), .Y(n1765) );
  OAI22X1 U1924 ( .A(n9267), .B(n11799), .C(n9316), .D(n10200), .Y(n8068) );
  OAI22X1 U1926 ( .A(n9267), .B(n11798), .C(n9314), .D(n10200), .Y(n8069) );
  OAI22X1 U1928 ( .A(n9267), .B(n11797), .C(n9312), .D(n10200), .Y(n8070) );
  OAI22X1 U1930 ( .A(n9267), .B(n11796), .C(n9310), .D(n10200), .Y(n8071) );
  OAI22X1 U1932 ( .A(n9267), .B(n11795), .C(n9308), .D(n10200), .Y(n8072) );
  OAI22X1 U1934 ( .A(n9267), .B(n11794), .C(n9306), .D(n10200), .Y(n8073) );
  OAI22X1 U1936 ( .A(n9267), .B(n11793), .C(n9304), .D(n10200), .Y(n8074) );
  OAI22X1 U1938 ( .A(n9267), .B(n11792), .C(n9302), .D(n10200), .Y(n8075) );
  OAI22X1 U1940 ( .A(n9266), .B(n11809), .C(n9316), .D(n10199), .Y(n8076) );
  OAI22X1 U1942 ( .A(n9266), .B(n11808), .C(n9314), .D(n10199), .Y(n8077) );
  OAI22X1 U1944 ( .A(n9266), .B(n11807), .C(n9312), .D(n10199), .Y(n8078) );
  OAI22X1 U1946 ( .A(n9266), .B(n11806), .C(n9310), .D(n10199), .Y(n8079) );
  OAI22X1 U1948 ( .A(n9266), .B(n11805), .C(n9308), .D(n10199), .Y(n8080) );
  OAI22X1 U1950 ( .A(n9266), .B(n11804), .C(n9306), .D(n10199), .Y(n8081) );
  OAI22X1 U1952 ( .A(n9266), .B(n11803), .C(n9304), .D(n10199), .Y(n8082) );
  OAI22X1 U1954 ( .A(n9266), .B(n11802), .C(n9302), .D(n10199), .Y(n8083) );
  OAI22X1 U1956 ( .A(n9265), .B(n11819), .C(n9316), .D(n10198), .Y(n8084) );
  OAI22X1 U1958 ( .A(n9265), .B(n11818), .C(n9314), .D(n10198), .Y(n8085) );
  OAI22X1 U1960 ( .A(n9265), .B(n11817), .C(n9312), .D(n10198), .Y(n8086) );
  OAI22X1 U1962 ( .A(n9265), .B(n11816), .C(n9310), .D(n10198), .Y(n8087) );
  OAI22X1 U1964 ( .A(n9265), .B(n11815), .C(n9308), .D(n10198), .Y(n8088) );
  OAI22X1 U1966 ( .A(n9265), .B(n11814), .C(n9306), .D(n10198), .Y(n8089) );
  OAI22X1 U1968 ( .A(n9265), .B(n11813), .C(n9304), .D(n10198), .Y(n8090) );
  OAI22X1 U1970 ( .A(n9265), .B(n11812), .C(n9302), .D(n10198), .Y(n8091) );
  OAI22X1 U1972 ( .A(n9264), .B(n11829), .C(n9306), .D(n10197), .Y(n8092) );
  OAI22X1 U1974 ( .A(n9264), .B(n11828), .C(n9304), .D(n10197), .Y(n8093) );
  OAI22X1 U1976 ( .A(n9264), .B(n11827), .C(n9302), .D(n10197), .Y(n8094) );
  OAI22X1 U1978 ( .A(n9264), .B(n11826), .C(n9316), .D(n10197), .Y(n8095) );
  OAI22X1 U1980 ( .A(n9264), .B(n11825), .C(n9314), .D(n10197), .Y(n8096) );
  OAI22X1 U1982 ( .A(n9264), .B(n11824), .C(n9312), .D(n10197), .Y(n8097) );
  OAI22X1 U1984 ( .A(n9264), .B(n11823), .C(n9310), .D(n10197), .Y(n8098) );
  OAI22X1 U1986 ( .A(n9264), .B(n11822), .C(n9308), .D(n10197), .Y(n8099) );
  AOI22X1 U1989 ( .A(n10196), .B(\U_1/U_1/U_1/memory[20][7] ), .C(n9317), .D(
        n9263), .Y(n1774) );
  AOI22X1 U1991 ( .A(n10196), .B(\U_1/U_1/U_1/memory[20][6] ), .C(n9315), .D(
        n9263), .Y(n1777) );
  AOI22X1 U1993 ( .A(n10196), .B(\U_1/U_1/U_1/memory[20][5] ), .C(n9313), .D(
        n9263), .Y(n1778) );
  AOI22X1 U1995 ( .A(n10196), .B(\U_1/U_1/U_1/memory[20][4] ), .C(
        \U_1/RCV_DATA [4]), .D(n9263), .Y(n1779) );
  AOI22X1 U1997 ( .A(n10196), .B(\U_1/U_1/U_1/memory[20][3] ), .C(
        \U_1/RCV_DATA [3]), .D(n9263), .Y(n1780) );
  AOI22X1 U1999 ( .A(n10196), .B(\U_1/U_1/U_1/memory[20][2] ), .C(n9307), .D(
        n9263), .Y(n1781) );
  AOI22X1 U2001 ( .A(n10196), .B(\U_1/U_1/U_1/memory[20][1] ), .C(n9305), .D(
        n9263), .Y(n1782) );
  AOI22X1 U2003 ( .A(n10196), .B(\U_1/U_1/U_1/memory[20][0] ), .C(
        \U_1/RCV_DATA [0]), .D(n9263), .Y(n1783) );
  AOI22X1 U2005 ( .A(n10187), .B(\U_1/U_1/U_1/memory[21][7] ), .C(
        \U_1/RCV_DATA [7]), .D(n9262), .Y(n1784) );
  AOI22X1 U2007 ( .A(n10187), .B(\U_1/U_1/U_1/memory[21][6] ), .C(n9315), .D(
        n9262), .Y(n1787) );
  AOI22X1 U2009 ( .A(n10187), .B(\U_1/U_1/U_1/memory[21][5] ), .C(
        \U_1/RCV_DATA [5]), .D(n9262), .Y(n1788) );
  AOI22X1 U2011 ( .A(n10187), .B(\U_1/U_1/U_1/memory[21][4] ), .C(
        \U_1/RCV_DATA [4]), .D(n9262), .Y(n1789) );
  AOI22X1 U2013 ( .A(n10187), .B(\U_1/U_1/U_1/memory[21][3] ), .C(
        \U_1/RCV_DATA [3]), .D(n9262), .Y(n1790) );
  AOI22X1 U2015 ( .A(n10187), .B(\U_1/U_1/U_1/memory[21][2] ), .C(
        \U_1/RCV_DATA [2]), .D(n9262), .Y(n1791) );
  AOI22X1 U2017 ( .A(n10187), .B(\U_1/U_1/U_1/memory[21][1] ), .C(
        \U_1/RCV_DATA [1]), .D(n9262), .Y(n1792) );
  AOI22X1 U2019 ( .A(n10187), .B(\U_1/U_1/U_1/memory[21][0] ), .C(
        \U_1/RCV_DATA [0]), .D(n9262), .Y(n1793) );
  AOI22X1 U2021 ( .A(n10178), .B(\U_1/U_1/U_1/memory[22][7] ), .C(n9317), .D(
        n9261), .Y(n1794) );
  AOI22X1 U2023 ( .A(n10178), .B(\U_1/U_1/U_1/memory[22][6] ), .C(n9315), .D(
        n9261), .Y(n1797) );
  AOI22X1 U2025 ( .A(n10178), .B(\U_1/U_1/U_1/memory[22][5] ), .C(n9313), .D(
        n9261), .Y(n1798) );
  AOI22X1 U2027 ( .A(n10178), .B(\U_1/U_1/U_1/memory[22][4] ), .C(
        \U_1/RCV_DATA [4]), .D(n9261), .Y(n1799) );
  AOI22X1 U2029 ( .A(n10178), .B(\U_1/U_1/U_1/memory[22][3] ), .C(
        \U_1/RCV_DATA [3]), .D(n9261), .Y(n1800) );
  AOI22X1 U2031 ( .A(n10178), .B(\U_1/U_1/U_1/memory[22][2] ), .C(n9307), .D(
        n9261), .Y(n1801) );
  AOI22X1 U2033 ( .A(n10178), .B(\U_1/U_1/U_1/memory[22][1] ), .C(n9305), .D(
        n9261), .Y(n1802) );
  AOI22X1 U2035 ( .A(n10178), .B(\U_1/U_1/U_1/memory[22][0] ), .C(
        \U_1/RCV_DATA [0]), .D(n9261), .Y(n1803) );
  AOI22X1 U2037 ( .A(n10169), .B(\U_1/U_1/U_1/memory[23][7] ), .C(
        \U_1/RCV_DATA [7]), .D(n9260), .Y(n1804) );
  AOI22X1 U2039 ( .A(n10169), .B(\U_1/U_1/U_1/memory[23][6] ), .C(n9315), .D(
        n9260), .Y(n1807) );
  AOI22X1 U2041 ( .A(n10169), .B(\U_1/U_1/U_1/memory[23][5] ), .C(
        \U_1/RCV_DATA [5]), .D(n9260), .Y(n1808) );
  AOI22X1 U2043 ( .A(n10169), .B(\U_1/U_1/U_1/memory[23][4] ), .C(
        \U_1/RCV_DATA [4]), .D(n9260), .Y(n1809) );
  AOI22X1 U2045 ( .A(n10169), .B(\U_1/U_1/U_1/memory[23][3] ), .C(
        \U_1/RCV_DATA [3]), .D(n9260), .Y(n1810) );
  AOI22X1 U2047 ( .A(n10169), .B(\U_1/U_1/U_1/memory[23][2] ), .C(
        \U_1/RCV_DATA [2]), .D(n9260), .Y(n1811) );
  AOI22X1 U2049 ( .A(n10169), .B(\U_1/U_1/U_1/memory[23][1] ), .C(
        \U_1/RCV_DATA [1]), .D(n9260), .Y(n1812) );
  AOI22X1 U2051 ( .A(n10169), .B(\U_1/U_1/U_1/memory[23][0] ), .C(
        \U_1/RCV_DATA [0]), .D(n9260), .Y(n1813) );
  AOI22X1 U2053 ( .A(n10160), .B(\U_1/U_1/U_1/memory[24][7] ), .C(n9317), .D(
        n9259), .Y(n1814) );
  AOI22X1 U2055 ( .A(n10160), .B(\U_1/U_1/U_1/memory[24][6] ), .C(n9315), .D(
        n9259), .Y(n1817) );
  AOI22X1 U2057 ( .A(n10160), .B(\U_1/U_1/U_1/memory[24][5] ), .C(n9313), .D(
        n9259), .Y(n1818) );
  AOI22X1 U2059 ( .A(n10160), .B(\U_1/U_1/U_1/memory[24][4] ), .C(
        \U_1/RCV_DATA [4]), .D(n9259), .Y(n1819) );
  AOI22X1 U2061 ( .A(n10160), .B(\U_1/U_1/U_1/memory[24][3] ), .C(
        \U_1/RCV_DATA [3]), .D(n9259), .Y(n1820) );
  AOI22X1 U2063 ( .A(n10160), .B(\U_1/U_1/U_1/memory[24][2] ), .C(n9307), .D(
        n9259), .Y(n1821) );
  AOI22X1 U2065 ( .A(n10160), .B(\U_1/U_1/U_1/memory[24][1] ), .C(n9305), .D(
        n9259), .Y(n1822) );
  AOI22X1 U2067 ( .A(n10160), .B(\U_1/U_1/U_1/memory[24][0] ), .C(
        \U_1/RCV_DATA [0]), .D(n9259), .Y(n1823) );
  AOI22X1 U2069 ( .A(n10151), .B(\U_1/U_1/U_1/memory[25][7] ), .C(
        \U_1/RCV_DATA [7]), .D(n9258), .Y(n1824) );
  AOI22X1 U2071 ( .A(n10151), .B(\U_1/U_1/U_1/memory[25][6] ), .C(n9315), .D(
        n9258), .Y(n1827) );
  AOI22X1 U2073 ( .A(n10151), .B(\U_1/U_1/U_1/memory[25][5] ), .C(
        \U_1/RCV_DATA [5]), .D(n9258), .Y(n1828) );
  AOI22X1 U2075 ( .A(n10151), .B(\U_1/U_1/U_1/memory[25][4] ), .C(
        \U_1/RCV_DATA [4]), .D(n9258), .Y(n1829) );
  AOI22X1 U2077 ( .A(n10151), .B(\U_1/U_1/U_1/memory[25][3] ), .C(
        \U_1/RCV_DATA [3]), .D(n9258), .Y(n1830) );
  AOI22X1 U2079 ( .A(n10151), .B(\U_1/U_1/U_1/memory[25][2] ), .C(
        \U_1/RCV_DATA [2]), .D(n9258), .Y(n1831) );
  AOI22X1 U2081 ( .A(n10151), .B(\U_1/U_1/U_1/memory[25][1] ), .C(
        \U_1/RCV_DATA [1]), .D(n9258), .Y(n1832) );
  AOI22X1 U2083 ( .A(n10151), .B(\U_1/U_1/U_1/memory[25][0] ), .C(
        \U_1/RCV_DATA [0]), .D(n9258), .Y(n1833) );
  AOI22X1 U2085 ( .A(n10142), .B(\U_1/U_1/U_1/memory[26][7] ), .C(n9317), .D(
        n9257), .Y(n1834) );
  AOI22X1 U2087 ( .A(n10142), .B(\U_1/U_1/U_1/memory[26][6] ), .C(n9315), .D(
        n9257), .Y(n1837) );
  AOI22X1 U2089 ( .A(n10142), .B(\U_1/U_1/U_1/memory[26][5] ), .C(n9313), .D(
        n9257), .Y(n1838) );
  AOI22X1 U2091 ( .A(n10142), .B(\U_1/U_1/U_1/memory[26][4] ), .C(n9311), .D(
        n9257), .Y(n1839) );
  AOI22X1 U2093 ( .A(n10142), .B(\U_1/U_1/U_1/memory[26][3] ), .C(n9309), .D(
        n9257), .Y(n1840) );
  AOI22X1 U2095 ( .A(n10142), .B(\U_1/U_1/U_1/memory[26][2] ), .C(n9307), .D(
        n9257), .Y(n1841) );
  AOI22X1 U2097 ( .A(n10142), .B(\U_1/U_1/U_1/memory[26][1] ), .C(n9305), .D(
        n9257), .Y(n1842) );
  AOI22X1 U2099 ( .A(n10142), .B(\U_1/U_1/U_1/memory[26][0] ), .C(n9303), .D(
        n9257), .Y(n1843) );
  AOI22X1 U2101 ( .A(n10133), .B(\U_1/U_1/U_1/memory[27][7] ), .C(n9317), .D(
        n9256), .Y(n1844) );
  AOI22X1 U2103 ( .A(n10133), .B(\U_1/U_1/U_1/memory[27][6] ), .C(n9315), .D(
        n9256), .Y(n1847) );
  AOI22X1 U2105 ( .A(n10133), .B(\U_1/U_1/U_1/memory[27][5] ), .C(n9313), .D(
        n9256), .Y(n1848) );
  AOI22X1 U2107 ( .A(n10133), .B(\U_1/U_1/U_1/memory[27][4] ), .C(n9311), .D(
        n9256), .Y(n1849) );
  AOI22X1 U2109 ( .A(n10133), .B(\U_1/U_1/U_1/memory[27][3] ), .C(n9309), .D(
        n9256), .Y(n1850) );
  AOI22X1 U2111 ( .A(n10133), .B(\U_1/U_1/U_1/memory[27][2] ), .C(n9307), .D(
        n9256), .Y(n1851) );
  AOI22X1 U2113 ( .A(n10133), .B(\U_1/U_1/U_1/memory[27][1] ), .C(n9305), .D(
        n9256), .Y(n1852) );
  AOI22X1 U2115 ( .A(n10133), .B(\U_1/U_1/U_1/memory[27][0] ), .C(n9303), .D(
        n9256), .Y(n1853) );
  OAI22X1 U2116 ( .A(n9255), .B(n11759), .C(n9316), .D(n10124), .Y(n8164) );
  OAI22X1 U2118 ( .A(n9255), .B(n11758), .C(n9314), .D(n10124), .Y(n8165) );
  OAI22X1 U2120 ( .A(n9255), .B(n11757), .C(n9312), .D(n10124), .Y(n8166) );
  OAI22X1 U2122 ( .A(n9255), .B(n11756), .C(n9310), .D(n10124), .Y(n8167) );
  OAI22X1 U2124 ( .A(n9255), .B(n11755), .C(n9308), .D(n10124), .Y(n8168) );
  OAI22X1 U2126 ( .A(n9255), .B(n11754), .C(n9306), .D(n10124), .Y(n8169) );
  OAI22X1 U2128 ( .A(n9255), .B(n11753), .C(n9304), .D(n10124), .Y(n8170) );
  OAI22X1 U2130 ( .A(n9255), .B(n11752), .C(n9302), .D(n10124), .Y(n8171) );
  OAI22X1 U2132 ( .A(n9254), .B(n11769), .C(n9316), .D(n10123), .Y(n8172) );
  OAI22X1 U2134 ( .A(n9254), .B(n11768), .C(n9314), .D(n10123), .Y(n8173) );
  OAI22X1 U2136 ( .A(n9254), .B(n11767), .C(n9312), .D(n10123), .Y(n8174) );
  OAI22X1 U2138 ( .A(n9254), .B(n11766), .C(n9310), .D(n10123), .Y(n8175) );
  OAI22X1 U2140 ( .A(n9254), .B(n11765), .C(n9308), .D(n10123), .Y(n8176) );
  OAI22X1 U2142 ( .A(n9254), .B(n11764), .C(n9306), .D(n10123), .Y(n8177) );
  OAI22X1 U2144 ( .A(n9254), .B(n11763), .C(n9304), .D(n10123), .Y(n8178) );
  OAI22X1 U2146 ( .A(n9254), .B(n11762), .C(n9302), .D(n10123), .Y(n8179) );
  OAI22X1 U2148 ( .A(n9253), .B(n11779), .C(n9316), .D(n10122), .Y(n8180) );
  OAI22X1 U2150 ( .A(n9253), .B(n11778), .C(n9314), .D(n10122), .Y(n8181) );
  OAI22X1 U2152 ( .A(n9253), .B(n11777), .C(n9312), .D(n10122), .Y(n8182) );
  OAI22X1 U2154 ( .A(n9253), .B(n11776), .C(n9310), .D(n10122), .Y(n8183) );
  OAI22X1 U2156 ( .A(n9253), .B(n11775), .C(n9308), .D(n10122), .Y(n8184) );
  OAI22X1 U2158 ( .A(n9253), .B(n11774), .C(n9306), .D(n10122), .Y(n8185) );
  OAI22X1 U2160 ( .A(n9253), .B(n11773), .C(n9304), .D(n10122), .Y(n8186) );
  OAI22X1 U2162 ( .A(n9253), .B(n11772), .C(n9302), .D(n10122), .Y(n8187) );
  OAI22X1 U2164 ( .A(n9252), .B(n11789), .C(n9316), .D(n10121), .Y(n8188) );
  OAI22X1 U2166 ( .A(n9252), .B(n11788), .C(n9314), .D(n10121), .Y(n8189) );
  OAI22X1 U2168 ( .A(n9252), .B(n11787), .C(n9312), .D(n10121), .Y(n8190) );
  OAI22X1 U2170 ( .A(n9252), .B(n11786), .C(n9310), .D(n10121), .Y(n8191) );
  OAI22X1 U2172 ( .A(n9252), .B(n11785), .C(n9308), .D(n10121), .Y(n8192) );
  OAI22X1 U2174 ( .A(n9252), .B(n11784), .C(n9306), .D(n10121), .Y(n8193) );
  OAI22X1 U2176 ( .A(n9252), .B(n11783), .C(n9304), .D(n10121), .Y(n8194) );
  OAI22X1 U2178 ( .A(n9252), .B(n11782), .C(n9302), .D(n10121), .Y(n8195) );
  AOI22X1 U2181 ( .A(n1863), .B(n11557), .C(\U_1/U_1/U_1/opcode[0][1] ), .D(
        n10073), .Y(n1862) );
  AOI22X1 U2183 ( .A(n9180), .B(n1863), .C(\U_1/U_1/U_1/opcode[0][0] ), .D(
        n10073), .Y(n1866) );
  OAI21X1 U2185 ( .A(n1868), .B(n1869), .C(n10280), .Y(n1863) );
  NOR2X1 U2187 ( .A(n1870), .B(n1871), .Y(n1662) );
  AOI22X1 U2189 ( .A(n1873), .B(n11557), .C(\U_1/U_1/U_1/opcode[1][1] ), .D(
        n10070), .Y(n1872) );
  AOI22X1 U2191 ( .A(n9180), .B(n1873), .C(\U_1/U_1/U_1/opcode[1][0] ), .D(
        n10070), .Y(n1875) );
  OAI21X1 U2193 ( .A(n1725), .B(n1869), .C(n10271), .Y(n1873) );
  NOR2X1 U2195 ( .A(n1876), .B(n1870), .Y(n1672) );
  AOI22X1 U2197 ( .A(n1878), .B(n11557), .C(\U_1/U_1/U_1/opcode[2][1] ), .D(
        n10067), .Y(n1877) );
  AOI22X1 U2199 ( .A(n9180), .B(n1878), .C(\U_1/U_1/U_1/opcode[2][0] ), .D(
        n10067), .Y(n1880) );
  OAI21X1 U2201 ( .A(n1881), .B(n1869), .C(n10262), .Y(n1878) );
  NOR2X1 U2203 ( .A(n1868), .B(n1870), .Y(n1682) );
  AOI22X1 U2205 ( .A(n1883), .B(n11557), .C(\U_1/U_1/U_1/opcode[3][1] ), .D(
        n10064), .Y(n1882) );
  AOI22X1 U2207 ( .A(n9180), .B(n1883), .C(\U_1/U_1/U_1/opcode[3][0] ), .D(
        n10064), .Y(n1885) );
  OAI21X1 U2209 ( .A(n1886), .B(n1869), .C(n10253), .Y(n1883) );
  NOR2X1 U2211 ( .A(n1725), .B(n1870), .Y(n1692) );
  OAI22X1 U2212 ( .A(n10061), .B(n9203), .C(n11671), .D(n1889), .Y(n8204) );
  OAI22X1 U2214 ( .A(n9248), .B(n10061), .C(n11670), .D(n1889), .Y(n8205) );
  OAI21X1 U2217 ( .A(n1891), .B(n1869), .C(n10244), .Y(n1889) );
  NOR2X1 U2219 ( .A(n1881), .B(n1870), .Y(n1700) );
  OAI22X1 U2220 ( .A(n10060), .B(n9204), .C(n11681), .D(n1893), .Y(n8206) );
  OAI22X1 U2222 ( .A(n9248), .B(n10060), .C(n11680), .D(n1893), .Y(n8207) );
  OAI21X1 U2225 ( .A(n1894), .B(n1869), .C(n10243), .Y(n1893) );
  NOR2X1 U2227 ( .A(n1886), .B(n1870), .Y(n1710) );
  OAI22X1 U2228 ( .A(n10120), .B(n9203), .C(n11709), .D(n1896), .Y(n8208) );
  OAI22X1 U2230 ( .A(n9248), .B(n10120), .C(n11708), .D(n1896), .Y(n8209) );
  OAI21X1 U2233 ( .A(n1871), .B(n1897), .C(n10242), .Y(n1896) );
  NOR2X1 U2235 ( .A(n1891), .B(n1870), .Y(n1712) );
  OAI22X1 U2236 ( .A(n10119), .B(n9205), .C(n11711), .D(n1899), .Y(n8210) );
  OAI22X1 U2238 ( .A(n9248), .B(n10119), .C(n11710), .D(n1899), .Y(n8211) );
  OAI21X1 U2241 ( .A(n1876), .B(n1897), .C(n10241), .Y(n1899) );
  NOR2X1 U2243 ( .A(n1894), .B(n1870), .Y(n1714) );
  NAND3X1 U2244 ( .A(n9291), .B(n9293), .C(n1902), .Y(n1870) );
  OAI22X1 U2245 ( .A(n10118), .B(n9203), .C(n11721), .D(n1904), .Y(n8212) );
  OAI22X1 U2247 ( .A(n9248), .B(n10118), .C(n11720), .D(n1904), .Y(n8213) );
  OAI21X1 U2250 ( .A(n1868), .B(n1897), .C(n10239), .Y(n1904) );
  NOR2X1 U2252 ( .A(n1724), .B(n1871), .Y(n1716) );
  OAI22X1 U2253 ( .A(n10117), .B(n9205), .C(n11731), .D(n1906), .Y(n8214) );
  OAI22X1 U2255 ( .A(n9248), .B(n10117), .C(n11730), .D(n1906), .Y(n8215) );
  OAI21X1 U2258 ( .A(n1725), .B(n1897), .C(n10238), .Y(n1906) );
  NOR2X1 U2260 ( .A(n1724), .B(n1876), .Y(n1718) );
  OAI22X1 U2261 ( .A(n10116), .B(n9204), .C(n11741), .D(n1908), .Y(n8216) );
  OAI22X1 U2263 ( .A(n9248), .B(n10116), .C(n11740), .D(n1908), .Y(n8217) );
  OAI21X1 U2266 ( .A(n1881), .B(n1897), .C(n10237), .Y(n1908) );
  NOR2X1 U2268 ( .A(n1724), .B(n1868), .Y(n1720) );
  OAI22X1 U2269 ( .A(n10281), .B(n11707), .C(n9248), .D(n1910), .Y(n8218) );
  OAI22X1 U2271 ( .A(n10281), .B(n11706), .C(n9204), .D(n1910), .Y(n8219) );
  NAND3X1 U2274 ( .A(n1911), .B(n9292), .C(n1912), .Y(n1910) );
  AOI21X1 U2275 ( .A(n1725), .B(n9205), .C(n1913), .Y(n1912) );
  NAND2X1 U2276 ( .A(n9509), .B(n9293), .Y(n1913) );
  AOI21X1 U2277 ( .A(n11557), .B(n1886), .C(n1914), .Y(n1911) );
  AOI22X1 U2279 ( .A(n1916), .B(n11557), .C(\U_1/U_1/U_1/opcode[12][1] ), .D(
        n10115), .Y(n1915) );
  AOI22X1 U2281 ( .A(n9180), .B(n1916), .C(\U_1/U_1/U_1/opcode[12][0] ), .D(
        n10115), .Y(n1918) );
  OAI21X1 U2283 ( .A(n1891), .B(n1897), .C(n10236), .Y(n1916) );
  NOR2X1 U2285 ( .A(n1724), .B(n1881), .Y(n1728) );
  AOI22X1 U2287 ( .A(n1920), .B(n11557), .C(\U_1/U_1/U_1/opcode[13][1] ), .D(
        n10112), .Y(n1919) );
  AOI22X1 U2289 ( .A(n9180), .B(n1920), .C(\U_1/U_1/U_1/opcode[13][0] ), .D(
        n10112), .Y(n1922) );
  OAI21X1 U2291 ( .A(n1894), .B(n1897), .C(n10227), .Y(n1920) );
  NOR2X1 U2293 ( .A(n1724), .B(n1886), .Y(n1738) );
  NAND3X1 U2294 ( .A(n9292), .B(n9293), .C(n1923), .Y(n1897) );
  AOI22X1 U2296 ( .A(n1925), .B(n11557), .C(\U_1/U_1/U_1/opcode[14][1] ), .D(
        n10109), .Y(n1924) );
  AOI22X1 U2298 ( .A(n9180), .B(n1925), .C(\U_1/U_1/U_1/opcode[14][0] ), .D(
        n10109), .Y(n1927) );
  OAI21X1 U2300 ( .A(n1871), .B(n1928), .C(n10218), .Y(n1925) );
  NOR2X1 U2302 ( .A(n1724), .B(n1891), .Y(n1748) );
  AOI22X1 U2304 ( .A(n1930), .B(n11557), .C(\U_1/U_1/U_1/opcode[15][1] ), .D(
        n10106), .Y(n1929) );
  AOI22X1 U2306 ( .A(n9180), .B(n1930), .C(\U_1/U_1/U_1/opcode[15][0] ), .D(
        n10106), .Y(n1932) );
  OAI21X1 U2308 ( .A(n1876), .B(n1928), .C(n10209), .Y(n1930) );
  NOR2X1 U2310 ( .A(n1724), .B(n1894), .Y(n1758) );
  NAND3X1 U2311 ( .A(n1902), .B(n9293), .C(n9292), .Y(n1724) );
  OAI22X1 U2312 ( .A(n10103), .B(n9205), .C(n11791), .D(n1934), .Y(n8228) );
  OAI22X1 U2314 ( .A(n9248), .B(n10103), .C(n11790), .D(n1934), .Y(n8229) );
  OAI21X1 U2317 ( .A(n1868), .B(n1928), .C(n10200), .Y(n1934) );
  NOR2X1 U2319 ( .A(n1935), .B(n1871), .Y(n1766) );
  OAI22X1 U2320 ( .A(n10102), .B(n9204), .C(n11801), .D(n1937), .Y(n8230) );
  OAI22X1 U2322 ( .A(n9248), .B(n10102), .C(n11800), .D(n1937), .Y(n8231) );
  OAI21X1 U2325 ( .A(n1725), .B(n1928), .C(n10199), .Y(n1937) );
  NOR2X1 U2327 ( .A(n1935), .B(n1876), .Y(n1768) );
  OAI22X1 U2328 ( .A(n10101), .B(n9203), .C(n11811), .D(n1939), .Y(n8232) );
  OAI22X1 U2330 ( .A(n9248), .B(n10101), .C(n11810), .D(n1939), .Y(n8233) );
  OAI21X1 U2333 ( .A(n1881), .B(n1928), .C(n10198), .Y(n1939) );
  NOR2X1 U2335 ( .A(n1935), .B(n1868), .Y(n1770) );
  OAI22X1 U2336 ( .A(n10100), .B(n9204), .C(n11821), .D(n1941), .Y(n8234) );
  OAI22X1 U2338 ( .A(n9248), .B(n10100), .C(n11820), .D(n1941), .Y(n8235) );
  OAI21X1 U2341 ( .A(n1886), .B(n1928), .C(n10197), .Y(n1941) );
  NOR2X1 U2343 ( .A(n1935), .B(n1725), .Y(n1772) );
  AOI22X1 U2345 ( .A(n1943), .B(n11557), .C(\U_1/U_1/U_1/opcode[20][1] ), .D(
        n10099), .Y(n1942) );
  AOI22X1 U2347 ( .A(n9180), .B(n1943), .C(\U_1/U_1/U_1/opcode[20][0] ), .D(
        n10099), .Y(n1945) );
  OAI21X1 U2349 ( .A(n1891), .B(n1928), .C(n10196), .Y(n1943) );
  NOR2X1 U2351 ( .A(n1935), .B(n1881), .Y(n1776) );
  AOI22X1 U2353 ( .A(n1947), .B(n11557), .C(\U_1/U_1/U_1/opcode[21][1] ), .D(
        n10096), .Y(n1946) );
  AOI22X1 U2355 ( .A(n9180), .B(n1947), .C(\U_1/U_1/U_1/opcode[21][0] ), .D(
        n10096), .Y(n1949) );
  OAI21X1 U2357 ( .A(n1894), .B(n1928), .C(n10187), .Y(n1947) );
  NOR2X1 U2359 ( .A(n1935), .B(n1886), .Y(n1786) );
  NAND3X1 U2360 ( .A(\U_1/U_1/U_1/writeptr[4] ), .B(n9291), .C(n1923), .Y(
        n1928) );
  AOI22X1 U2362 ( .A(n1951), .B(n11557), .C(\U_1/U_1/U_1/opcode[22][1] ), .D(
        n10093), .Y(n1950) );
  AOI22X1 U2364 ( .A(n9180), .B(n1951), .C(\U_1/U_1/U_1/opcode[22][0] ), .D(
        n10093), .Y(n1953) );
  OAI21X1 U2366 ( .A(n1871), .B(n1954), .C(n10178), .Y(n1951) );
  NOR2X1 U2368 ( .A(n1935), .B(n1891), .Y(n1796) );
  AOI22X1 U2370 ( .A(n1956), .B(n11557), .C(\U_1/U_1/U_1/opcode[23][1] ), .D(
        n10090), .Y(n1955) );
  AOI22X1 U2372 ( .A(n9180), .B(n1956), .C(\U_1/U_1/U_1/opcode[23][0] ), .D(
        n10090), .Y(n1958) );
  OAI21X1 U2374 ( .A(n1876), .B(n1954), .C(n10169), .Y(n1956) );
  NOR2X1 U2376 ( .A(n1935), .B(n1894), .Y(n1806) );
  NAND3X1 U2377 ( .A(n1902), .B(n9291), .C(n9294), .Y(n1935) );
  AOI22X1 U2379 ( .A(n1960), .B(n11557), .C(\U_1/U_1/U_1/opcode[24][1] ), .D(
        n10087), .Y(n1959) );
  AOI22X1 U2381 ( .A(n9180), .B(n1960), .C(\U_1/U_1/U_1/opcode[24][0] ), .D(
        n10087), .Y(n1962) );
  OAI21X1 U2383 ( .A(n1868), .B(n1954), .C(n10160), .Y(n1960) );
  NOR2X1 U2385 ( .A(n1963), .B(n1871), .Y(n1816) );
  AOI22X1 U2387 ( .A(n1965), .B(n11557), .C(\U_1/U_1/U_1/opcode[25][1] ), .D(
        n10084), .Y(n1964) );
  AOI22X1 U2389 ( .A(n9180), .B(n1965), .C(\U_1/U_1/U_1/opcode[25][0] ), .D(
        n10084), .Y(n1967) );
  OAI21X1 U2391 ( .A(n1725), .B(n1954), .C(n10151), .Y(n1965) );
  NOR2X1 U2393 ( .A(n1963), .B(n1876), .Y(n1826) );
  AOI22X1 U2395 ( .A(n1969), .B(n11557), .C(\U_1/U_1/U_1/opcode[26][1] ), .D(
        n10081), .Y(n1968) );
  AOI22X1 U2397 ( .A(n9180), .B(n1969), .C(\U_1/U_1/U_1/opcode[26][0] ), .D(
        n10081), .Y(n1971) );
  OAI21X1 U2399 ( .A(n1881), .B(n1954), .C(n10142), .Y(n1969) );
  NOR2X1 U2401 ( .A(n1963), .B(n1868), .Y(n1836) );
  NAND3X1 U2402 ( .A(n11669), .B(n9287), .C(n9290), .Y(n1868) );
  AOI22X1 U2404 ( .A(n1975), .B(n11557), .C(\U_1/U_1/U_1/opcode[27][1] ), .D(
        n10078), .Y(n1974) );
  AOI22X1 U2406 ( .A(n9180), .B(n1975), .C(\U_1/U_1/U_1/opcode[27][0] ), .D(
        n10078), .Y(n1977) );
  OAI21X1 U2408 ( .A(n1886), .B(n1954), .C(n10133), .Y(n1975) );
  NOR2X1 U2410 ( .A(n1963), .B(n1725), .Y(n1846) );
  NAND3X1 U2411 ( .A(\U_1/U_1/U_1/writeptr[0] ), .B(n9287), .C(n9290), .Y(
        n1725) );
  OAI22X1 U2412 ( .A(n10075), .B(n9203), .C(n11751), .D(n1979), .Y(n8252) );
  OAI22X1 U2414 ( .A(n9248), .B(n10075), .C(n11750), .D(n1979), .Y(n8253) );
  OAI21X1 U2417 ( .A(n1891), .B(n1954), .C(n10124), .Y(n1979) );
  NOR2X1 U2419 ( .A(n1963), .B(n1881), .Y(n1854) );
  NAND3X1 U2420 ( .A(n11669), .B(n9289), .C(\U_1/U_1/U_1/writeptr[2] ), .Y(
        n1881) );
  OAI22X1 U2421 ( .A(n10074), .B(n9205), .C(n11761), .D(n1982), .Y(n8254) );
  OAI22X1 U2423 ( .A(n9248), .B(n10074), .C(n11760), .D(n1982), .Y(n8255) );
  OAI21X1 U2426 ( .A(n1894), .B(n1954), .C(n10123), .Y(n1982) );
  NOR2X1 U2428 ( .A(n1963), .B(n1886), .Y(n1856) );
  NAND3X1 U2429 ( .A(\U_1/U_1/U_1/writeptr[0] ), .B(n9289), .C(n9288), .Y(
        n1886) );
  NAND3X1 U2430 ( .A(\U_1/U_1/U_1/writeptr[4] ), .B(n9292), .C(n1923), .Y(
        n1954) );
  OAI22X1 U2431 ( .A(n10059), .B(n9203), .C(n11771), .D(n1984), .Y(n8256) );
  OAI22X1 U2433 ( .A(n9248), .B(n10059), .C(n11770), .D(n1984), .Y(n8257) );
  OAI21X1 U2436 ( .A(n1871), .B(n1869), .C(n10122), .Y(n1984) );
  NOR2X1 U2438 ( .A(n1963), .B(n1891), .Y(n1858) );
  NAND3X1 U2439 ( .A(n9290), .B(n11669), .C(\U_1/U_1/U_1/writeptr[2] ), .Y(
        n1891) );
  NAND3X1 U2440 ( .A(n9289), .B(n9287), .C(n11669), .Y(n1871) );
  OAI22X1 U2441 ( .A(n10058), .B(n9205), .C(n11781), .D(n1986), .Y(n8258) );
  OAI22X1 U2443 ( .A(n9248), .B(n10058), .C(n11780), .D(n1986), .Y(n8259) );
  OAI21X1 U2446 ( .A(n1876), .B(n1869), .C(n10121), .Y(n1986) );
  NOR2X1 U2448 ( .A(n1963), .B(n1894), .Y(n1860) );
  NAND3X1 U2449 ( .A(n9290), .B(\U_1/U_1/U_1/writeptr[0] ), .C(
        \U_1/U_1/U_1/writeptr[2] ), .Y(n1894) );
  NAND3X1 U2450 ( .A(n9292), .B(n1902), .C(n9294), .Y(n1963) );
  NAND3X1 U2452 ( .A(n9291), .B(n9293), .C(n1923), .Y(n1869) );
  NAND3X1 U2454 ( .A(n9289), .B(n9287), .C(\U_1/U_1/U_1/writeptr[0] ), .Y(
        n1876) );
  OAI21X1 U2455 ( .A(n11545), .B(n9291), .C(n1990), .Y(n8260) );
  AOI22X1 U2456 ( .A(\U_1/U_1/U_1/N50 ), .B(n1987), .C(\U_1/U_1/U_1/N45 ), .D(
        n1988), .Y(n1990) );
  OAI21X1 U2458 ( .A(n11545), .B(n9287), .C(n1991), .Y(n8261) );
  AOI22X1 U2459 ( .A(\U_1/U_1/U_1/N49 ), .B(n1987), .C(\U_1/U_1/U_1/N44 ), .D(
        n1988), .Y(n1991) );
  OAI21X1 U2461 ( .A(n11545), .B(n9289), .C(n1992), .Y(n8262) );
  AOI22X1 U2462 ( .A(\U_1/U_1/U_1/N48 ), .B(n1987), .C(\U_1/U_1/U_1/N43 ), .D(
        n1988), .Y(n1992) );
  OAI21X1 U2464 ( .A(n11545), .B(n11669), .C(n1993), .Y(n8263) );
  AOI22X1 U2465 ( .A(n11669), .B(n1987), .C(n11669), .D(n1988), .Y(n1993) );
  OAI21X1 U2467 ( .A(n11545), .B(n9293), .C(n1994), .Y(n8264) );
  AOI22X1 U2468 ( .A(\U_1/U_1/U_1/N51 ), .B(n1987), .C(\U_1/U_1/U_1/N46 ), .D(
        n1988), .Y(n1994) );
  NOR2X1 U2469 ( .A(n1914), .B(n9204), .Y(n1988) );
  NOR2X1 U2470 ( .A(n1914), .B(n11557), .Y(n1987) );
  NAND2X1 U2473 ( .A(\U_1/U_1/U_1/N36 ), .B(n9453), .Y(n1914) );
  OAI21X1 U2474 ( .A(n11866), .B(n879), .C(n1996), .Y(n8265) );
  AOI22X1 U2475 ( .A(\U_1/U_3/U_3/N84 ), .B(n881), .C(\U_1/U_3/U_3/N59 ), .D(
        n882), .Y(n1996) );
  OAI21X1 U2477 ( .A(n11653), .B(n1999), .C(n2000), .Y(n1997) );
  NOR2X1 U2478 ( .A(n11648), .B(n11643), .Y(n2000) );
  NAND2X1 U2479 ( .A(n11646), .B(n11656), .Y(n1999) );
  OAI21X1 U2480 ( .A(n2004), .B(n237), .C(n2005), .Y(n881) );
  OAI21X1 U2481 ( .A(n11646), .B(n11845), .C(n11654), .Y(n2005) );
  NAND2X1 U2482 ( .A(n11648), .B(n11623), .Y(n879) );
  OAI21X1 U2483 ( .A(RST), .B(n9719), .C(n2010), .Y(n8266) );
  NAND2X1 U2484 ( .A(CRCE_S), .B(RST), .Y(n2010) );
  OAI22X1 U2485 ( .A(n9531), .B(n11619), .C(RST), .D(n9719), .Y(n8267) );
  OAI21X1 U2487 ( .A(n9720), .B(n11619), .C(n2014), .Y(n2012) );
  NAND3X1 U2488 ( .A(n11557), .B(n11570), .C(n2016), .Y(n2014) );
  OAI21X1 U2490 ( .A(n9452), .B(n11571), .C(n2019), .Y(n8268) );
  NAND2X1 U2491 ( .A(\U_1/U_2/rx_CHECK_CRC [15]), .B(n9452), .Y(n2019) );
  OAI21X1 U2492 ( .A(n9452), .B(n11615), .C(n2021), .Y(n8269) );
  NAND2X1 U2493 ( .A(\U_1/U_2/rx_CHECK_CRC [14]), .B(n9452), .Y(n2021) );
  OAI21X1 U2494 ( .A(n9452), .B(n11614), .C(n2023), .Y(n8270) );
  NAND2X1 U2495 ( .A(\U_1/U_2/rx_CHECK_CRC [13]), .B(n9452), .Y(n2023) );
  OAI21X1 U2496 ( .A(n9452), .B(n11613), .C(n2025), .Y(n8271) );
  NAND2X1 U2497 ( .A(\U_1/U_2/rx_CHECK_CRC [12]), .B(n9452), .Y(n2025) );
  OAI21X1 U2498 ( .A(n9452), .B(n11612), .C(n2027), .Y(n8272) );
  NAND2X1 U2499 ( .A(\U_1/U_2/rx_CHECK_CRC [11]), .B(n9452), .Y(n2027) );
  OAI21X1 U2500 ( .A(n9452), .B(n11611), .C(n2029), .Y(n8273) );
  NAND2X1 U2501 ( .A(\U_1/U_2/rx_CHECK_CRC [10]), .B(n9452), .Y(n2029) );
  OAI21X1 U2502 ( .A(n9452), .B(n9636), .C(n2031), .Y(n8274) );
  NAND2X1 U2503 ( .A(\U_1/U_2/rx_CHECK_CRC [9]), .B(n9452), .Y(n2031) );
  OAI21X1 U2504 ( .A(n9452), .B(n11610), .C(n2033), .Y(n8275) );
  NAND2X1 U2505 ( .A(\U_1/U_2/rx_CHECK_CRC [8]), .B(n9452), .Y(n2033) );
  OAI22X1 U2506 ( .A(n11571), .B(n9453), .C(n9452), .D(n9316), .Y(n8276) );
  OAI22X1 U2508 ( .A(n9454), .B(n11615), .C(n9452), .D(n9314), .Y(n8277) );
  OAI22X1 U2510 ( .A(n9453), .B(n11614), .C(n9452), .D(n9312), .Y(n8278) );
  OAI22X1 U2512 ( .A(n9454), .B(n11613), .C(n9452), .D(n9310), .Y(n8279) );
  OAI22X1 U2514 ( .A(n9454), .B(n11612), .C(n9452), .D(n9308), .Y(n8280) );
  OAI22X1 U2516 ( .A(n9455), .B(n11611), .C(n9452), .D(n9306), .Y(n8281) );
  OAI22X1 U2518 ( .A(n9455), .B(n9636), .C(n9452), .D(n9304), .Y(n8282) );
  OAI22X1 U2520 ( .A(n9453), .B(n11610), .C(n9452), .D(n9302), .Y(n8283) );
  OAI21X1 U2524 ( .A(n9376), .B(n11598), .C(n2037), .Y(n8284) );
  NAND2X1 U2525 ( .A(\U_1/U_2/RX_CRC [14]), .B(n9378), .Y(n2037) );
  OAI22X1 U2526 ( .A(n9375), .B(n11597), .C(n9251), .D(n11598), .Y(n8285) );
  OAI22X1 U2528 ( .A(n9249), .B(n11595), .C(n11597), .D(n9250), .Y(n8286) );
  OAI21X1 U2529 ( .A(n9376), .B(n11601), .C(n2044), .Y(n8287) );
  NAND2X1 U2530 ( .A(\U_1/U_2/RX_CRC [13]), .B(n9378), .Y(n2044) );
  OAI22X1 U2531 ( .A(n9375), .B(n11594), .C(n9251), .D(n11601), .Y(n8288) );
  OAI22X1 U2533 ( .A(n9249), .B(n11592), .C(n9250), .D(n11594), .Y(n8289) );
  OAI21X1 U2535 ( .A(n9376), .B(n11591), .C(n2048), .Y(n8290) );
  NAND2X1 U2536 ( .A(\U_1/U_2/RX_CRC [12]), .B(n9378), .Y(n2048) );
  OAI22X1 U2537 ( .A(n9375), .B(n11590), .C(n9251), .D(n11591), .Y(n8291) );
  OAI22X1 U2539 ( .A(n9249), .B(n11588), .C(n9250), .D(n11590), .Y(n8292) );
  OAI21X1 U2541 ( .A(n9376), .B(n11602), .C(n2052), .Y(n8293) );
  NAND2X1 U2542 ( .A(\U_1/U_2/RX_CRC [11]), .B(n9377), .Y(n2052) );
  OAI22X1 U2543 ( .A(n9375), .B(n11587), .C(n9251), .D(n11602), .Y(n8294) );
  OAI22X1 U2545 ( .A(n9249), .B(n11585), .C(n9250), .D(n11587), .Y(n8295) );
  OAI21X1 U2547 ( .A(n9376), .B(n11607), .C(n2056), .Y(n8296) );
  NAND2X1 U2548 ( .A(\U_1/U_2/RX_CRC [10]), .B(n9377), .Y(n2056) );
  OAI22X1 U2549 ( .A(n9375), .B(n11584), .C(n9251), .D(n11607), .Y(n8297) );
  OAI22X1 U2551 ( .A(n9249), .B(n11582), .C(n9250), .D(n11584), .Y(n8298) );
  OAI21X1 U2553 ( .A(n9376), .B(n11606), .C(n2060), .Y(n8299) );
  NAND2X1 U2554 ( .A(\U_1/U_2/RX_CRC [9]), .B(n9377), .Y(n2060) );
  OAI22X1 U2555 ( .A(n9376), .B(n11605), .C(n9251), .D(n11606), .Y(n8300) );
  OAI22X1 U2557 ( .A(n9250), .B(n11605), .C(n2062), .D(n9249), .Y(n8301) );
  XNOR2X1 U2558 ( .A(\U_1/U_2/U_2/current_crc[1] ), .B(n2063), .Y(n2062) );
  OAI21X1 U2560 ( .A(n9376), .B(n11608), .C(n2065), .Y(n8302) );
  NAND2X1 U2561 ( .A(\U_1/U_2/RX_CRC [8]), .B(n9377), .Y(n2065) );
  OAI22X1 U2562 ( .A(n9376), .B(n11581), .C(n9251), .D(n11608), .Y(n8303) );
  OAI22X1 U2564 ( .A(n9250), .B(n11581), .C(n2067), .D(n9249), .Y(n8304) );
  XOR2X1 U2565 ( .A(n2068), .B(n2069), .Y(n2067) );
  XNOR2X1 U2566 ( .A(\U_1/U_2/U_2/current_crc[0] ), .B(n2063), .Y(n2068) );
  OAI21X1 U2568 ( .A(n9376), .B(n11600), .C(n2071), .Y(n8305) );
  NAND2X1 U2569 ( .A(\U_1/U_2/RX_CRC [7]), .B(n9377), .Y(n2071) );
  OAI22X1 U2570 ( .A(n9375), .B(n11599), .C(n9251), .D(n11600), .Y(n8306) );
  OAI22X1 U2572 ( .A(n9250), .B(n11599), .C(n2073), .D(n9249), .Y(n8307) );
  OAI21X1 U2573 ( .A(n9376), .B(n11596), .C(n2075), .Y(n8308) );
  NAND2X1 U2574 ( .A(\U_1/U_2/RX_CRC [6]), .B(n9377), .Y(n2075) );
  OAI22X1 U2575 ( .A(n9376), .B(n11595), .C(n9251), .D(n11596), .Y(n8309) );
  OAI22X1 U2577 ( .A(n9250), .B(n11595), .C(n2076), .D(n9249), .Y(n8310) );
  XNOR2X1 U2578 ( .A(n2077), .B(n2078), .Y(n2076) );
  OAI21X1 U2580 ( .A(n9377), .B(n11593), .C(n2080), .Y(n8311) );
  NAND2X1 U2581 ( .A(\U_1/U_2/RX_CRC [5]), .B(n9377), .Y(n2080) );
  OAI22X1 U2582 ( .A(n9375), .B(n11592), .C(n9251), .D(n11593), .Y(n8312) );
  OAI22X1 U2584 ( .A(n9250), .B(n11592), .C(n2081), .D(n9249), .Y(n8313) );
  OAI21X1 U2586 ( .A(n9377), .B(n11589), .C(n2083), .Y(n8314) );
  NAND2X1 U2587 ( .A(\U_1/U_2/RX_CRC [4]), .B(n9377), .Y(n2083) );
  OAI22X1 U2588 ( .A(n9376), .B(n11588), .C(n9251), .D(n11589), .Y(n8315) );
  OAI22X1 U2590 ( .A(n9250), .B(n11588), .C(n2084), .D(n9249), .Y(n8316) );
  XNOR2X1 U2591 ( .A(n2085), .B(n2086), .Y(n2084) );
  OAI21X1 U2593 ( .A(n9377), .B(n11586), .C(n2088), .Y(n8317) );
  NAND2X1 U2594 ( .A(\U_1/U_2/RX_CRC [3]), .B(n9378), .Y(n2088) );
  OAI22X1 U2595 ( .A(n9375), .B(n11585), .C(n9251), .D(n11586), .Y(n8318) );
  OAI22X1 U2597 ( .A(n9250), .B(n11585), .C(n2089), .D(n9249), .Y(n8319) );
  OAI21X1 U2599 ( .A(n9377), .B(n11583), .C(n2091), .Y(n8320) );
  NAND2X1 U2600 ( .A(\U_1/U_2/RX_CRC [2]), .B(n9378), .Y(n2091) );
  OAI22X1 U2601 ( .A(n9375), .B(n11582), .C(n9251), .D(n11583), .Y(n8321) );
  OAI22X1 U2603 ( .A(n9250), .B(n11582), .C(n2092), .D(n9249), .Y(n8322) );
  XNOR2X1 U2604 ( .A(n2093), .B(n2094), .Y(n2092) );
  OAI21X1 U2606 ( .A(n9377), .B(n11604), .C(n2096), .Y(n8323) );
  NAND2X1 U2607 ( .A(\U_1/U_2/RX_CRC [1]), .B(n9378), .Y(n2096) );
  OAI22X1 U2608 ( .A(n9375), .B(n11603), .C(n9251), .D(n11604), .Y(n8324) );
  OAI22X1 U2610 ( .A(n9250), .B(n11603), .C(n2098), .D(n9249), .Y(n8325) );
  XOR2X1 U2611 ( .A(n2099), .B(n2100), .Y(n2098) );
  OAI21X1 U2613 ( .A(n9377), .B(n11580), .C(n2102), .Y(n8326) );
  NAND2X1 U2614 ( .A(\U_1/U_2/RX_CRC [0]), .B(n9378), .Y(n2102) );
  OAI22X1 U2615 ( .A(n9375), .B(n11579), .C(n9251), .D(n11580), .Y(n8327) );
  OAI22X1 U2617 ( .A(n9250), .B(n11579), .C(n2104), .D(n9249), .Y(n8328) );
  OAI22X1 U2619 ( .A(n9532), .B(n11618), .C(RST), .D(n761), .Y(n8329) );
  NOR2X1 U2620 ( .A(n2106), .B(n2107), .Y(n761) );
  OAI21X1 U2621 ( .A(n2108), .B(n9698), .C(n2109), .Y(n2107) );
  OAI21X1 U2622 ( .A(n9720), .B(n11618), .C(n2110), .Y(n2106) );
  OAI21X1 U2624 ( .A(n2112), .B(n2113), .C(n2114), .Y(n2111) );
  NAND2X1 U2625 ( .A(n2115), .B(n11577), .Y(n2113) );
  OAI21X1 U2627 ( .A(n9701), .B(n11573), .C(n2119), .Y(n8330) );
  NAND3X1 U2628 ( .A(n9247), .B(n11573), .C(n9700), .Y(n2119) );
  OAI21X1 U2630 ( .A(n2123), .B(n11574), .C(n2125), .Y(n8331) );
  NAND3X1 U2631 ( .A(n9247), .B(n11574), .C(n2126), .Y(n2125) );
  NOR2X1 U2632 ( .A(n2127), .B(n11573), .Y(n2126) );
  AOI21X1 U2633 ( .A(n2128), .B(n11573), .C(n2122), .Y(n2123) );
  OAI21X1 U2634 ( .A(n9247), .B(n11548), .C(n2130), .Y(n2122) );
  OAI21X1 U2635 ( .A(n9699), .B(n11575), .C(n2133), .Y(n8332) );
  NAND3X1 U2636 ( .A(n9700), .B(n11575), .C(n9717), .Y(n2133) );
  OAI21X1 U2638 ( .A(n2136), .B(n11576), .C(n2138), .Y(n8333) );
  NAND3X1 U2639 ( .A(n9700), .B(n11576), .C(n2139), .Y(n2138) );
  NOR2X1 U2640 ( .A(n2140), .B(n11575), .Y(n2139) );
  NAND2X1 U2642 ( .A(n2128), .B(n2130), .Y(n2127) );
  AOI21X1 U2643 ( .A(n2128), .B(n11575), .C(n2135), .Y(n2136) );
  OAI21X1 U2644 ( .A(n9717), .B(n11548), .C(n2130), .Y(n2135) );
  NAND3X1 U2647 ( .A(\U_1/U_2/U_5/count[0] ), .B(n9247), .C(
        \U_1/U_2/U_5/count[1] ), .Y(n2140) );
  NOR2X1 U2648 ( .A(n11549), .B(n2142), .Y(n2128) );
  OAI21X1 U2649 ( .A(n9377), .B(n11609), .C(n2144), .Y(n8334) );
  NAND2X1 U2650 ( .A(\U_1/U_2/RX_CRC [15]), .B(n9378), .Y(n2144) );
  OAI22X1 U2651 ( .A(n9375), .B(n11578), .C(n9251), .D(n11609), .Y(n8335) );
  OAI22X1 U2655 ( .A(n9250), .B(n11578), .C(n2146), .D(n9249), .Y(n8336) );
  XNOR2X1 U2656 ( .A(n2104), .B(n11599), .Y(n2146) );
  XOR2X1 U2658 ( .A(n2147), .B(n2100), .Y(n2104) );
  XOR2X1 U2659 ( .A(n2089), .B(n2081), .Y(n2100) );
  XNOR2X1 U2660 ( .A(n2086), .B(n2077), .Y(n2081) );
  XNOR2X1 U2661 ( .A(\U_1/U_2/U_2/current_crc[12] ), .B(n9310), .Y(n2077) );
  XNOR2X1 U2662 ( .A(\U_1/U_2/U_2/current_crc[11] ), .B(n9308), .Y(n2086) );
  XNOR2X1 U2663 ( .A(n2094), .B(n2085), .Y(n2089) );
  XNOR2X1 U2664 ( .A(\U_1/U_2/U_2/current_crc[10] ), .B(n9306), .Y(n2085) );
  XNOR2X1 U2665 ( .A(\U_1/U_2/U_2/current_crc[9] ), .B(n9304), .Y(n2094) );
  XOR2X1 U2666 ( .A(n2099), .B(n2093), .Y(n2147) );
  XNOR2X1 U2667 ( .A(\U_1/U_2/U_2/current_crc[8] ), .B(n9302), .Y(n2093) );
  XOR2X1 U2668 ( .A(n2063), .B(n2073), .Y(n2099) );
  XNOR2X1 U2669 ( .A(n2078), .B(n2069), .Y(n2073) );
  XNOR2X1 U2670 ( .A(n11597), .B(n9315), .Y(n2069) );
  XNOR2X1 U2672 ( .A(\U_1/U_2/U_2/current_crc[13] ), .B(n9312), .Y(n2078) );
  XNOR2X1 U2673 ( .A(\U_1/U_2/U_2/current_crc[15] ), .B(n9316), .Y(n2063) );
  OAI22X1 U2679 ( .A(n9247), .B(n9302), .C(n9304), .D(n9182), .Y(n8337) );
  OAI22X1 U2680 ( .A(n9247), .B(n9304), .C(n9306), .D(n9182), .Y(n8338) );
  OAI22X1 U2682 ( .A(n9247), .B(n9306), .C(n9308), .D(n9182), .Y(n8339) );
  OAI22X1 U2684 ( .A(n9247), .B(n9308), .C(n9310), .D(n9182), .Y(n8340) );
  OAI22X1 U2685 ( .A(n9247), .B(n9310), .C(n9312), .D(n9182), .Y(n8341) );
  OAI22X1 U2686 ( .A(n9247), .B(n9312), .C(n9314), .D(n9182), .Y(n8342) );
  OAI22X1 U2688 ( .A(n9247), .B(n9314), .C(n9316), .D(n9182), .Y(n8343) );
  OAI22X1 U2690 ( .A(n9247), .B(n9316), .C(n9182), .D(n2150), .Y(n8344) );
  XNOR2X1 U2691 ( .A(n11566), .B(\U_1/U_2/U_1/DP_hold1 ), .Y(n2150) );
  NAND2X1 U2694 ( .A(n2152), .B(n2153), .Y(n8345) );
  AOI22X1 U2695 ( .A(DPRS), .B(n11563), .C(\U_1/U_2/U_1/DP_hold1 ), .D(n2155), 
        .Y(n2152) );
  OAI21X1 U2696 ( .A(n11566), .B(n2156), .C(n2157), .Y(n8346) );
  OAI21X1 U2697 ( .A(\U_1/U_2/U_1/DP_hold1 ), .B(n9702), .C(n2156), .Y(n2157)
         );
  NOR2X1 U2699 ( .A(\U_1/U_2/U_1/state[3] ), .B(n9202), .Y(n2153) );
  OAI21X1 U2700 ( .A(n2155), .B(n11563), .C(n2160), .Y(n2156) );
  NOR2X1 U2701 ( .A(n9202), .B(n9247), .Y(n2160) );
  NOR3X1 U2704 ( .A(n2163), .B(n2164), .C(n2165), .Y(n2162) );
  OAI21X1 U2705 ( .A(n9442), .B(n11542), .C(n2167), .Y(n8347) );
  AOI22X1 U2706 ( .A(n2168), .B(n2169), .C(n9447), .D(n11397), .Y(n2167) );
  OAI22X1 U2707 ( .A(n2172), .B(n2173), .C(n9246), .D(n2175), .Y(n2168) );
  OAI21X1 U2708 ( .A(\U_1/U_0/U_1/RCV_DATA [5]), .B(n2176), .C(n9446), .Y(
        n2173) );
  OAI21X1 U2709 ( .A(n11379), .B(n2179), .C(n9246), .Y(n2172) );
  AOI22X1 U2710 ( .A(n2180), .B(n2181), .C(n11501), .D(n11518), .Y(n2179) );
  OAI22X1 U2711 ( .A(\U_1/U_0/U_1/RCV_DATA [3]), .B(n2183), .C(n11432), .D(
        n2185), .Y(n2180) );
  AOI22X1 U2712 ( .A(n2186), .B(n2187), .C(n11483), .D(n9475), .Y(n2185) );
  OAI22X1 U2714 ( .A(n2189), .B(n11415), .C(\U_1/U_0/U_1/RCV_DATA [1]), .D(
        n2191), .Y(n2186) );
  NAND2X1 U2716 ( .A(n2192), .B(n2193), .Y(n2191) );
  AOI22X1 U2717 ( .A(n2194), .B(n9480), .C(n11466), .D(n11542), .Y(n2189) );
  NOR2X1 U2720 ( .A(n2196), .B(n2197), .Y(n2194) );
  NAND2X1 U2722 ( .A(n10057), .B(n2199), .Y(n8348) );
  AOI22X1 U2723 ( .A(n9443), .B(\U_1/U_0/U_1/U_8/currentPlainKey[62] ), .C(
        n9447), .D(n11450), .Y(n2199) );
  OAI22X1 U2725 ( .A(n2175), .B(n2169), .C(n2203), .D(n2204), .Y(n2202) );
  OAI21X1 U2726 ( .A(n2205), .B(n2206), .C(n9446), .Y(n2204) );
  OAI22X1 U2727 ( .A(n11516), .B(n9246), .C(n11518), .D(n2176), .Y(n2206) );
  OAI21X1 U2728 ( .A(n9393), .B(n2181), .C(n2207), .Y(n2205) );
  AOI22X1 U2729 ( .A(n11432), .B(n9474), .C(n11380), .D(n2209), .Y(n2207) );
  OAI21X1 U2730 ( .A(n9402), .B(n2187), .C(n2210), .Y(n2209) );
  NAND2X1 U2731 ( .A(n2211), .B(n2187), .Y(n2210) );
  OAI21X1 U2732 ( .A(n2212), .B(n2213), .C(n2214), .Y(n2211) );
  OAI21X1 U2733 ( .A(n2212), .B(n2196), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[62] ), .Y(n2214) );
  NAND2X1 U2734 ( .A(n2215), .B(n2193), .Y(n2187) );
  NAND2X1 U2736 ( .A(n2217), .B(n2169), .Y(n2203) );
  NAND2X1 U2737 ( .A(n2218), .B(n2219), .Y(n8349) );
  AOI22X1 U2738 ( .A(n2220), .B(n2221), .C(n11450), .D(n9370), .Y(n2219) );
  OAI21X1 U2739 ( .A(n11516), .B(n2169), .C(n2223), .Y(n2221) );
  OAI21X1 U2740 ( .A(n2224), .B(n2225), .C(n2169), .Y(n2223) );
  OAI22X1 U2741 ( .A(n11518), .B(n9246), .C(n9475), .D(n2181), .Y(n2225) );
  OAI21X1 U2742 ( .A(n2226), .B(n2216), .C(n2227), .Y(n2224) );
  AOI22X1 U2743 ( .A(n11432), .B(\U_1/U_0/U_1/RCV_DATA [1]), .C(n11379), .D(
        \U_1/U_0/U_1/RCV_DATA [3]), .Y(n2227) );
  NAND2X1 U2746 ( .A(n2228), .B(n2183), .Y(n2216) );
  NAND2X1 U2747 ( .A(n2229), .B(n2193), .Y(n2183) );
  AOI22X1 U2748 ( .A(n2230), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[61] ), .D(n11484), .Y(n2226) );
  NOR2X1 U2750 ( .A(n2196), .B(n2232), .Y(n2230) );
  AOI22X1 U2751 ( .A(n11399), .B(n9447), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[61] ), .D(n9441), .Y(n2218) );
  NAND2X1 U2752 ( .A(n2234), .B(n2235), .Y(n8350) );
  AOI22X1 U2753 ( .A(n2236), .B(n2237), .C(n11399), .D(n9370), .Y(n2235) );
  OAI21X1 U2754 ( .A(n10054), .B(n2239), .C(n2240), .Y(n2236) );
  AOI22X1 U2755 ( .A(n9440), .B(n11397), .C(n2242), .D(n11450), .Y(n2240) );
  OAI21X1 U2756 ( .A(n2243), .B(n2244), .C(n2169), .Y(n2239) );
  OAI22X1 U2757 ( .A(n9393), .B(n9246), .C(n9476), .D(n2176), .Y(n2244) );
  OAI21X1 U2758 ( .A(n9402), .B(n2181), .C(n2245), .Y(n2243) );
  NAND2X1 U2759 ( .A(n2228), .B(n2246), .Y(n2245) );
  OAI21X1 U2760 ( .A(n2247), .B(n2213), .C(n2248), .Y(n2246) );
  OAI21X1 U2761 ( .A(n2247), .B(n2196), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[60] ), .Y(n2248) );
  NOR2X1 U2762 ( .A(n2249), .B(n11501), .Y(n2228) );
  NAND2X1 U2764 ( .A(n2250), .B(n2193), .Y(n2181) );
  AOI22X1 U2766 ( .A(n11467), .B(n9447), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[60] ), .D(n9441), .Y(n2234) );
  NAND2X1 U2767 ( .A(n2252), .B(n2253), .Y(n8351) );
  AOI22X1 U2768 ( .A(n2254), .B(n2255), .C(n11467), .D(n9370), .Y(n2253) );
  OAI21X1 U2769 ( .A(n2256), .B(n9365), .C(n2258), .Y(n2255) );
  AOI22X1 U2770 ( .A(n2220), .B(n2259), .C(n9439), .D(n11450), .Y(n2258) );
  OAI21X1 U2771 ( .A(n9393), .B(n2169), .C(n2260), .Y(n2259) );
  OAI21X1 U2772 ( .A(n2261), .B(n2262), .C(n2169), .Y(n2260) );
  OAI22X1 U2773 ( .A(n9398), .B(n2176), .C(n2263), .D(n2249), .Y(n2262) );
  NAND2X1 U2774 ( .A(n2176), .B(n9246), .Y(n2249) );
  AOI22X1 U2775 ( .A(n2264), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[59] ), .D(n11502), .Y(n2263) );
  NOR2X1 U2777 ( .A(n2196), .B(n2266), .Y(n2264) );
  NAND2X1 U2778 ( .A(n2267), .B(n2193), .Y(n2176) );
  NOR2X1 U2779 ( .A(n9477), .B(n9246), .Y(n2261) );
  NOR2X1 U2780 ( .A(n11398), .B(n9444), .Y(n2220) );
  AOI22X1 U2781 ( .A(n11416), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[59] ), .D(n9441), .Y(n2252) );
  NAND2X1 U2782 ( .A(n2271), .B(n2272), .Y(n8352) );
  AOI22X1 U2783 ( .A(n2273), .B(n2274), .C(n11416), .D(n9370), .Y(n2272) );
  OAI21X1 U2784 ( .A(n9365), .B(n2237), .C(n2275), .Y(n2274) );
  AOI22X1 U2785 ( .A(n2276), .B(n2277), .C(n9438), .D(n11399), .Y(n2275) );
  NOR2X1 U2786 ( .A(n11399), .B(n11467), .Y(n2277) );
  NOR2X1 U2787 ( .A(n2278), .B(n9444), .Y(n2276) );
  AOI21X1 U2788 ( .A(n11450), .B(\U_1/U_0/U_1/RCV_DATA [3]), .C(n2279), .Y(
        n2278) );
  OAI21X1 U2789 ( .A(n9477), .B(n2169), .C(n2280), .Y(n2279) );
  NAND3X1 U2790 ( .A(n2217), .B(n2169), .C(n2281), .Y(n2280) );
  OAI22X1 U2791 ( .A(n9398), .B(n9246), .C(n9170), .D(n2283), .Y(n2281) );
  AOI22X1 U2792 ( .A(n2284), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[58] ), .D(n11381), .Y(n2283) );
  NOR2X1 U2794 ( .A(n2196), .B(n2286), .Y(n2284) );
  AOI22X1 U2797 ( .A(n11485), .B(n9447), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[58] ), .D(n9441), .Y(n2271) );
  NAND2X1 U2798 ( .A(n2289), .B(n2290), .Y(n8353) );
  AOI22X1 U2799 ( .A(n2291), .B(n2292), .C(n11485), .D(n9370), .Y(n2290) );
  OAI21X1 U2800 ( .A(n9365), .B(n2293), .C(n2294), .Y(n2292) );
  AOI22X1 U2801 ( .A(n2295), .B(n2254), .C(n11467), .D(n9440), .Y(n2294) );
  NOR2X1 U2802 ( .A(n2296), .B(n9444), .Y(n2295) );
  AOI21X1 U2803 ( .A(n11399), .B(\U_1/U_0/U_1/RCV_DATA [3]), .C(n2297), .Y(
        n2296) );
  OAI22X1 U2804 ( .A(n9476), .B(n2217), .C(n2298), .D(n11398), .Y(n2297) );
  AOI22X1 U2806 ( .A(n2300), .B(n2169), .C(n11397), .D(
        \U_1/U_0/U_1/RCV_DATA [1]), .Y(n2298) );
  NAND2X1 U2808 ( .A(n2193), .B(n2301), .Y(n2169) );
  OAI21X1 U2809 ( .A(n2302), .B(n2213), .C(n2303), .Y(n2300) );
  OAI21X1 U2810 ( .A(n2302), .B(n2196), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[57] ), .Y(n2303) );
  AOI22X1 U2811 ( .A(n11363), .B(n9447), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[57] ), .D(n9441), .Y(n2289) );
  NAND2X1 U2812 ( .A(n2305), .B(n2306), .Y(n8354) );
  AOI22X1 U2813 ( .A(n2307), .B(n2308), .C(n11363), .D(n9370), .Y(n2306) );
  OAI21X1 U2814 ( .A(n9365), .B(n2309), .C(n2310), .Y(n2308) );
  AOI22X1 U2815 ( .A(n2311), .B(n2273), .C(n11416), .D(n9439), .Y(n2310) );
  NOR2X1 U2816 ( .A(n2312), .B(n9444), .Y(n2311) );
  AOI21X1 U2817 ( .A(n11467), .B(\U_1/U_0/U_1/RCV_DATA [3]), .C(n2313), .Y(
        n2312) );
  OAI22X1 U2818 ( .A(n9476), .B(n2256), .C(n11467), .D(n2314), .Y(n2313) );
  AOI22X1 U2819 ( .A(n11450), .B(\U_1/U_0/U_1/RCV_DATA [1]), .C(n2299), .D(
        n2315), .Y(n2314) );
  OAI21X1 U2820 ( .A(n2316), .B(n2213), .C(n2317), .Y(n2315) );
  OAI21X1 U2821 ( .A(n2316), .B(n2196), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[56] ), .Y(n2317) );
  NAND2X1 U2822 ( .A(n11509), .B(n9479), .Y(n2213) );
  NAND2X1 U2824 ( .A(\U_1/U_0/U_1/U_8/address[3] ), .B(n2319), .Y(n2196) );
  NOR2X1 U2825 ( .A(n11399), .B(n11450), .Y(n2299) );
  NAND2X1 U2827 ( .A(n2320), .B(n11461), .Y(n2217) );
  AOI22X1 U2829 ( .A(n11434), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[56] ), .D(n2200), .Y(n2305) );
  NAND2X1 U2830 ( .A(n2323), .B(n2324), .Y(n8355) );
  AOI22X1 U2831 ( .A(n2325), .B(n2326), .C(n11434), .D(n9370), .Y(n2324) );
  OAI21X1 U2832 ( .A(n9365), .B(n2327), .C(n2328), .Y(n2326) );
  AOI22X1 U2833 ( .A(n2329), .B(n2291), .C(n11485), .D(n9440), .Y(n2328) );
  OAI21X1 U2835 ( .A(n9393), .B(n2293), .C(n2331), .Y(n2330) );
  AOI22X1 U2836 ( .A(n2254), .B(n2332), .C(n11467), .D(n9474), .Y(n2331) );
  OAI22X1 U2837 ( .A(n9398), .B(n2256), .C(n11399), .D(n2333), .Y(n2332) );
  AOI22X1 U2838 ( .A(n11451), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[55] ), .D(n2335), .Y(n2333) );
  NAND2X1 U2840 ( .A(n2336), .B(n11461), .Y(n2335) );
  NAND2X1 U2842 ( .A(n2320), .B(n11410), .Y(n2256) );
  NOR2X1 U2843 ( .A(n11416), .B(n11467), .Y(n2254) );
  AOI22X1 U2844 ( .A(n11382), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[55] ), .D(n9443), .Y(n2323) );
  NAND2X1 U2845 ( .A(n2339), .B(n2340), .Y(n8356) );
  AOI22X1 U2846 ( .A(n2341), .B(n2342), .C(n11382), .D(n9370), .Y(n2340) );
  OAI21X1 U2847 ( .A(n9365), .B(n2343), .C(n2344), .Y(n2342) );
  AOI22X1 U2848 ( .A(n2345), .B(n2307), .C(n11363), .D(n9440), .Y(n2344) );
  OAI21X1 U2850 ( .A(n9393), .B(n2309), .C(n2347), .Y(n2346) );
  AOI22X1 U2851 ( .A(n2273), .B(n2348), .C(n11416), .D(n9474), .Y(n2347) );
  OAI22X1 U2852 ( .A(n9398), .B(n2237), .C(n11467), .D(n2349), .Y(n2348) );
  AOI22X1 U2853 ( .A(n11400), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[54] ), .D(n2351), .Y(n2349) );
  NAND2X1 U2855 ( .A(n2336), .B(n11410), .Y(n2351) );
  NAND2X1 U2857 ( .A(n2320), .B(n11478), .Y(n2237) );
  NOR2X1 U2858 ( .A(n11485), .B(n11416), .Y(n2273) );
  AOI22X1 U2859 ( .A(n11465), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[54] ), .D(n9441), .Y(n2339) );
  NAND2X1 U2860 ( .A(n2354), .B(n2355), .Y(n8357) );
  AOI22X1 U2861 ( .A(n2356), .B(n2357), .C(n11465), .D(n9370), .Y(n2355) );
  OAI21X1 U2862 ( .A(n9365), .B(n2358), .C(n2359), .Y(n2357) );
  AOI22X1 U2863 ( .A(n2360), .B(n2325), .C(n11434), .D(n9440), .Y(n2359) );
  OAI21X1 U2865 ( .A(n9393), .B(n2327), .C(n2362), .Y(n2361) );
  AOI22X1 U2866 ( .A(n2291), .B(n2363), .C(n11485), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2362) );
  OAI22X1 U2867 ( .A(n9398), .B(n2293), .C(n11416), .D(n2364), .Y(n2363) );
  AOI22X1 U2868 ( .A(n11468), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[53] ), .D(n2366), .Y(n2364) );
  NAND2X1 U2870 ( .A(n2336), .B(n11478), .Y(n2366) );
  NAND2X1 U2872 ( .A(n2320), .B(n11427), .Y(n2293) );
  NOR2X1 U2873 ( .A(n11363), .B(n11485), .Y(n2291) );
  AOI22X1 U2874 ( .A(n11414), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[53] ), .D(n9441), .Y(n2354) );
  NAND2X1 U2875 ( .A(n2369), .B(n2370), .Y(n8358) );
  AOI22X1 U2876 ( .A(n2371), .B(n2372), .C(n11414), .D(n9370), .Y(n2370) );
  OAI21X1 U2877 ( .A(n9365), .B(n2373), .C(n2374), .Y(n2372) );
  AOI22X1 U2878 ( .A(n2375), .B(n2341), .C(n11382), .D(n9440), .Y(n2374) );
  OAI21X1 U2880 ( .A(n9393), .B(n2343), .C(n2377), .Y(n2376) );
  AOI22X1 U2881 ( .A(n2307), .B(n2378), .C(n11363), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2377) );
  OAI22X1 U2882 ( .A(n9398), .B(n2309), .C(n11485), .D(n2379), .Y(n2378) );
  AOI22X1 U2883 ( .A(n11417), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[52] ), .D(n2381), .Y(n2379) );
  NAND2X1 U2885 ( .A(n2336), .B(n11427), .Y(n2381) );
  NAND2X1 U2887 ( .A(n2320), .B(n11496), .Y(n2309) );
  NOR2X1 U2888 ( .A(n11434), .B(n11363), .Y(n2307) );
  AOI22X1 U2889 ( .A(n11482), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[52] ), .D(n9441), .Y(n2369) );
  NAND2X1 U2890 ( .A(n2384), .B(n2385), .Y(n8359) );
  AOI22X1 U2891 ( .A(n2386), .B(n2387), .C(n11482), .D(n9370), .Y(n2385) );
  OAI21X1 U2892 ( .A(n9365), .B(n2388), .C(n2389), .Y(n2387) );
  AOI22X1 U2893 ( .A(n2390), .B(n2356), .C(n11465), .D(n9440), .Y(n2389) );
  OAI21X1 U2895 ( .A(n9393), .B(n2358), .C(n2392), .Y(n2391) );
  AOI22X1 U2896 ( .A(n2325), .B(n2393), .C(n11434), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2392) );
  OAI22X1 U2897 ( .A(n9398), .B(n2327), .C(n11363), .D(n2394), .Y(n2393) );
  AOI22X1 U2898 ( .A(n11486), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[51] ), .D(n2396), .Y(n2394) );
  NAND2X1 U2900 ( .A(n2336), .B(n11496), .Y(n2396) );
  NAND2X1 U2902 ( .A(n2320), .B(n11374), .Y(n2327) );
  NOR2X1 U2903 ( .A(n11382), .B(n11434), .Y(n2325) );
  AOI22X1 U2904 ( .A(n11431), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[51] ), .D(n9441), .Y(n2384) );
  NAND2X1 U2905 ( .A(n2399), .B(n2400), .Y(n8360) );
  AOI22X1 U2906 ( .A(n2401), .B(n2402), .C(n11431), .D(n9370), .Y(n2400) );
  OAI21X1 U2907 ( .A(n9365), .B(n2403), .C(n2404), .Y(n2402) );
  AOI22X1 U2908 ( .A(n2405), .B(n2371), .C(n11414), .D(n9440), .Y(n2404) );
  OAI21X1 U2910 ( .A(n9393), .B(n2373), .C(n2407), .Y(n2406) );
  AOI22X1 U2911 ( .A(n2341), .B(n2408), .C(n11382), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2407) );
  OAI22X1 U2912 ( .A(n9398), .B(n2343), .C(n11434), .D(n2409), .Y(n2408) );
  AOI22X1 U2913 ( .A(n11364), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[50] ), .D(n2411), .Y(n2409) );
  NAND2X1 U2915 ( .A(n2336), .B(n11374), .Y(n2411) );
  NAND2X1 U2917 ( .A(n2320), .B(n11445), .Y(n2343) );
  NOR2X1 U2918 ( .A(n11465), .B(n11382), .Y(n2341) );
  AOI22X1 U2919 ( .A(n11500), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[50] ), .D(n9441), .Y(n2399) );
  NAND2X1 U2920 ( .A(n2414), .B(n2415), .Y(n8361) );
  AOI22X1 U2921 ( .A(n2416), .B(n2417), .C(n11500), .D(n9370), .Y(n2415) );
  OAI21X1 U2922 ( .A(n9365), .B(n2418), .C(n2419), .Y(n2417) );
  AOI22X1 U2923 ( .A(n2420), .B(n2386), .C(n11482), .D(n9440), .Y(n2419) );
  OAI21X1 U2925 ( .A(n9393), .B(n2388), .C(n2422), .Y(n2421) );
  AOI22X1 U2926 ( .A(n2356), .B(n2423), .C(n11465), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2422) );
  OAI22X1 U2927 ( .A(n9398), .B(n2358), .C(n11382), .D(n2424), .Y(n2423) );
  AOI22X1 U2928 ( .A(n11435), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[49] ), .D(n2426), .Y(n2424) );
  NAND2X1 U2930 ( .A(n2336), .B(n11445), .Y(n2426) );
  NAND2X1 U2932 ( .A(n2320), .B(n11393), .Y(n2358) );
  NOR2X1 U2935 ( .A(n11414), .B(n11465), .Y(n2356) );
  AOI22X1 U2936 ( .A(n11378), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[49] ), .D(n9441), .Y(n2414) );
  NAND2X1 U2937 ( .A(n2431), .B(n2432), .Y(n8362) );
  AOI22X1 U2938 ( .A(n2433), .B(n2434), .C(n11378), .D(n9371), .Y(n2432) );
  OAI21X1 U2939 ( .A(n9365), .B(n2435), .C(n2436), .Y(n2434) );
  AOI22X1 U2940 ( .A(n2437), .B(n2401), .C(n11431), .D(n9440), .Y(n2436) );
  OAI21X1 U2942 ( .A(n9393), .B(n2403), .C(n2439), .Y(n2438) );
  AOI22X1 U2943 ( .A(n2371), .B(n2440), .C(n11414), .D(n9474), .Y(n2439) );
  OAI22X1 U2944 ( .A(n9398), .B(n2373), .C(n11465), .D(n2441), .Y(n2440) );
  AOI22X1 U2945 ( .A(n11383), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[48] ), .D(n2443), .Y(n2441) );
  NAND2X1 U2947 ( .A(n2336), .B(n11393), .Y(n2443) );
  NAND2X1 U2950 ( .A(n2444), .B(n2445), .Y(n2373) );
  NOR2X1 U2951 ( .A(n11482), .B(n11414), .Y(n2371) );
  AOI22X1 U2952 ( .A(n11449), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[48] ), .D(n2200), .Y(n2431) );
  NAND2X1 U2953 ( .A(n2447), .B(n2448), .Y(n8363) );
  AOI22X1 U2954 ( .A(n2449), .B(n2450), .C(n11449), .D(n9371), .Y(n2448) );
  OAI21X1 U2955 ( .A(n9365), .B(n2451), .C(n2452), .Y(n2450) );
  AOI22X1 U2956 ( .A(n2453), .B(n2416), .C(n11500), .D(n9440), .Y(n2452) );
  OAI21X1 U2958 ( .A(n9394), .B(n2418), .C(n2455), .Y(n2454) );
  AOI22X1 U2959 ( .A(n2386), .B(n2456), .C(n11482), .D(n9474), .Y(n2455) );
  OAI22X1 U2960 ( .A(n9398), .B(n2388), .C(n11414), .D(n2457), .Y(n2456) );
  AOI22X1 U2961 ( .A(n11452), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[47] ), .D(n2459), .Y(n2457) );
  NAND2X1 U2963 ( .A(n2460), .B(n11461), .Y(n2459) );
  NAND2X1 U2965 ( .A(n2444), .B(n2192), .Y(n2388) );
  NOR2X1 U2966 ( .A(n11431), .B(n11482), .Y(n2386) );
  AOI22X1 U2967 ( .A(n11396), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[47] ), .D(n9443), .Y(n2447) );
  NAND2X1 U2968 ( .A(n2462), .B(n2463), .Y(n8364) );
  AOI22X1 U2969 ( .A(n2464), .B(n2465), .C(n11396), .D(n9371), .Y(n2463) );
  OAI21X1 U2970 ( .A(n9366), .B(n2466), .C(n2467), .Y(n2465) );
  AOI22X1 U2971 ( .A(n2468), .B(n2433), .C(n11378), .D(n9440), .Y(n2467) );
  OAI21X1 U2973 ( .A(n9394), .B(n2435), .C(n2470), .Y(n2469) );
  AOI22X1 U2974 ( .A(n2401), .B(n2471), .C(n11431), .D(n9474), .Y(n2470) );
  OAI22X1 U2975 ( .A(n9400), .B(n2403), .C(n11482), .D(n2472), .Y(n2471) );
  AOI22X1 U2976 ( .A(n11401), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[46] ), .D(n2474), .Y(n2472) );
  NAND2X1 U2978 ( .A(n2460), .B(n11410), .Y(n2474) );
  NAND2X1 U2980 ( .A(n2444), .B(n2215), .Y(n2403) );
  NOR2X1 U2981 ( .A(n11500), .B(n11431), .Y(n2401) );
  AOI22X1 U2982 ( .A(n11453), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[46] ), .D(n9443), .Y(n2462) );
  NAND2X1 U2983 ( .A(n2476), .B(n2477), .Y(n8365) );
  AOI22X1 U2984 ( .A(n2478), .B(n2479), .C(n11453), .D(n9371), .Y(n2477) );
  OAI21X1 U2985 ( .A(n9366), .B(n2480), .C(n2481), .Y(n2479) );
  AOI22X1 U2986 ( .A(n2482), .B(n2449), .C(n11449), .D(n9440), .Y(n2481) );
  OAI21X1 U2988 ( .A(n9395), .B(n2451), .C(n2484), .Y(n2483) );
  AOI22X1 U2989 ( .A(n2416), .B(n2485), .C(n11500), .D(n9474), .Y(n2484) );
  OAI22X1 U2990 ( .A(n9399), .B(n2418), .C(n11431), .D(n2486), .Y(n2485) );
  AOI22X1 U2991 ( .A(n11469), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[45] ), .D(n2488), .Y(n2486) );
  NAND2X1 U2993 ( .A(n2460), .B(n11478), .Y(n2488) );
  NAND2X1 U2995 ( .A(n2444), .B(n2229), .Y(n2418) );
  NOR2X1 U2996 ( .A(n11378), .B(n11500), .Y(n2416) );
  AOI22X1 U2997 ( .A(n11402), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[45] ), .D(n9443), .Y(n2476) );
  NAND2X1 U2998 ( .A(n2490), .B(n2491), .Y(n8366) );
  AOI22X1 U2999 ( .A(n2492), .B(n2493), .C(n11402), .D(n9371), .Y(n2491) );
  OAI21X1 U3000 ( .A(n9366), .B(n2494), .C(n2495), .Y(n2493) );
  AOI22X1 U3001 ( .A(n2496), .B(n2464), .C(n11396), .D(n9440), .Y(n2495) );
  OAI21X1 U3003 ( .A(n9394), .B(n2466), .C(n2498), .Y(n2497) );
  AOI22X1 U3004 ( .A(n2433), .B(n2499), .C(n11378), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2498) );
  OAI22X1 U3005 ( .A(n9399), .B(n2435), .C(n11500), .D(n2500), .Y(n2499) );
  AOI22X1 U3006 ( .A(n11418), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[44] ), .D(n2502), .Y(n2500) );
  NAND2X1 U3008 ( .A(n2460), .B(n11427), .Y(n2502) );
  NAND2X1 U3010 ( .A(n2444), .B(n2250), .Y(n2435) );
  NOR2X1 U3011 ( .A(n11449), .B(n11378), .Y(n2433) );
  AOI22X1 U3012 ( .A(n11470), .B(n9448), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[44] ), .D(n9443), .Y(n2490) );
  NAND2X1 U3013 ( .A(n2504), .B(n2505), .Y(n8367) );
  AOI22X1 U3014 ( .A(n2506), .B(n2507), .C(n11470), .D(n9371), .Y(n2505) );
  OAI21X1 U3015 ( .A(n9366), .B(n2508), .C(n2509), .Y(n2507) );
  AOI22X1 U3016 ( .A(n2510), .B(n2478), .C(n11453), .D(n9440), .Y(n2509) );
  OAI21X1 U3018 ( .A(n9394), .B(n2480), .C(n2512), .Y(n2511) );
  AOI22X1 U3019 ( .A(n2449), .B(n2513), .C(n11449), .D(n9474), .Y(n2512) );
  OAI22X1 U3020 ( .A(n9399), .B(n2451), .C(n11378), .D(n2514), .Y(n2513) );
  AOI22X1 U3021 ( .A(n11487), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[43] ), .D(n2516), .Y(n2514) );
  NAND2X1 U3023 ( .A(n2460), .B(n11496), .Y(n2516) );
  NAND2X1 U3025 ( .A(n2444), .B(n2267), .Y(n2451) );
  NOR2X1 U3026 ( .A(n11396), .B(n11449), .Y(n2449) );
  AOI22X1 U3027 ( .A(n11419), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[43] ), .D(n9443), .Y(n2504) );
  NAND2X1 U3028 ( .A(n2518), .B(n2519), .Y(n8368) );
  AOI22X1 U3029 ( .A(n2520), .B(n2521), .C(n11419), .D(n9371), .Y(n2519) );
  OAI21X1 U3030 ( .A(n9366), .B(n2522), .C(n2523), .Y(n2521) );
  AOI22X1 U3031 ( .A(n2524), .B(n2492), .C(n11402), .D(n9439), .Y(n2523) );
  OAI21X1 U3033 ( .A(n9394), .B(n2494), .C(n2526), .Y(n2525) );
  AOI22X1 U3034 ( .A(n2464), .B(n2527), .C(n11396), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2526) );
  OAI22X1 U3035 ( .A(n9399), .B(n2466), .C(n11449), .D(n2528), .Y(n2527) );
  AOI22X1 U3036 ( .A(n11365), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[42] ), .D(n2530), .Y(n2528) );
  NAND2X1 U3038 ( .A(n2460), .B(n11374), .Y(n2530) );
  NAND2X1 U3040 ( .A(n2444), .B(n2287), .Y(n2466) );
  NOR2X1 U3041 ( .A(n11453), .B(n11396), .Y(n2464) );
  AOI22X1 U3042 ( .A(n11488), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[42] ), .D(n9443), .Y(n2518) );
  NAND2X1 U3043 ( .A(n2532), .B(n2533), .Y(n8369) );
  AOI22X1 U3044 ( .A(n2534), .B(n2535), .C(n11488), .D(n9371), .Y(n2533) );
  OAI21X1 U3045 ( .A(n9366), .B(n2536), .C(n2537), .Y(n2535) );
  AOI22X1 U3046 ( .A(n2538), .B(n2506), .C(n11470), .D(n9439), .Y(n2537) );
  OAI21X1 U3048 ( .A(n9394), .B(n2508), .C(n2540), .Y(n2539) );
  AOI22X1 U3049 ( .A(n2478), .B(n2541), .C(n11453), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2540) );
  OAI22X1 U3050 ( .A(n9399), .B(n2480), .C(n11396), .D(n2542), .Y(n2541) );
  AOI22X1 U3051 ( .A(n11436), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[41] ), .D(n2544), .Y(n2542) );
  NAND2X1 U3053 ( .A(n2460), .B(n11445), .Y(n2544) );
  NAND2X1 U3055 ( .A(n2444), .B(n2301), .Y(n2480) );
  NOR2X1 U3056 ( .A(n11402), .B(n11453), .Y(n2478) );
  AOI22X1 U3057 ( .A(n11366), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[41] ), .D(n9443), .Y(n2532) );
  NAND2X1 U3058 ( .A(n2546), .B(n2547), .Y(n8370) );
  AOI22X1 U3059 ( .A(n2548), .B(n2549), .C(n11366), .D(n9371), .Y(n2547) );
  OAI21X1 U3060 ( .A(n9366), .B(n2550), .C(n2551), .Y(n2549) );
  AOI22X1 U3061 ( .A(n2552), .B(n2520), .C(n11419), .D(n9439), .Y(n2551) );
  OAI21X1 U3063 ( .A(n9394), .B(n2522), .C(n2554), .Y(n2553) );
  AOI22X1 U3064 ( .A(n2492), .B(n2555), .C(n11402), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2554) );
  OAI22X1 U3065 ( .A(n9399), .B(n2494), .C(n11453), .D(n2556), .Y(n2555) );
  AOI22X1 U3066 ( .A(n11384), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[40] ), .D(n2558), .Y(n2556) );
  NAND2X1 U3068 ( .A(n2460), .B(n11393), .Y(n2558) );
  NAND2X1 U3071 ( .A(n2560), .B(n11461), .Y(n2494) );
  NOR2X1 U3072 ( .A(n11470), .B(n11402), .Y(n2492) );
  AOI22X1 U3073 ( .A(n11437), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[40] ), .D(n9443), .Y(n2546) );
  NAND2X1 U3074 ( .A(n2562), .B(n2563), .Y(n8371) );
  AOI22X1 U3075 ( .A(n2564), .B(n2565), .C(n11437), .D(n9371), .Y(n2563) );
  OAI21X1 U3076 ( .A(n9366), .B(n2566), .C(n2567), .Y(n2565) );
  AOI22X1 U3077 ( .A(n2568), .B(n2534), .C(n11488), .D(n9439), .Y(n2567) );
  OAI21X1 U3079 ( .A(n9394), .B(n2536), .C(n2570), .Y(n2569) );
  AOI22X1 U3080 ( .A(n2506), .B(n2571), .C(n11470), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2570) );
  OAI22X1 U3081 ( .A(n9399), .B(n2508), .C(n11402), .D(n2572), .Y(n2571) );
  AOI22X1 U3082 ( .A(n11454), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[39] ), .D(n2574), .Y(n2572) );
  NAND2X1 U3084 ( .A(n2575), .B(n11461), .Y(n2574) );
  NAND2X1 U3086 ( .A(n2560), .B(n11410), .Y(n2508) );
  NOR2X1 U3087 ( .A(n11419), .B(n11470), .Y(n2506) );
  AOI22X1 U3088 ( .A(n11385), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[39] ), .D(n9443), .Y(n2562) );
  NAND2X1 U3089 ( .A(n2577), .B(n2578), .Y(n8372) );
  AOI22X1 U3090 ( .A(n2579), .B(n2580), .C(n11385), .D(n9371), .Y(n2578) );
  OAI21X1 U3091 ( .A(n9366), .B(n2581), .C(n2582), .Y(n2580) );
  AOI22X1 U3092 ( .A(n2583), .B(n2548), .C(n11366), .D(n9439), .Y(n2582) );
  OAI21X1 U3094 ( .A(n9394), .B(n2550), .C(n2585), .Y(n2584) );
  AOI22X1 U3095 ( .A(n2520), .B(n2586), .C(n11419), .D(
        \U_1/U_0/U_1/RCV_DATA [2]), .Y(n2585) );
  OAI22X1 U3096 ( .A(n9399), .B(n2522), .C(n11470), .D(n2587), .Y(n2586) );
  AOI22X1 U3097 ( .A(n11403), .B(\U_1/U_0/U_1/RCV_DATA [0]), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[38] ), .D(n2589), .Y(n2587) );
  NAND2X1 U3099 ( .A(n2575), .B(n11410), .Y(n2589) );
  NAND2X1 U3101 ( .A(n2560), .B(n11478), .Y(n2522) );
  NOR2X1 U3102 ( .A(n11488), .B(n11419), .Y(n2520) );
  AOI22X1 U3103 ( .A(n11464), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[38] ), .D(n9443), .Y(n2577) );
  NAND2X1 U3104 ( .A(n2591), .B(n2592), .Y(n8373) );
  AOI22X1 U3105 ( .A(n2593), .B(n2594), .C(n11464), .D(n9371), .Y(n2592) );
  OAI21X1 U3106 ( .A(n9366), .B(n2595), .C(n2596), .Y(n2594) );
  AOI22X1 U3107 ( .A(n2597), .B(n2564), .C(n11437), .D(n9439), .Y(n2596) );
  OAI21X1 U3109 ( .A(n9394), .B(n2566), .C(n2599), .Y(n2598) );
  AOI22X1 U3110 ( .A(n2534), .B(n2600), .C(n11488), .D(n9474), .Y(n2599) );
  OAI22X1 U3111 ( .A(n9399), .B(n2536), .C(n11419), .D(n2601), .Y(n2600) );
  AOI22X1 U3112 ( .A(n11471), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[37] ), .D(n2603), .Y(n2601) );
  NAND2X1 U3114 ( .A(n2575), .B(n11478), .Y(n2603) );
  NAND2X1 U3116 ( .A(n2560), .B(n11427), .Y(n2536) );
  NOR2X1 U3117 ( .A(n11366), .B(n11488), .Y(n2534) );
  AOI22X1 U3118 ( .A(n11413), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[37] ), .D(n9443), .Y(n2591) );
  NAND2X1 U3119 ( .A(n2605), .B(n2606), .Y(n8374) );
  AOI22X1 U3120 ( .A(n2607), .B(n2608), .C(n11413), .D(n9371), .Y(n2606) );
  OAI21X1 U3121 ( .A(n9366), .B(n2609), .C(n2610), .Y(n2608) );
  AOI22X1 U3122 ( .A(n2611), .B(n2579), .C(n11385), .D(n9439), .Y(n2610) );
  OAI21X1 U3124 ( .A(n9394), .B(n2581), .C(n2613), .Y(n2612) );
  AOI22X1 U3125 ( .A(n2548), .B(n2614), .C(n11366), .D(n9474), .Y(n2613) );
  OAI22X1 U3126 ( .A(n9399), .B(n2550), .C(n11488), .D(n2615), .Y(n2614) );
  AOI22X1 U3127 ( .A(n11420), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[36] ), .D(n2617), .Y(n2615) );
  NAND2X1 U3129 ( .A(n2575), .B(n11427), .Y(n2617) );
  NAND2X1 U3131 ( .A(n2560), .B(n11496), .Y(n2550) );
  NOR2X1 U3132 ( .A(n11437), .B(n11366), .Y(n2548) );
  AOI22X1 U3133 ( .A(n11481), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[36] ), .D(n9443), .Y(n2605) );
  NAND2X1 U3134 ( .A(n2619), .B(n2620), .Y(n8375) );
  AOI22X1 U3135 ( .A(n2621), .B(n2622), .C(n11481), .D(n9372), .Y(n2620) );
  OAI21X1 U3136 ( .A(n9366), .B(n2623), .C(n2624), .Y(n2622) );
  AOI22X1 U3137 ( .A(n2625), .B(n2593), .C(n11464), .D(n9439), .Y(n2624) );
  OAI21X1 U3139 ( .A(n9394), .B(n2595), .C(n2627), .Y(n2626) );
  AOI22X1 U3140 ( .A(n2564), .B(n2628), .C(n11437), .D(n9474), .Y(n2627) );
  OAI22X1 U3141 ( .A(n9399), .B(n2566), .C(n11366), .D(n2629), .Y(n2628) );
  AOI22X1 U3142 ( .A(n11489), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[35] ), .D(n2631), .Y(n2629) );
  NAND2X1 U3144 ( .A(n2575), .B(n11496), .Y(n2631) );
  NAND2X1 U3146 ( .A(n2560), .B(n11374), .Y(n2566) );
  NOR2X1 U3147 ( .A(n11385), .B(n11437), .Y(n2564) );
  AOI22X1 U3148 ( .A(n11430), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[35] ), .D(n9443), .Y(n2619) );
  NAND2X1 U3149 ( .A(n2633), .B(n2634), .Y(n8376) );
  AOI22X1 U3150 ( .A(n2635), .B(n2636), .C(n11430), .D(n9372), .Y(n2634) );
  OAI21X1 U3151 ( .A(n9366), .B(n2637), .C(n2638), .Y(n2636) );
  AOI22X1 U3152 ( .A(n2639), .B(n2607), .C(n11413), .D(n9439), .Y(n2638) );
  OAI21X1 U3154 ( .A(n9394), .B(n2609), .C(n2641), .Y(n2640) );
  AOI22X1 U3155 ( .A(n2579), .B(n2642), .C(n11385), .D(n9474), .Y(n2641) );
  OAI22X1 U3156 ( .A(n9399), .B(n2581), .C(n11437), .D(n2643), .Y(n2642) );
  AOI22X1 U3157 ( .A(n11367), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[34] ), .D(n2645), .Y(n2643) );
  NAND2X1 U3159 ( .A(n2575), .B(n11374), .Y(n2645) );
  NAND2X1 U3161 ( .A(n2560), .B(n11445), .Y(n2581) );
  NOR2X1 U3162 ( .A(n11464), .B(n11385), .Y(n2579) );
  AOI22X1 U3163 ( .A(n11499), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[34] ), .D(n2200), .Y(n2633) );
  NAND2X1 U3164 ( .A(n2647), .B(n2648), .Y(n8377) );
  AOI22X1 U3165 ( .A(n2649), .B(n2650), .C(n11499), .D(n9372), .Y(n2648) );
  OAI21X1 U3166 ( .A(n9367), .B(n2651), .C(n2652), .Y(n2650) );
  AOI22X1 U3167 ( .A(n2653), .B(n2621), .C(n11481), .D(n9439), .Y(n2652) );
  OAI21X1 U3169 ( .A(n9395), .B(n2623), .C(n2655), .Y(n2654) );
  AOI22X1 U3170 ( .A(n2593), .B(n2656), .C(n11464), .D(n9474), .Y(n2655) );
  OAI22X1 U3171 ( .A(n9399), .B(n2595), .C(n11385), .D(n2657), .Y(n2656) );
  AOI22X1 U3172 ( .A(n11438), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[33] ), .D(n2659), .Y(n2657) );
  NAND2X1 U3174 ( .A(n2575), .B(n11445), .Y(n2659) );
  NAND2X1 U3176 ( .A(n2560), .B(n11393), .Y(n2595) );
  NOR2X1 U3179 ( .A(n11413), .B(n11464), .Y(n2593) );
  AOI22X1 U3180 ( .A(n11377), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[33] ), .D(n2200), .Y(n2647) );
  NAND2X1 U3181 ( .A(n2661), .B(n2662), .Y(n8378) );
  AOI22X1 U3182 ( .A(n2663), .B(n2664), .C(n11377), .D(n9372), .Y(n2662) );
  OAI21X1 U3183 ( .A(n9367), .B(n2665), .C(n2666), .Y(n2664) );
  AOI22X1 U3184 ( .A(n2667), .B(n2635), .C(n11430), .D(n9439), .Y(n2666) );
  OAI21X1 U3186 ( .A(n9395), .B(n2637), .C(n2669), .Y(n2668) );
  AOI22X1 U3187 ( .A(n2607), .B(n2670), .C(n11413), .D(n9474), .Y(n2669) );
  OAI22X1 U3188 ( .A(n9400), .B(n2609), .C(n11464), .D(n2671), .Y(n2670) );
  AOI22X1 U3189 ( .A(n11386), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[32] ), .D(n2673), .Y(n2671) );
  NAND2X1 U3191 ( .A(n2575), .B(n11393), .Y(n2673) );
  NOR2X1 U3193 ( .A(n11510), .B(\U_1/U_0/U_1/U_8/address[4] ), .Y(n2559) );
  NAND2X1 U3195 ( .A(n2675), .B(n2445), .Y(n2609) );
  NOR2X1 U3196 ( .A(n11481), .B(n11413), .Y(n2607) );
  AOI22X1 U3197 ( .A(n11448), .B(n9449), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[32] ), .D(n2200), .Y(n2661) );
  NAND2X1 U3198 ( .A(n2677), .B(n2678), .Y(n8379) );
  AOI22X1 U3199 ( .A(n2679), .B(n2680), .C(n11448), .D(n9372), .Y(n2678) );
  OAI21X1 U3200 ( .A(n9367), .B(n2681), .C(n2682), .Y(n2680) );
  AOI22X1 U3201 ( .A(n2683), .B(n2649), .C(n11499), .D(n9439), .Y(n2682) );
  OAI21X1 U3203 ( .A(n9395), .B(n2651), .C(n2685), .Y(n2684) );
  AOI22X1 U3204 ( .A(n2621), .B(n2686), .C(n11481), .D(n9474), .Y(n2685) );
  OAI22X1 U3205 ( .A(n9400), .B(n2623), .C(n11413), .D(n2687), .Y(n2686) );
  AOI22X1 U3206 ( .A(n11455), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[31] ), .D(n2689), .Y(n2687) );
  NAND2X1 U3208 ( .A(n2690), .B(n11461), .Y(n2689) );
  NAND2X1 U3210 ( .A(n2675), .B(n2192), .Y(n2623) );
  NOR2X1 U3211 ( .A(n11430), .B(n11481), .Y(n2621) );
  AOI22X1 U3212 ( .A(n11395), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[31] ), .D(n2200), .Y(n2677) );
  NAND2X1 U3213 ( .A(n2692), .B(n2693), .Y(n8380) );
  AOI22X1 U3214 ( .A(n2694), .B(n2695), .C(n11395), .D(n9372), .Y(n2693) );
  OAI21X1 U3215 ( .A(n9367), .B(n2696), .C(n2697), .Y(n2695) );
  AOI22X1 U3216 ( .A(n2698), .B(n2663), .C(n11377), .D(n9439), .Y(n2697) );
  OAI21X1 U3218 ( .A(n9395), .B(n2665), .C(n2700), .Y(n2699) );
  AOI22X1 U3219 ( .A(n2635), .B(n2701), .C(n11430), .D(n9474), .Y(n2700) );
  OAI22X1 U3220 ( .A(n9400), .B(n2637), .C(n11481), .D(n2702), .Y(n2701) );
  AOI22X1 U3221 ( .A(n11404), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[30] ), .D(n2704), .Y(n2702) );
  NAND2X1 U3223 ( .A(n2690), .B(n11410), .Y(n2704) );
  NAND2X1 U3225 ( .A(n2675), .B(n2215), .Y(n2637) );
  NOR2X1 U3226 ( .A(n11499), .B(n11430), .Y(n2635) );
  AOI22X1 U3227 ( .A(n11456), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[30] ), .D(n9441), .Y(n2692) );
  NAND2X1 U3228 ( .A(n2706), .B(n2707), .Y(n8381) );
  AOI22X1 U3229 ( .A(n2708), .B(n2709), .C(n11456), .D(n9372), .Y(n2707) );
  OAI21X1 U3230 ( .A(n9367), .B(n2710), .C(n2711), .Y(n2709) );
  AOI22X1 U3231 ( .A(n2712), .B(n2679), .C(n11448), .D(n9438), .Y(n2711) );
  OAI21X1 U3233 ( .A(n9395), .B(n2681), .C(n2714), .Y(n2713) );
  AOI22X1 U3234 ( .A(n2649), .B(n2715), .C(n11499), .D(n9474), .Y(n2714) );
  OAI22X1 U3235 ( .A(n9400), .B(n2651), .C(n11430), .D(n2716), .Y(n2715) );
  AOI22X1 U3236 ( .A(n11472), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[29] ), .D(n2718), .Y(n2716) );
  NAND2X1 U3238 ( .A(n2690), .B(n11478), .Y(n2718) );
  NAND2X1 U3240 ( .A(n2675), .B(n2229), .Y(n2651) );
  NOR2X1 U3241 ( .A(n11377), .B(n11499), .Y(n2649) );
  AOI22X1 U3242 ( .A(n11405), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[29] ), .D(n2200), .Y(n2706) );
  NAND2X1 U3243 ( .A(n2720), .B(n2721), .Y(n8382) );
  AOI22X1 U3244 ( .A(n2722), .B(n2723), .C(n11405), .D(n9372), .Y(n2721) );
  OAI21X1 U3245 ( .A(n9367), .B(n2724), .C(n2725), .Y(n2723) );
  AOI22X1 U3246 ( .A(n2726), .B(n2694), .C(n11395), .D(n9438), .Y(n2725) );
  OAI21X1 U3248 ( .A(n9395), .B(n2696), .C(n2728), .Y(n2727) );
  AOI22X1 U3249 ( .A(n2663), .B(n2729), .C(n11377), .D(n9474), .Y(n2728) );
  OAI22X1 U3250 ( .A(n9400), .B(n2665), .C(n11499), .D(n2730), .Y(n2729) );
  AOI22X1 U3251 ( .A(n11421), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[28] ), .D(n2732), .Y(n2730) );
  NAND2X1 U3253 ( .A(n2690), .B(n11427), .Y(n2732) );
  NAND2X1 U3255 ( .A(n2675), .B(n2250), .Y(n2665) );
  NOR2X1 U3256 ( .A(n11448), .B(n11377), .Y(n2663) );
  AOI22X1 U3257 ( .A(n11473), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[28] ), .D(n9441), .Y(n2720) );
  NAND2X1 U3258 ( .A(n2734), .B(n2735), .Y(n8383) );
  AOI22X1 U3259 ( .A(n2736), .B(n2737), .C(n11473), .D(n9372), .Y(n2735) );
  OAI21X1 U3260 ( .A(n9367), .B(n2738), .C(n2739), .Y(n2737) );
  AOI22X1 U3261 ( .A(n2740), .B(n2708), .C(n11456), .D(n9440), .Y(n2739) );
  OAI21X1 U3263 ( .A(n9395), .B(n2710), .C(n2742), .Y(n2741) );
  AOI22X1 U3264 ( .A(n2679), .B(n2743), .C(n11448), .D(n9474), .Y(n2742) );
  OAI22X1 U3265 ( .A(n9400), .B(n2681), .C(n11377), .D(n2744), .Y(n2743) );
  AOI22X1 U3266 ( .A(n11490), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[27] ), .D(n2746), .Y(n2744) );
  NAND2X1 U3268 ( .A(n2690), .B(n11496), .Y(n2746) );
  NAND2X1 U3270 ( .A(n2675), .B(n2267), .Y(n2681) );
  NOR2X1 U3271 ( .A(n11395), .B(n11448), .Y(n2679) );
  AOI22X1 U3272 ( .A(n11422), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[27] ), .D(n2200), .Y(n2734) );
  NAND2X1 U3273 ( .A(n2748), .B(n2749), .Y(n8384) );
  AOI22X1 U3274 ( .A(n2750), .B(n2751), .C(n11422), .D(n9372), .Y(n2749) );
  OAI21X1 U3275 ( .A(n9367), .B(n2752), .C(n2753), .Y(n2751) );
  AOI22X1 U3276 ( .A(n2754), .B(n2722), .C(n11405), .D(n9439), .Y(n2753) );
  OAI21X1 U3278 ( .A(n9395), .B(n2724), .C(n2756), .Y(n2755) );
  AOI22X1 U3279 ( .A(n2694), .B(n2757), .C(n11395), .D(n9474), .Y(n2756) );
  OAI22X1 U3280 ( .A(n9400), .B(n2696), .C(n11448), .D(n2758), .Y(n2757) );
  AOI22X1 U3281 ( .A(n11368), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[26] ), .D(n2760), .Y(n2758) );
  NAND2X1 U3283 ( .A(n2690), .B(n11374), .Y(n2760) );
  NAND2X1 U3285 ( .A(n2675), .B(n2287), .Y(n2696) );
  NOR2X1 U3286 ( .A(n11456), .B(n11395), .Y(n2694) );
  AOI22X1 U3287 ( .A(n11491), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[26] ), .D(n9441), .Y(n2748) );
  NAND2X1 U3288 ( .A(n2762), .B(n2763), .Y(n8385) );
  AOI22X1 U3289 ( .A(n2764), .B(n2765), .C(n11491), .D(n9372), .Y(n2763) );
  OAI21X1 U3290 ( .A(n9367), .B(n2766), .C(n2767), .Y(n2765) );
  AOI22X1 U3291 ( .A(n2768), .B(n2736), .C(n11473), .D(n9440), .Y(n2767) );
  OAI21X1 U3293 ( .A(n9395), .B(n2738), .C(n2770), .Y(n2769) );
  AOI22X1 U3294 ( .A(n2708), .B(n2771), .C(n11456), .D(n9474), .Y(n2770) );
  OAI22X1 U3295 ( .A(n9400), .B(n2710), .C(n11395), .D(n2772), .Y(n2771) );
  AOI22X1 U3296 ( .A(n11439), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[25] ), .D(n2774), .Y(n2772) );
  NAND2X1 U3298 ( .A(n2690), .B(n11445), .Y(n2774) );
  NAND2X1 U3300 ( .A(n2675), .B(n2301), .Y(n2710) );
  NOR2X1 U3301 ( .A(n11405), .B(n11456), .Y(n2708) );
  AOI22X1 U3302 ( .A(n11369), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[25] ), .D(n9441), .Y(n2762) );
  NAND2X1 U3303 ( .A(n2776), .B(n2777), .Y(n8386) );
  AOI22X1 U3304 ( .A(n2778), .B(n2779), .C(n11369), .D(n9372), .Y(n2777) );
  OAI21X1 U3305 ( .A(n9367), .B(n2780), .C(n2781), .Y(n2779) );
  AOI22X1 U3306 ( .A(n2782), .B(n2750), .C(n11422), .D(n9438), .Y(n2781) );
  OAI21X1 U3308 ( .A(n9395), .B(n2752), .C(n2784), .Y(n2783) );
  AOI22X1 U3309 ( .A(n2722), .B(n2785), .C(n11405), .D(n9474), .Y(n2784) );
  OAI22X1 U3310 ( .A(n9400), .B(n2724), .C(n11456), .D(n2786), .Y(n2785) );
  AOI22X1 U3311 ( .A(n11387), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[24] ), .D(n2788), .Y(n2786) );
  NAND2X1 U3313 ( .A(n2690), .B(n11393), .Y(n2788) );
  NAND2X1 U3316 ( .A(n2790), .B(n11461), .Y(n2724) );
  NOR2X1 U3317 ( .A(n11473), .B(n11405), .Y(n2722) );
  AOI22X1 U3318 ( .A(n11440), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[24] ), .D(n9441), .Y(n2776) );
  NAND2X1 U3319 ( .A(n2792), .B(n2793), .Y(n8387) );
  AOI22X1 U3320 ( .A(n2794), .B(n2795), .C(n11440), .D(n9372), .Y(n2793) );
  OAI21X1 U3321 ( .A(n9367), .B(n2796), .C(n2797), .Y(n2795) );
  AOI22X1 U3322 ( .A(n2798), .B(n2764), .C(n11491), .D(n9439), .Y(n2797) );
  OAI21X1 U3324 ( .A(n9395), .B(n2766), .C(n2800), .Y(n2799) );
  AOI22X1 U3325 ( .A(n2736), .B(n2801), .C(n11473), .D(n9474), .Y(n2800) );
  OAI22X1 U3326 ( .A(n9400), .B(n2738), .C(n11405), .D(n2802), .Y(n2801) );
  AOI22X1 U3327 ( .A(n11457), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[23] ), .D(n2804), .Y(n2802) );
  NAND2X1 U3329 ( .A(n2805), .B(n11461), .Y(n2804) );
  NAND2X1 U3331 ( .A(n2790), .B(n11410), .Y(n2738) );
  NOR2X1 U3332 ( .A(n11422), .B(n11473), .Y(n2736) );
  AOI22X1 U3333 ( .A(n11388), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[23] ), .D(n9441), .Y(n2792) );
  NAND2X1 U3334 ( .A(n2807), .B(n2808), .Y(n8388) );
  AOI22X1 U3335 ( .A(n2809), .B(n2810), .C(n11388), .D(n9373), .Y(n2808) );
  OAI21X1 U3336 ( .A(n9367), .B(n2811), .C(n2812), .Y(n2810) );
  AOI22X1 U3337 ( .A(n2813), .B(n2778), .C(n11369), .D(n9440), .Y(n2812) );
  OAI21X1 U3339 ( .A(n9395), .B(n2780), .C(n2815), .Y(n2814) );
  AOI22X1 U3340 ( .A(n2750), .B(n2816), .C(n11422), .D(n9474), .Y(n2815) );
  OAI22X1 U3341 ( .A(n9400), .B(n2752), .C(n11473), .D(n2817), .Y(n2816) );
  AOI22X1 U3342 ( .A(n11406), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[22] ), .D(n2819), .Y(n2817) );
  NAND2X1 U3344 ( .A(n2805), .B(n11410), .Y(n2819) );
  NAND2X1 U3346 ( .A(n2790), .B(n11478), .Y(n2752) );
  NOR2X1 U3347 ( .A(n11491), .B(n11422), .Y(n2750) );
  AOI22X1 U3348 ( .A(n11463), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[22] ), .D(n9441), .Y(n2807) );
  NAND2X1 U3349 ( .A(n2821), .B(n2822), .Y(n8389) );
  AOI22X1 U3350 ( .A(n2823), .B(n2824), .C(n11463), .D(n9373), .Y(n2822) );
  OAI21X1 U3351 ( .A(n9367), .B(n2825), .C(n2826), .Y(n2824) );
  AOI22X1 U3352 ( .A(n2827), .B(n2794), .C(n11440), .D(n9438), .Y(n2826) );
  OAI21X1 U3354 ( .A(n9396), .B(n2796), .C(n2829), .Y(n2828) );
  AOI22X1 U3355 ( .A(n2764), .B(n2830), .C(n11491), .D(n9474), .Y(n2829) );
  OAI22X1 U3356 ( .A(n9400), .B(n2766), .C(n11422), .D(n2831), .Y(n2830) );
  AOI22X1 U3357 ( .A(n11474), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[21] ), .D(n2833), .Y(n2831) );
  NAND2X1 U3359 ( .A(n2805), .B(n11478), .Y(n2833) );
  NAND2X1 U3361 ( .A(n2790), .B(n11427), .Y(n2766) );
  NOR2X1 U3362 ( .A(n11369), .B(n11491), .Y(n2764) );
  AOI22X1 U3363 ( .A(n11412), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[21] ), .D(n9441), .Y(n2821) );
  NAND2X1 U3364 ( .A(n2835), .B(n2836), .Y(n8390) );
  AOI22X1 U3365 ( .A(n2837), .B(n2838), .C(n11412), .D(n9373), .Y(n2836) );
  OAI21X1 U3366 ( .A(n9368), .B(n2839), .C(n2840), .Y(n2838) );
  AOI22X1 U3367 ( .A(n2841), .B(n2809), .C(n11388), .D(n9439), .Y(n2840) );
  OAI21X1 U3369 ( .A(n9396), .B(n2811), .C(n2843), .Y(n2842) );
  AOI22X1 U3370 ( .A(n2778), .B(n2844), .C(n11369), .D(n9474), .Y(n2843) );
  OAI22X1 U3371 ( .A(n9401), .B(n2780), .C(n11491), .D(n2845), .Y(n2844) );
  AOI22X1 U3372 ( .A(n11423), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[20] ), .D(n2847), .Y(n2845) );
  NAND2X1 U3374 ( .A(n2805), .B(n11427), .Y(n2847) );
  NAND2X1 U3376 ( .A(n2790), .B(n11496), .Y(n2780) );
  NOR2X1 U3377 ( .A(n11440), .B(n11369), .Y(n2778) );
  AOI22X1 U3378 ( .A(n11480), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[20] ), .D(n9441), .Y(n2835) );
  NAND2X1 U3379 ( .A(n2849), .B(n2850), .Y(n8391) );
  AOI22X1 U3380 ( .A(n2851), .B(n2852), .C(n11480), .D(n9373), .Y(n2850) );
  OAI21X1 U3381 ( .A(n9368), .B(n2853), .C(n2854), .Y(n2852) );
  AOI22X1 U3382 ( .A(n2855), .B(n2823), .C(n11463), .D(n9440), .Y(n2854) );
  OAI21X1 U3384 ( .A(n9396), .B(n2825), .C(n2857), .Y(n2856) );
  AOI22X1 U3385 ( .A(n2794), .B(n2858), .C(n11440), .D(n9474), .Y(n2857) );
  OAI22X1 U3386 ( .A(n9401), .B(n2796), .C(n11369), .D(n2859), .Y(n2858) );
  AOI22X1 U3387 ( .A(n11492), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[19] ), .D(n2861), .Y(n2859) );
  NAND2X1 U3389 ( .A(n2805), .B(n11496), .Y(n2861) );
  NAND2X1 U3391 ( .A(n2790), .B(n11374), .Y(n2796) );
  NOR2X1 U3392 ( .A(n11388), .B(n11440), .Y(n2794) );
  AOI22X1 U3393 ( .A(n11429), .B(n9450), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[19] ), .D(n9441), .Y(n2849) );
  NAND2X1 U3394 ( .A(n2863), .B(n2864), .Y(n8392) );
  AOI22X1 U3395 ( .A(n2865), .B(n2866), .C(n11429), .D(n9373), .Y(n2864) );
  OAI21X1 U3396 ( .A(n9368), .B(n2867), .C(n2868), .Y(n2866) );
  AOI22X1 U3397 ( .A(n2869), .B(n2837), .C(n11412), .D(n9438), .Y(n2868) );
  OAI21X1 U3399 ( .A(n9396), .B(n2839), .C(n2871), .Y(n2870) );
  AOI22X1 U3400 ( .A(n2809), .B(n2872), .C(n11388), .D(n9474), .Y(n2871) );
  OAI22X1 U3401 ( .A(n9401), .B(n2811), .C(n11440), .D(n2873), .Y(n2872) );
  AOI22X1 U3402 ( .A(n11370), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[18] ), .D(n2875), .Y(n2873) );
  NAND2X1 U3404 ( .A(n2805), .B(n11374), .Y(n2875) );
  NAND2X1 U3406 ( .A(n2790), .B(n11445), .Y(n2811) );
  NOR2X1 U3407 ( .A(n11463), .B(n11388), .Y(n2809) );
  AOI22X1 U3408 ( .A(n11498), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[18] ), .D(n9441), .Y(n2863) );
  NAND2X1 U3409 ( .A(n2877), .B(n2878), .Y(n8393) );
  AOI22X1 U3410 ( .A(n2879), .B(n2880), .C(n11498), .D(n9373), .Y(n2878) );
  OAI21X1 U3411 ( .A(n9368), .B(n2881), .C(n2882), .Y(n2880) );
  AOI22X1 U3412 ( .A(n2883), .B(n2851), .C(n11480), .D(n9439), .Y(n2882) );
  OAI21X1 U3414 ( .A(n9396), .B(n2853), .C(n2885), .Y(n2884) );
  AOI22X1 U3415 ( .A(n2823), .B(n2886), .C(n11463), .D(n9474), .Y(n2885) );
  OAI22X1 U3416 ( .A(n9401), .B(n2825), .C(n11388), .D(n2887), .Y(n2886) );
  AOI22X1 U3417 ( .A(n11441), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[17] ), .D(n2889), .Y(n2887) );
  NAND2X1 U3419 ( .A(n2805), .B(n11445), .Y(n2889) );
  NAND2X1 U3421 ( .A(n2790), .B(n11393), .Y(n2825) );
  NOR2X1 U3424 ( .A(n11412), .B(n11463), .Y(n2823) );
  AOI22X1 U3425 ( .A(n11376), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[17] ), .D(n9441), .Y(n2877) );
  NAND2X1 U3426 ( .A(n2891), .B(n2892), .Y(n8394) );
  AOI22X1 U3427 ( .A(n2893), .B(n2894), .C(n11376), .D(n9373), .Y(n2892) );
  OAI21X1 U3428 ( .A(n9368), .B(n2895), .C(n2896), .Y(n2894) );
  AOI22X1 U3429 ( .A(n2897), .B(n2865), .C(n11429), .D(n9438), .Y(n2896) );
  OAI21X1 U3431 ( .A(n9396), .B(n2867), .C(n2899), .Y(n2898) );
  AOI22X1 U3432 ( .A(n2837), .B(n2900), .C(n11412), .D(n9474), .Y(n2899) );
  OAI22X1 U3433 ( .A(n9401), .B(n2839), .C(n11463), .D(n2901), .Y(n2900) );
  AOI22X1 U3434 ( .A(n11389), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[16] ), .D(n2903), .Y(n2901) );
  NAND2X1 U3436 ( .A(n2805), .B(n11393), .Y(n2903) );
  NOR2X1 U3438 ( .A(n11511), .B(\U_1/U_0/U_1/U_8/address[5] ), .Y(n2789) );
  NAND2X1 U3440 ( .A(n2905), .B(n2445), .Y(n2839) );
  NOR2X1 U3441 ( .A(n11480), .B(n11412), .Y(n2837) );
  AOI22X1 U3442 ( .A(n11447), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[16] ), .D(n9441), .Y(n2891) );
  NAND2X1 U3443 ( .A(n2907), .B(n2908), .Y(n8395) );
  AOI22X1 U3444 ( .A(n2909), .B(n2910), .C(n11447), .D(n9373), .Y(n2908) );
  OAI21X1 U3445 ( .A(n9368), .B(n2911), .C(n2912), .Y(n2910) );
  AOI22X1 U3446 ( .A(n2913), .B(n2879), .C(n11498), .D(n9438), .Y(n2912) );
  OAI21X1 U3448 ( .A(n9396), .B(n2881), .C(n2915), .Y(n2914) );
  AOI22X1 U3449 ( .A(n2851), .B(n2916), .C(n11480), .D(n9474), .Y(n2915) );
  OAI22X1 U3450 ( .A(n9401), .B(n2853), .C(n11412), .D(n2917), .Y(n2916) );
  AOI22X1 U3451 ( .A(n11458), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[15] ), .D(n2919), .Y(n2917) );
  NAND2X1 U3453 ( .A(n2920), .B(n11461), .Y(n2919) );
  NAND2X1 U3455 ( .A(n2905), .B(n2192), .Y(n2853) );
  NOR2X1 U3456 ( .A(n11429), .B(n11480), .Y(n2851) );
  AOI22X1 U3457 ( .A(n11394), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[15] ), .D(n9441), .Y(n2907) );
  NAND2X1 U3458 ( .A(n2922), .B(n2923), .Y(n8396) );
  AOI22X1 U3459 ( .A(n2924), .B(n2925), .C(n11394), .D(n9373), .Y(n2923) );
  OAI21X1 U3460 ( .A(n9368), .B(n2926), .C(n2927), .Y(n2925) );
  AOI22X1 U3461 ( .A(n2928), .B(n2893), .C(n11376), .D(n9438), .Y(n2927) );
  OAI21X1 U3463 ( .A(n9396), .B(n2895), .C(n2930), .Y(n2929) );
  AOI22X1 U3464 ( .A(n2865), .B(n2931), .C(n11429), .D(n9474), .Y(n2930) );
  OAI22X1 U3465 ( .A(n9401), .B(n2867), .C(n11480), .D(n2932), .Y(n2931) );
  AOI22X1 U3466 ( .A(n11407), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[14] ), .D(n2934), .Y(n2932) );
  NAND2X1 U3468 ( .A(n2920), .B(n11410), .Y(n2934) );
  NAND2X1 U3470 ( .A(n2905), .B(n2215), .Y(n2867) );
  NOR2X1 U3471 ( .A(n11498), .B(n11429), .Y(n2865) );
  AOI22X1 U3472 ( .A(n11459), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[14] ), .D(n2200), .Y(n2922) );
  NAND2X1 U3473 ( .A(n2936), .B(n2937), .Y(n8397) );
  AOI22X1 U3474 ( .A(n2938), .B(n2939), .C(n11459), .D(n9373), .Y(n2937) );
  OAI21X1 U3475 ( .A(n9368), .B(n2940), .C(n2941), .Y(n2939) );
  AOI22X1 U3476 ( .A(n2942), .B(n2909), .C(n11447), .D(n9438), .Y(n2941) );
  OAI21X1 U3478 ( .A(n9396), .B(n2911), .C(n2944), .Y(n2943) );
  AOI22X1 U3479 ( .A(n2879), .B(n2945), .C(n11498), .D(n9474), .Y(n2944) );
  OAI22X1 U3480 ( .A(n9401), .B(n2881), .C(n11429), .D(n2946), .Y(n2945) );
  AOI22X1 U3481 ( .A(n11475), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[13] ), .D(n2948), .Y(n2946) );
  NAND2X1 U3483 ( .A(n2920), .B(n11478), .Y(n2948) );
  NAND2X1 U3485 ( .A(n2905), .B(n2229), .Y(n2881) );
  NOR2X1 U3486 ( .A(n11376), .B(n11498), .Y(n2879) );
  AOI22X1 U3487 ( .A(n11408), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[13] ), .D(n9441), .Y(n2936) );
  NAND2X1 U3488 ( .A(n2950), .B(n2951), .Y(n8398) );
  AOI22X1 U3489 ( .A(n2952), .B(n2953), .C(n11408), .D(n9373), .Y(n2951) );
  OAI21X1 U3490 ( .A(n9368), .B(n2954), .C(n2955), .Y(n2953) );
  AOI22X1 U3491 ( .A(n2956), .B(n2924), .C(n11394), .D(n9438), .Y(n2955) );
  OAI21X1 U3493 ( .A(n9396), .B(n2926), .C(n2958), .Y(n2957) );
  AOI22X1 U3494 ( .A(n2893), .B(n2959), .C(n11376), .D(n9474), .Y(n2958) );
  OAI22X1 U3495 ( .A(n9401), .B(n2895), .C(n11498), .D(n2960), .Y(n2959) );
  AOI22X1 U3496 ( .A(n11424), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[12] ), .D(n2962), .Y(n2960) );
  NAND2X1 U3498 ( .A(n2920), .B(n11427), .Y(n2962) );
  NAND2X1 U3500 ( .A(n2905), .B(n2250), .Y(n2895) );
  NOR2X1 U3501 ( .A(n11447), .B(n11376), .Y(n2893) );
  AOI22X1 U3502 ( .A(n11476), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[12] ), .D(n2200), .Y(n2950) );
  NAND2X1 U3503 ( .A(n2964), .B(n2965), .Y(n8399) );
  AOI22X1 U3504 ( .A(n2966), .B(n2967), .C(n11476), .D(n9373), .Y(n2965) );
  OAI21X1 U3505 ( .A(n9368), .B(n2968), .C(n2969), .Y(n2967) );
  AOI22X1 U3506 ( .A(n2970), .B(n2938), .C(n11459), .D(n9438), .Y(n2969) );
  OAI21X1 U3508 ( .A(n9396), .B(n2940), .C(n2972), .Y(n2971) );
  AOI22X1 U3509 ( .A(n2909), .B(n2973), .C(n11447), .D(n9474), .Y(n2972) );
  OAI22X1 U3510 ( .A(n9401), .B(n2911), .C(n11376), .D(n2974), .Y(n2973) );
  AOI22X1 U3511 ( .A(n11493), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[11] ), .D(n2976), .Y(n2974) );
  NAND2X1 U3513 ( .A(n2920), .B(n11496), .Y(n2976) );
  NAND2X1 U3515 ( .A(n2905), .B(n2267), .Y(n2911) );
  NOR2X1 U3516 ( .A(n11394), .B(n11447), .Y(n2909) );
  AOI22X1 U3517 ( .A(n11425), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[11] ), .D(n2200), .Y(n2964) );
  NAND2X1 U3518 ( .A(n2978), .B(n2979), .Y(n8400) );
  AOI22X1 U3519 ( .A(n2980), .B(n2981), .C(n11425), .D(n9373), .Y(n2979) );
  OAI21X1 U3520 ( .A(n9368), .B(n2982), .C(n2983), .Y(n2981) );
  AOI22X1 U3521 ( .A(n2984), .B(n2952), .C(n11408), .D(n9438), .Y(n2983) );
  OAI21X1 U3523 ( .A(n9396), .B(n2954), .C(n2986), .Y(n2985) );
  AOI22X1 U3524 ( .A(n2924), .B(n2987), .C(n11394), .D(n9474), .Y(n2986) );
  OAI22X1 U3525 ( .A(n9401), .B(n2926), .C(n11447), .D(n2988), .Y(n2987) );
  AOI22X1 U3526 ( .A(n11371), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[10] ), .D(n2990), .Y(n2988) );
  NAND2X1 U3528 ( .A(n2920), .B(n11374), .Y(n2990) );
  NAND2X1 U3530 ( .A(n2905), .B(n2287), .Y(n2926) );
  NOR2X1 U3531 ( .A(n11459), .B(n11394), .Y(n2924) );
  AOI22X1 U3532 ( .A(n11494), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[10] ), .D(n9443), .Y(n2978) );
  NAND2X1 U3533 ( .A(n2992), .B(n2993), .Y(n8401) );
  AOI22X1 U3534 ( .A(n2994), .B(n2995), .C(n11494), .D(n9374), .Y(n2993) );
  OAI21X1 U3535 ( .A(n9368), .B(n2996), .C(n2997), .Y(n2995) );
  AOI22X1 U3536 ( .A(n2998), .B(n2966), .C(n11476), .D(n9438), .Y(n2997) );
  OAI21X1 U3538 ( .A(n9396), .B(n2968), .C(n3000), .Y(n2999) );
  AOI22X1 U3539 ( .A(n2938), .B(n3001), .C(n11459), .D(n9474), .Y(n3000) );
  OAI22X1 U3540 ( .A(n9401), .B(n2940), .C(n11394), .D(n3002), .Y(n3001) );
  AOI22X1 U3541 ( .A(n11442), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[9] ), .D(n3004), .Y(n3002) );
  NAND2X1 U3543 ( .A(n2920), .B(n11445), .Y(n3004) );
  NAND2X1 U3545 ( .A(n2905), .B(n2301), .Y(n2940) );
  NOR2X1 U3546 ( .A(n11508), .B(n2316), .Y(n2301) );
  NOR2X1 U3547 ( .A(n11408), .B(n11459), .Y(n2938) );
  AOI22X1 U3548 ( .A(n11372), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[9] ), .D(n2200), .Y(n2992) );
  NAND2X1 U3549 ( .A(n3006), .B(n3007), .Y(n8402) );
  AOI22X1 U3550 ( .A(n3008), .B(n3009), .C(n11372), .D(n9374), .Y(n3007) );
  OAI21X1 U3551 ( .A(n9368), .B(n3010), .C(n3011), .Y(n3009) );
  AOI22X1 U3552 ( .A(n3012), .B(n2980), .C(n11425), .D(n9438), .Y(n3011) );
  OAI21X1 U3554 ( .A(n9397), .B(n2982), .C(n3014), .Y(n3013) );
  AOI22X1 U3555 ( .A(n2952), .B(n3015), .C(n11408), .D(n9474), .Y(n3014) );
  OAI22X1 U3556 ( .A(n9401), .B(n2954), .C(n11459), .D(n3016), .Y(n3015) );
  AOI22X1 U3557 ( .A(n11390), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[8] ), .D(n3018), .Y(n3016) );
  NAND2X1 U3559 ( .A(n2920), .B(n11393), .Y(n3018) );
  NAND2X1 U3562 ( .A(n3020), .B(n11461), .Y(n2954) );
  NOR2X1 U3563 ( .A(n11476), .B(n11408), .Y(n2952) );
  AOI22X1 U3564 ( .A(n11443), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[8] ), .D(n9443), .Y(n3006) );
  NAND2X1 U3565 ( .A(n3022), .B(n3023), .Y(n8403) );
  AOI22X1 U3566 ( .A(n3024), .B(n3025), .C(n11443), .D(n9374), .Y(n3023) );
  OAI21X1 U3567 ( .A(n9369), .B(n3026), .C(n3027), .Y(n3025) );
  AOI22X1 U3568 ( .A(n3028), .B(n2994), .C(n11494), .D(n9438), .Y(n3027) );
  OAI21X1 U3570 ( .A(n9397), .B(n2996), .C(n3030), .Y(n3029) );
  AOI22X1 U3571 ( .A(n2966), .B(n3031), .C(n11476), .D(n9474), .Y(n3030) );
  OAI22X1 U3572 ( .A(n9402), .B(n2968), .C(n11408), .D(n3032), .Y(n3031) );
  AOI22X1 U3573 ( .A(n11460), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[7] ), .D(n3034), .Y(n3032) );
  NAND2X1 U3575 ( .A(n3035), .B(n11461), .Y(n3034) );
  NAND2X1 U3578 ( .A(n3020), .B(n11410), .Y(n2968) );
  NOR2X1 U3579 ( .A(n11425), .B(n11476), .Y(n2966) );
  AOI22X1 U3580 ( .A(n11391), .B(n9451), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[7] ), .D(n9443), .Y(n3022) );
  NAND2X1 U3581 ( .A(n3037), .B(n3038), .Y(n8404) );
  AOI22X1 U3582 ( .A(n3039), .B(n3040), .C(n11391), .D(n9374), .Y(n3038) );
  OAI21X1 U3583 ( .A(n9369), .B(n3041), .C(n3042), .Y(n3040) );
  AOI22X1 U3584 ( .A(n3043), .B(n3008), .C(n11372), .D(n9438), .Y(n3042) );
  OAI21X1 U3586 ( .A(n9397), .B(n3010), .C(n3045), .Y(n3044) );
  AOI22X1 U3587 ( .A(n2980), .B(n3046), .C(n11425), .D(n9474), .Y(n3045) );
  OAI22X1 U3588 ( .A(n9402), .B(n2982), .C(n11476), .D(n3047), .Y(n3046) );
  AOI22X1 U3589 ( .A(n11409), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[6] ), .D(n3049), .Y(n3047) );
  NAND2X1 U3591 ( .A(n3035), .B(n11410), .Y(n3049) );
  NAND2X1 U3594 ( .A(n3020), .B(n11478), .Y(n2982) );
  NOR2X1 U3595 ( .A(n11494), .B(n11425), .Y(n2980) );
  AOI22X1 U3596 ( .A(n11462), .B(n9447), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[6] ), .D(n9443), .Y(n3037) );
  NAND2X1 U3597 ( .A(n3051), .B(n3052), .Y(n8405) );
  AOI22X1 U3598 ( .A(n3053), .B(n3054), .C(n11411), .D(n9447), .Y(n3052) );
  OAI21X1 U3599 ( .A(n9369), .B(n3056), .C(n3057), .Y(n3054) );
  AOI22X1 U3600 ( .A(n3058), .B(n3024), .C(n11443), .D(n9438), .Y(n3057) );
  OAI21X1 U3602 ( .A(n9397), .B(n3026), .C(n3060), .Y(n3059) );
  AOI22X1 U3603 ( .A(n2994), .B(n3061), .C(n11494), .D(n9474), .Y(n3060) );
  OAI22X1 U3604 ( .A(n9402), .B(n2996), .C(n11425), .D(n3062), .Y(n3061) );
  AOI22X1 U3605 ( .A(n11477), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[5] ), .D(n3064), .Y(n3062) );
  NAND2X1 U3607 ( .A(n3035), .B(n11478), .Y(n3064) );
  NAND2X1 U3610 ( .A(n3020), .B(n11427), .Y(n2996) );
  NOR2X1 U3611 ( .A(n11372), .B(n11494), .Y(n2994) );
  AOI22X1 U3612 ( .A(n11462), .B(n9374), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[5] ), .D(n9443), .Y(n3051) );
  NAND2X1 U3613 ( .A(n3065), .B(n3066), .Y(n8406) );
  AOI22X1 U3614 ( .A(n3067), .B(n3068), .C(n11479), .D(n9447), .Y(n3066) );
  OAI21X1 U3615 ( .A(n9369), .B(n3070), .C(n3071), .Y(n3068) );
  AOI22X1 U3616 ( .A(n3072), .B(n3039), .C(n11391), .D(n9438), .Y(n3071) );
  OAI21X1 U3618 ( .A(n9397), .B(n3041), .C(n3074), .Y(n3073) );
  AOI22X1 U3619 ( .A(n3008), .B(n3075), .C(n11372), .D(n9474), .Y(n3074) );
  OAI22X1 U3620 ( .A(n9402), .B(n3010), .C(n11494), .D(n3076), .Y(n3075) );
  AOI22X1 U3621 ( .A(n11426), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[4] ), .D(n3078), .Y(n3076) );
  NAND2X1 U3623 ( .A(n3035), .B(n11427), .Y(n3078) );
  NAND2X1 U3626 ( .A(n3020), .B(n11496), .Y(n3010) );
  NOR2X1 U3627 ( .A(n11443), .B(n11372), .Y(n3008) );
  AOI22X1 U3628 ( .A(n11411), .B(n9374), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[4] ), .D(n9443), .Y(n3065) );
  OAI21X1 U3630 ( .A(n9442), .B(n11540), .C(n3079), .Y(n8407) );
  AOI22X1 U3631 ( .A(n3080), .B(n3081), .C(n11428), .D(n9447), .Y(n3079) );
  OAI21X1 U3632 ( .A(n2175), .B(n3083), .C(n3084), .Y(n3080) );
  OAI21X1 U3633 ( .A(n3085), .B(n3086), .C(n3083), .Y(n3084) );
  OAI21X1 U3634 ( .A(n9165), .B(n3070), .C(n3088), .Y(n3086) );
  NAND3X1 U3635 ( .A(n9445), .B(n3089), .C(n3053), .Y(n3088) );
  OAI21X1 U3636 ( .A(n9397), .B(n3056), .C(n3090), .Y(n3089) );
  AOI22X1 U3637 ( .A(n3024), .B(n3091), .C(n11443), .D(n9474), .Y(n3090) );
  OAI22X1 U3638 ( .A(n9402), .B(n3026), .C(n11372), .D(n3092), .Y(n3091) );
  AOI22X1 U3639 ( .A(n11495), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[3] ), .D(n3094), .Y(n3092) );
  NAND2X1 U3641 ( .A(n3035), .B(n11496), .Y(n3094) );
  NAND2X1 U3644 ( .A(n3020), .B(n11374), .Y(n3026) );
  NOR2X1 U3645 ( .A(n11391), .B(n11443), .Y(n3024) );
  NOR2X1 U3646 ( .A(n9369), .B(n3095), .Y(n3085) );
  OAI21X1 U3648 ( .A(n9442), .B(n11538), .C(n3096), .Y(n8408) );
  AOI22X1 U3649 ( .A(n3097), .B(n3098), .C(n11497), .D(n9447), .Y(n3096) );
  OAI21X1 U3650 ( .A(n2175), .B(n3081), .C(n3100), .Y(n3097) );
  OAI21X1 U3651 ( .A(n3101), .B(n3102), .C(n3081), .Y(n3100) );
  OAI21X1 U3652 ( .A(n9165), .B(n3095), .C(n3103), .Y(n3102) );
  NAND3X1 U3653 ( .A(n9445), .B(n3104), .C(n3067), .Y(n3103) );
  OAI21X1 U3654 ( .A(n9397), .B(n3070), .C(n3105), .Y(n3104) );
  AOI22X1 U3655 ( .A(n3039), .B(n3106), .C(n11391), .D(n9474), .Y(n3105) );
  OAI22X1 U3656 ( .A(n9402), .B(n3041), .C(n11443), .D(n3107), .Y(n3106) );
  AOI22X1 U3657 ( .A(n11373), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[2] ), .D(n3109), .Y(n3107) );
  NAND2X1 U3659 ( .A(n3035), .B(n11374), .Y(n3109) );
  NAND2X1 U3662 ( .A(n3020), .B(n11445), .Y(n3041) );
  NOR2X1 U3663 ( .A(n11462), .B(n11391), .Y(n3039) );
  NOR2X1 U3664 ( .A(n9369), .B(n3083), .Y(n3101) );
  OAI21X1 U3667 ( .A(n9442), .B(n11536), .C(n3110), .Y(n8409) );
  AOI22X1 U3668 ( .A(n3111), .B(n3112), .C(n11375), .D(n9447), .Y(n3110) );
  OAI22X1 U3670 ( .A(n2175), .B(n3098), .C(n11497), .D(n3114), .Y(n3111) );
  AOI22X1 U3671 ( .A(n3115), .B(n3081), .C(n11428), .D(n2242), .Y(n3114) );
  NOR2X1 U3672 ( .A(n9444), .B(n11516), .Y(n2242) );
  OAI21X1 U3674 ( .A(n9165), .B(n3083), .C(n3116), .Y(n3115) );
  NAND3X1 U3675 ( .A(n3117), .B(n3083), .C(n9445), .Y(n3116) );
  OAI21X1 U3676 ( .A(n9393), .B(n3095), .C(n3118), .Y(n3117) );
  AOI22X1 U3677 ( .A(n3053), .B(n3119), .C(n11462), .D(n9474), .Y(n3118) );
  OAI22X1 U3678 ( .A(n9402), .B(n3056), .C(n11391), .D(n3120), .Y(n3119) );
  AOI22X1 U3679 ( .A(n11444), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[1] ), .D(n3122), .Y(n3120) );
  NAND2X1 U3681 ( .A(n3035), .B(n11445), .Y(n3122) );
  NAND2X1 U3684 ( .A(n3020), .B(n11393), .Y(n3056) );
  NOR2X1 U3687 ( .A(\U_1/U_0/U_1/U_8/address[6] ), .B(
        \U_1/U_0/U_1/U_8/address[7] ), .Y(n2429) );
  NOR2X1 U3688 ( .A(n11411), .B(n11462), .Y(n3053) );
  OAI21X1 U3693 ( .A(n9442), .B(n11534), .C(n3123), .Y(n8410) );
  AOI22X1 U3694 ( .A(n3124), .B(n3125), .C(n11446), .D(n9447), .Y(n3123) );
  NOR2X1 U3695 ( .A(n9444), .B(n11513), .Y(n2170) );
  NAND2X1 U3699 ( .A(n11506), .B(n2287), .Y(n3125) );
  NOR2X1 U3700 ( .A(n2302), .B(n11508), .Y(n2287) );
  NAND3X1 U3701 ( .A(n11503), .B(n11504), .C(\U_1/U_0/U_1/U_8/address[0] ), 
        .Y(n2302) );
  OAI22X1 U3702 ( .A(n3130), .B(n3131), .C(n2175), .D(n3112), .Y(n3124) );
  NAND2X1 U3703 ( .A(n9446), .B(\U_1/U_0/U_1/RCV_DATA [6]), .Y(n2175) );
  OAI21X1 U3704 ( .A(\U_1/U_0/U_1/RCV_DATA [5]), .B(n3098), .C(n9446), .Y(
        n3131) );
  NOR2X1 U3705 ( .A(n3132), .B(n9443), .Y(n2177) );
  OAI21X1 U3706 ( .A(n11497), .B(n3133), .C(n3112), .Y(n3130) );
  NAND2X1 U3707 ( .A(n11506), .B(n2267), .Y(n3112) );
  NOR2X1 U3708 ( .A(n2286), .B(n11508), .Y(n2267) );
  NAND3X1 U3709 ( .A(n11433), .B(n11504), .C(\U_1/U_0/U_1/U_8/address[1] ), 
        .Y(n2286) );
  AOI22X1 U3710 ( .A(n11428), .B(n11518), .C(n3135), .D(n3136), .Y(n3133) );
  AOI21X1 U3711 ( .A(n3067), .B(n3137), .C(n11428), .Y(n3136) );
  OAI22X1 U3712 ( .A(n9398), .B(n3070), .C(n11462), .D(n3138), .Y(n3137) );
  AOI22X1 U3713 ( .A(n11392), .B(n9479), .C(
        \U_1/U_0/U_1/U_8/currentPlainKey[0] ), .D(n3140), .Y(n3138) );
  NAND2X1 U3715 ( .A(n3035), .B(n11393), .Y(n3140) );
  NAND3X1 U3717 ( .A(n11503), .B(n11504), .C(n11433), .Y(n2316) );
  NOR2X1 U3719 ( .A(\U_1/U_0/U_1/U_8/address[4] ), .B(
        \U_1/U_0/U_1/U_8/address[5] ), .Y(n3019) );
  NAND2X1 U3721 ( .A(n11506), .B(n2445), .Y(n3070) );
  NOR2X1 U3722 ( .A(n2197), .B(n11508), .Y(n2445) );
  NAND3X1 U3723 ( .A(\U_1/U_0/U_1/U_8/address[1] ), .B(
        \U_1/U_0/U_1/U_8/address[0] ), .C(\U_1/U_0/U_1/U_8/address[2] ), .Y(
        n2197) );
  NOR2X1 U3725 ( .A(n11479), .B(n11411), .Y(n3067) );
  AOI22X1 U3726 ( .A(n11411), .B(n9474), .C(n11479), .D(
        \U_1/U_0/U_1/RCV_DATA [3]), .Y(n3135) );
  NAND2X1 U3728 ( .A(n11506), .B(n2215), .Y(n3083) );
  NOR2X1 U3729 ( .A(n2232), .B(n11508), .Y(n2215) );
  NAND3X1 U3730 ( .A(\U_1/U_0/U_1/U_8/address[0] ), .B(n11503), .C(
        \U_1/U_0/U_1/U_8/address[2] ), .Y(n2232) );
  NAND2X1 U3732 ( .A(n11506), .B(n2192), .Y(n3095) );
  NOR2X1 U3733 ( .A(n2212), .B(n11508), .Y(n2192) );
  NAND3X1 U3734 ( .A(\U_1/U_0/U_1/U_8/address[1] ), .B(n11433), .C(
        \U_1/U_0/U_1/U_8/address[2] ), .Y(n2212) );
  NAND2X1 U3737 ( .A(n11506), .B(n2229), .Y(n3081) );
  NOR2X1 U3738 ( .A(n2247), .B(n11508), .Y(n2229) );
  NAND3X1 U3739 ( .A(n11433), .B(n11503), .C(\U_1/U_0/U_1/U_8/address[2] ), 
        .Y(n2247) );
  NAND2X1 U3741 ( .A(n11506), .B(n2250), .Y(n3098) );
  NOR2X1 U3742 ( .A(n2266), .B(n11508), .Y(n2250) );
  NAND3X1 U3744 ( .A(\U_1/U_0/U_1/U_8/address[0] ), .B(n11504), .C(
        \U_1/U_0/U_1/U_8/address[1] ), .Y(n2266) );
  NAND3X1 U3746 ( .A(\U_1/U_0/U_1/U_8/address[6] ), .B(n2319), .C(
        \U_1/U_0/U_1/U_8/address[7] ), .Y(n3141) );
  NOR2X1 U3747 ( .A(n11510), .B(n11511), .Y(n2319) );
  NAND2X1 U3752 ( .A(n3142), .B(n11354), .Y(n2200) );
  OAI21X1 U3753 ( .A(n9245), .B(n11532), .C(n3146), .Y(n8411) );
  NAND2X1 U3754 ( .A(\U_1/U_0/U_1/U_8/N1799 ), .B(n3147), .Y(n3146) );
  OAI21X1 U3755 ( .A(n9245), .B(n11531), .C(n3149), .Y(n8412) );
  NAND2X1 U3756 ( .A(\U_1/U_0/U_1/U_8/N1798 ), .B(n3147), .Y(n3149) );
  OAI21X1 U3757 ( .A(n9245), .B(n11530), .C(n3151), .Y(n8413) );
  NAND2X1 U3758 ( .A(\U_1/U_0/U_1/U_8/N1797 ), .B(n3147), .Y(n3151) );
  OAI21X1 U3760 ( .A(n9245), .B(n11529), .C(n3153), .Y(n8414) );
  NAND2X1 U3761 ( .A(\U_1/U_0/U_1/U_8/N1796 ), .B(n3147), .Y(n3153) );
  OAI21X1 U3763 ( .A(n9245), .B(n11528), .C(n3155), .Y(n8415) );
  NAND2X1 U3764 ( .A(\U_1/U_0/U_1/U_8/N1795 ), .B(n3147), .Y(n3155) );
  OAI21X1 U3765 ( .A(n9245), .B(n11527), .C(n3157), .Y(n8416) );
  NAND2X1 U3766 ( .A(\U_1/U_0/U_1/U_8/N1794 ), .B(n3147), .Y(n3157) );
  OAI21X1 U3767 ( .A(n9245), .B(n11526), .C(n3159), .Y(n8417) );
  NAND2X1 U3768 ( .A(\U_1/U_0/U_1/U_8/N1793 ), .B(n3147), .Y(n3159) );
  OAI21X1 U3770 ( .A(n9245), .B(n11525), .C(n3161), .Y(n8418) );
  NAND2X1 U3771 ( .A(\U_1/U_0/U_1/U_8/N1792 ), .B(n3147), .Y(n3161) );
  OAI22X1 U3774 ( .A(n9244), .B(n11524), .C(n11522), .D(n3164), .Y(n8419) );
  OAI22X1 U3776 ( .A(n9244), .B(n11522), .C(n11521), .D(n3164), .Y(n8420) );
  OAI22X1 U3778 ( .A(n9244), .B(n11521), .C(n11519), .D(n3164), .Y(n8421) );
  OAI22X1 U3780 ( .A(n9244), .B(n11519), .C(n11517), .D(n3164), .Y(n8422) );
  OAI22X1 U3782 ( .A(n9244), .B(n11517), .C(n11515), .D(n3164), .Y(n8423) );
  OAI22X1 U3784 ( .A(n9244), .B(n11515), .C(n11514), .D(n3164), .Y(n8424) );
  OAI22X1 U3786 ( .A(n9244), .B(n11514), .C(n11512), .D(n3164), .Y(n8425) );
  OAI22X1 U3788 ( .A(n9244), .B(n11512), .C(n3164), .D(n11319), .Y(n8426) );
  OAI21X1 U3790 ( .A(n3167), .B(n11433), .C(n3168), .Y(n8427) );
  OAI21X1 U3792 ( .A(n3167), .B(n11503), .C(n3168), .Y(n8428) );
  OAI21X1 U3794 ( .A(n3167), .B(n11504), .C(n3168), .Y(n8429) );
  OAI21X1 U3796 ( .A(n10539), .B(n11358), .C(n3171), .Y(n8430) );
  AOI21X1 U3797 ( .A(\U_1/U_0/U_1/U_8/address[3] ), .B(n10539), .C(n10540), 
        .Y(n3171) );
  OAI21X1 U3798 ( .A(n10539), .B(n11355), .C(n3174), .Y(n8431) );
  AOI21X1 U3799 ( .A(\U_1/U_0/U_1/U_8/address[4] ), .B(n10539), .C(n10540), 
        .Y(n3174) );
  OAI21X1 U3800 ( .A(n10539), .B(n11356), .C(n3176), .Y(n8432) );
  AOI21X1 U3801 ( .A(\U_1/U_0/U_1/U_8/address[5] ), .B(n10539), .C(n10540), 
        .Y(n3176) );
  OAI21X1 U3804 ( .A(n3167), .B(n11505), .C(n3168), .Y(n8433) );
  OAI21X1 U3806 ( .A(n3167), .B(n11507), .C(n3168), .Y(n8434) );
  NAND2X1 U3807 ( .A(\U_1/U_0/U_1/U_8/keyCount[3] ), .B(n3167), .Y(n3168) );
  NOR2X1 U3809 ( .A(n3179), .B(n3180), .Y(n3167) );
  NAND3X1 U3810 ( .A(n3181), .B(n11352), .C(n7749), .Y(n3180) );
  NOR2X1 U3811 ( .A(n3162), .B(RST), .Y(n7749) );
  NAND3X1 U3812 ( .A(n3183), .B(n11354), .C(n3184), .Y(n3179) );
  OAI21X1 U3813 ( .A(n3185), .B(n3186), .C(n3187), .Y(n8435) );
  NAND2X1 U3814 ( .A(\U_1/U_0/U_1/U_8/keyCount[3] ), .B(n3188), .Y(n3187) );
  OAI21X1 U3815 ( .A(\U_1/U_0/U_1/U_8/keyCount[2] ), .B(n3132), .C(n3189), .Y(
        n3188) );
  OAI21X1 U3816 ( .A(n3189), .B(n11356), .C(n3190), .Y(n8436) );
  NAND3X1 U3817 ( .A(\U_1/U_0/U_1/U_8/keyCount[0] ), .B(n11356), .C(n3191), 
        .Y(n3190) );
  NOR2X1 U3818 ( .A(n11355), .B(n3186), .Y(n3191) );
  AOI21X1 U3820 ( .A(n11355), .B(n11342), .C(n3193), .Y(n3189) );
  OAI21X1 U3821 ( .A(n10053), .B(n11355), .C(n3195), .Y(n8437) );
  NAND3X1 U3822 ( .A(\U_1/U_0/U_1/U_8/keyCount[0] ), .B(n11355), .C(n10052), 
        .Y(n3195) );
  OAI21X1 U3826 ( .A(\U_1/U_0/U_1/U_8/keyCount[0] ), .B(n3132), .C(n3142), .Y(
        n3193) );
  OAI22X1 U3827 ( .A(n3142), .B(n11358), .C(\U_1/U_0/U_1/U_8/keyCount[0] ), 
        .D(n3186), .Y(n8438) );
  NAND2X1 U3828 ( .A(n11342), .B(n3142), .Y(n3186) );
  NOR2X1 U3830 ( .A(n3198), .B(n3199), .Y(n3144) );
  NAND3X1 U3831 ( .A(n3200), .B(n3184), .C(n11352), .Y(n3199) );
  NAND3X1 U3832 ( .A(n3183), .B(n9518), .C(n3201), .Y(n3198) );
  NAND3X1 U3833 ( .A(n3201), .B(n3132), .C(n3202), .Y(n8439) );
  AOI21X1 U3834 ( .A(\U_1/U_0/U_1/U_8/state[1] ), .B(n3203), .C(n11348), .Y(
        n3202) );
  OAI21X1 U3835 ( .A(n11340), .B(n11359), .C(n3197), .Y(n8440) );
  OAI21X1 U3837 ( .A(n3207), .B(n3208), .C(n3209), .Y(n3203) );
  OAI21X1 U3838 ( .A(n11361), .B(\U_1/U_0/U_1/U_8/keyCount[3] ), .C(n11350), 
        .Y(n3208) );
  NAND2X1 U3840 ( .A(n11362), .B(n11341), .Y(n3207) );
  NAND3X1 U3841 ( .A(n3215), .B(n3216), .C(n3217), .Y(n8441) );
  AOI21X1 U3842 ( .A(n11342), .B(n3185), .C(n3218), .Y(n3217) );
  OAI21X1 U3843 ( .A(n11349), .B(n3209), .C(n3220), .Y(n3218) );
  OAI21X1 U3844 ( .A(n11351), .B(n11348), .C(\U_1/RBUF_FULL ), .Y(n3220) );
  NAND3X1 U3846 ( .A(n11362), .B(n11341), .C(n11350), .Y(n3216) );
  NOR2X1 U3849 ( .A(n3222), .B(n3223), .Y(n3215) );
  OAI21X1 U3851 ( .A(\U_1/RBUF_FULL ), .B(n11354), .C(n11347), .Y(n3225) );
  OAI22X1 U3853 ( .A(n3209), .B(n11357), .C(n3185), .D(n3132), .Y(n3227) );
  NAND3X1 U3854 ( .A(\U_1/U_0/U_1/U_8/keyCount[2] ), .B(
        \U_1/U_0/U_1/U_8/keyCount[1] ), .C(n3229), .Y(n3185) );
  NOR2X1 U3855 ( .A(\U_1/U_0/U_1/U_8/keyCount[3] ), .B(n11358), .Y(n3229) );
  OAI21X1 U3857 ( .A(\U_1/U_0/U_1/U_8/state[3] ), .B(n3230), .C(n3231), .Y(
        n3209) );
  NAND3X1 U3859 ( .A(n11352), .B(n3200), .C(n3232), .Y(n3224) );
  OAI21X1 U3860 ( .A(\U_1/U_0/U_1/OE ), .B(\U_1/U_0/U_1/SBE ), .C(n11350), .Y(
        n3232) );
  OAI21X1 U3862 ( .A(n11320), .B(n3234), .C(n3235), .Y(n8443) );
  NAND3X1 U3863 ( .A(n3236), .B(n3237), .C(\U_1/U_0/U_1/SET_RBUF_FULL ), .Y(
        n3235) );
  XNOR2X1 U3864 ( .A(n11322), .B(\U_1/U_0/U_1/U_2/nextState[0] ), .Y(n3234) );
  OAI21X1 U3865 ( .A(n3239), .B(n11329), .C(n3237), .Y(n8444) );
  OAI21X1 U3866 ( .A(n3239), .B(n11330), .C(n3237), .Y(n8445) );
  NAND2X1 U3867 ( .A(n3236), .B(n3242), .Y(n3239) );
  OAI21X1 U3868 ( .A(n11322), .B(n3243), .C(n3244), .Y(n8446) );
  NAND3X1 U3869 ( .A(n3236), .B(n3237), .C(\U_1/U_0/U_1/RBUF_LOAD ), .Y(n3244)
         );
  NAND2X1 U3870 ( .A(\U_1/U_0/U_1/U_2/nextState[2] ), .B(n11312), .Y(n3243) );
  OAI21X1 U3871 ( .A(n11328), .B(n3247), .C(n3248), .Y(n8447) );
  NAND2X1 U3872 ( .A(n3236), .B(n3237), .Y(n3247) );
  OAI21X1 U3873 ( .A(n11339), .B(n3250), .C(n3242), .Y(n8448) );
  NAND3X1 U3874 ( .A(n11312), .B(n11320), .C(\U_1/U_0/U_1/U_2/nextState[1] ), 
        .Y(n3242) );
  NAND2X1 U3875 ( .A(n3248), .B(n3236), .Y(n3250) );
  NAND2X1 U3876 ( .A(\U_1/U_0/U_1/U_2/nextState[2] ), .B(n11322), .Y(n3248) );
  OAI21X1 U3877 ( .A(n3251), .B(n11323), .C(n3237), .Y(n8449) );
  NAND3X1 U3878 ( .A(n11322), .B(n11320), .C(\U_1/U_0/U_1/U_2/nextState[0] ), 
        .Y(n3237) );
  NAND3X1 U3880 ( .A(n11322), .B(n11320), .C(n11312), .Y(n3236) );
  OAI22X1 U3884 ( .A(n9244), .B(n11319), .C(n3164), .D(n11318), .Y(n8450) );
  OAI22X1 U3885 ( .A(n9244), .B(n11318), .C(n3164), .D(n10543), .Y(n8451) );
  OAI21X1 U3888 ( .A(n3255), .B(n3256), .C(n3257), .Y(n3164) );
  NOR2X1 U3889 ( .A(\U_1/U_0/U_1/U_7/state[7] ), .B(\U_1/U_0/U_1/U_7/state[0] ), .Y(n3257) );
  OAI21X1 U3890 ( .A(n11335), .B(n3259), .C(n3260), .Y(n3256) );
  NAND3X1 U3891 ( .A(\U_1/U_0/U_1/U_7/state[6] ), .B(
        \U_1/U_0/U_1/U_7/state[1] ), .C(n3261), .Y(n3260) );
  AOI21X1 U3892 ( .A(n3262), .B(n3263), .C(\U_1/U_0/U_1/U_7/state[3] ), .Y(
        n3261) );
  NAND3X1 U3893 ( .A(n11335), .B(n11317), .C(\U_1/U_0/U_1/U_7/state[4] ), .Y(
        n3263) );
  NAND3X1 U3895 ( .A(\U_1/U_0/U_1/U_7/state[2] ), .B(n11338), .C(
        \U_1/U_0/U_1/U_7/state[5] ), .Y(n3262) );
  NAND2X1 U3896 ( .A(\U_1/U_0/U_1/U_7/state[4] ), .B(n3266), .Y(n3259) );
  AOI21X1 U3897 ( .A(n11315), .B(n11335), .C(n3268), .Y(n3255) );
  NAND2X1 U3898 ( .A(n3269), .B(n11338), .Y(n3268) );
  OAI21X1 U3900 ( .A(n3270), .B(n3271), .C(\U_1/U_0/U_1/U_7/state[2] ), .Y(
        n3269) );
  NAND2X1 U3901 ( .A(\U_1/U_0/U_1/U_7/state[3] ), .B(n11333), .Y(n3271) );
  OAI21X1 U3906 ( .A(\U_1/U_0/U_1/U_7/state[6] ), .B(n3273), .C(n3274), .Y(
        n3266) );
  NAND3X1 U3907 ( .A(\U_1/U_0/U_1/U_7/state[3] ), .B(
        \U_1/U_0/U_1/U_7/state[6] ), .C(n3275), .Y(n3274) );
  NOR2X1 U3908 ( .A(\U_1/U_0/U_1/U_7/state[5] ), .B(\U_1/U_0/U_1/U_7/state[1] ), .Y(n3275) );
  AOI22X1 U3909 ( .A(n3276), .B(\U_1/U_0/U_1/U_7/state[1] ), .C(n3277), .D(
        \U_1/U_0/U_1/U_7/state[5] ), .Y(n3273) );
  XNOR2X1 U3910 ( .A(\U_1/U_0/U_1/U_7/state[1] ), .B(
        \U_1/U_0/U_1/U_7/state[3] ), .Y(n3277) );
  NOR2X1 U3911 ( .A(\U_1/U_0/U_1/U_7/state[5] ), .B(\U_1/U_0/U_1/U_7/state[3] ), .Y(n3276) );
  OAI21X1 U3912 ( .A(n11331), .B(n3279), .C(n3280), .Y(n8452) );
  NAND2X1 U3913 ( .A(\U_1/U_0/U_1/U_7/N26 ), .B(n3281), .Y(n3280) );
  OAI21X1 U3915 ( .A(n3279), .B(n11332), .C(n3283), .Y(n8453) );
  NAND2X1 U3916 ( .A(\U_1/U_0/U_1/U_7/N27 ), .B(n3281), .Y(n3283) );
  OAI21X1 U3917 ( .A(n11334), .B(n3279), .C(n3285), .Y(n8454) );
  NAND2X1 U3918 ( .A(\U_1/U_0/U_1/U_7/N28 ), .B(n3281), .Y(n3285) );
  OAI21X1 U3919 ( .A(n11336), .B(n3279), .C(n3287), .Y(n8455) );
  NAND2X1 U3920 ( .A(\U_1/U_0/U_1/U_7/N29 ), .B(n3281), .Y(n3287) );
  OAI21X1 U3921 ( .A(n3279), .B(n11337), .C(n3289), .Y(n8456) );
  NAND2X1 U3922 ( .A(\U_1/U_0/U_1/U_7/N30 ), .B(n3281), .Y(n3289) );
  OAI21X1 U3924 ( .A(n11316), .B(n3279), .C(n3291), .Y(n8457) );
  NAND2X1 U3925 ( .A(\U_1/U_0/U_1/U_7/N31 ), .B(n3281), .Y(n3291) );
  OAI21X1 U3927 ( .A(n11314), .B(n3279), .C(n3293), .Y(n8458) );
  NAND2X1 U3928 ( .A(\U_1/U_0/U_1/U_7/N32 ), .B(n3281), .Y(n3293) );
  OAI21X1 U3930 ( .A(n3279), .B(n11313), .C(n3295), .Y(n8459) );
  NAND2X1 U3931 ( .A(\U_1/U_0/U_1/U_7/N33 ), .B(n3281), .Y(n3295) );
  NAND2X1 U3934 ( .A(n11330), .B(n3296), .Y(n3279) );
  NAND3X1 U3936 ( .A(\U_1/U_0/U_1/U_7/nextState[6] ), .B(
        \U_1/U_0/U_1/U_7/nextState[5] ), .C(n3299), .Y(n3298) );
  NOR2X1 U3937 ( .A(n11334), .B(n11336), .Y(n3299) );
  NAND3X1 U3940 ( .A(\U_1/U_0/U_1/U_7/nextState[0] ), .B(n11332), .C(n3300), 
        .Y(n3297) );
  NOR2X1 U3941 ( .A(\U_1/U_0/U_1/U_7/nextState[7] ), .B(
        \U_1/U_0/U_1/U_7/nextState[4] ), .Y(n3300) );
  OAI22X1 U3944 ( .A(n10868), .B(n11311), .C(n10879), .D(n3303), .Y(n8460) );
  NAND3X1 U3946 ( .A(\U_0/U_3/U_0/N59 ), .B(n10875), .C(n3305), .Y(n3303) );
  NOR2X1 U3947 ( .A(n3306), .B(n3307), .Y(n3305) );
  AOI22X1 U3949 ( .A(\U_0/U_3/send_data [7]), .B(n10889), .C(n3310), .D(
        \U_0/U_3/U_2/present_val [7]), .Y(n3308) );
  OAI21X1 U3950 ( .A(n11290), .B(n3312), .C(n3313), .Y(n8462) );
  AOI22X1 U3951 ( .A(n9243), .B(\U_0/U_3/U_2/present_val [7]), .C(
        \U_0/U_3/U_2/present_val [6]), .D(n3310), .Y(n3313) );
  OAI21X1 U3953 ( .A(n11292), .B(n3312), .C(n3316), .Y(n8463) );
  AOI22X1 U3954 ( .A(\U_0/U_3/U_2/present_val [6]), .B(n9243), .C(
        \U_0/U_3/U_2/present_val [5]), .D(n3310), .Y(n3316) );
  OAI21X1 U3956 ( .A(n11294), .B(n3312), .C(n3318), .Y(n8464) );
  AOI22X1 U3957 ( .A(\U_0/U_3/U_2/present_val [5]), .B(n9243), .C(
        \U_0/U_3/U_2/present_val [4]), .D(n3310), .Y(n3318) );
  OAI21X1 U3959 ( .A(n11296), .B(n3312), .C(n3320), .Y(n8465) );
  AOI22X1 U3960 ( .A(\U_0/U_3/U_2/present_val [4]), .B(n9243), .C(
        \U_0/U_3/U_2/present_val [3]), .D(n3310), .Y(n3320) );
  OAI21X1 U3962 ( .A(n11298), .B(n3312), .C(n3322), .Y(n8466) );
  AOI22X1 U3963 ( .A(\U_0/U_3/U_2/present_val [3]), .B(n9243), .C(
        \U_0/U_3/U_2/present_val [2]), .D(n3310), .Y(n3322) );
  OAI21X1 U3965 ( .A(n11300), .B(n3312), .C(n3324), .Y(n8467) );
  AOI22X1 U3966 ( .A(\U_0/U_3/U_2/present_val [2]), .B(n9243), .C(
        \U_0/U_3/U_2/present_val [1]), .D(n3310), .Y(n3324) );
  OAI21X1 U3968 ( .A(n11302), .B(n3312), .C(n3326), .Y(n8468) );
  AOI22X1 U3969 ( .A(\U_0/U_3/U_2/present_val [1]), .B(n9243), .C(
        \U_0/U_3/d_encode ), .D(n3310), .Y(n3326) );
  OAI21X1 U3971 ( .A(n10889), .B(n11308), .C(n3328), .Y(n8469) );
  NAND3X1 U3972 ( .A(\U_0/U_3/U_2/count[1] ), .B(\U_0/U_3/U_2/count[0] ), .C(
        n9243), .Y(n3328) );
  OAI21X1 U3973 ( .A(n10872), .B(n3330), .C(n3331), .Y(n8470) );
  OAI21X1 U3974 ( .A(n3310), .B(n11309), .C(\U_0/U_3/U_2/count[1] ), .Y(n3331)
         );
  NAND2X1 U3975 ( .A(\U_0/U_3/U_2/count[0] ), .B(n11307), .Y(n3330) );
  AOI22X1 U3978 ( .A(\U_0/U_3/U_2/count[0] ), .B(n3310), .C(n11309), .D(n9243), 
        .Y(n3334) );
  NOR2X1 U3979 ( .A(n10889), .B(n3310), .Y(n3314) );
  AOI21X1 U3981 ( .A(\U_0/U_3/U_0/N59 ), .B(n7754), .C(n10889), .Y(n3310) );
  NAND3X1 U3983 ( .A(\U_0/U_3/U_2/count[0] ), .B(n7754), .C(n3335), .Y(n3312)
         );
  NOR2X1 U3984 ( .A(n11307), .B(n11308), .Y(n3335) );
  NOR2X1 U3987 ( .A(n3336), .B(n3337), .Y(n7754) );
  NAND3X1 U3988 ( .A(\U_0/U_3/U_4/count[3] ), .B(host_is_sending), .C(
        \U_0/U_3/U_4/state ), .Y(n3337) );
  OAI22X1 U3989 ( .A(n11218), .B(n9242), .C(n3340), .D(n9241), .Y(n8472) );
  XNOR2X1 U3990 ( .A(n3342), .B(n11231), .Y(n3340) );
  OAI22X1 U3992 ( .A(n11229), .B(n9241), .C(n11230), .D(n9242), .Y(n8473) );
  OAI22X1 U3994 ( .A(n11227), .B(n9241), .C(n11228), .D(n9242), .Y(n8474) );
  OAI22X1 U3996 ( .A(n11225), .B(n9241), .C(n11226), .D(n9242), .Y(n8475) );
  OAI22X1 U3998 ( .A(n11223), .B(n9241), .C(n11224), .D(n9242), .Y(n8476) );
  OAI22X1 U3999 ( .A(n11221), .B(n9241), .C(n11222), .D(n9242), .Y(n8477) );
  OAI22X1 U4001 ( .A(n11220), .B(n9242), .C(n3355), .D(n9241), .Y(n8478) );
  XNOR2X1 U4002 ( .A(\U_0/U_3/TX_CRC [1]), .B(n3356), .Y(n3355) );
  OAI22X1 U4004 ( .A(n11233), .B(n9242), .C(n3358), .D(n9241), .Y(n8479) );
  XOR2X1 U4005 ( .A(n3359), .B(n3360), .Y(n3358) );
  XNOR2X1 U4006 ( .A(\U_0/U_3/TX_CRC [0]), .B(n3356), .Y(n3359) );
  OAI22X1 U4007 ( .A(n11231), .B(n9242), .C(n3361), .D(n9241), .Y(n8480) );
  OAI22X1 U4009 ( .A(n11229), .B(n9242), .C(n3362), .D(n3341), .Y(n8481) );
  XNOR2X1 U4010 ( .A(n3363), .B(n3364), .Y(n3362) );
  OAI22X1 U4012 ( .A(n11227), .B(n9242), .C(n3365), .D(n3341), .Y(n8482) );
  OAI22X1 U4014 ( .A(n11225), .B(n9242), .C(n3366), .D(n3341), .Y(n8483) );
  XNOR2X1 U4015 ( .A(n3367), .B(n3368), .Y(n3366) );
  OAI22X1 U4017 ( .A(n11223), .B(n9242), .C(n3369), .D(n3341), .Y(n8484) );
  OAI22X1 U4019 ( .A(n11221), .B(n9242), .C(n3370), .D(n3341), .Y(n8485) );
  XOR2X1 U4020 ( .A(n3371), .B(n3372), .Y(n3370) );
  OAI22X1 U4022 ( .A(n11219), .B(n9242), .C(n3374), .D(n3341), .Y(n8486) );
  XNOR2X1 U4023 ( .A(n3375), .B(n3361), .Y(n3374) );
  XNOR2X1 U4024 ( .A(n3356), .B(n3376), .Y(n3375) );
  OAI22X1 U4026 ( .A(n11232), .B(n9242), .C(n3342), .D(n3341), .Y(n8487) );
  XOR2X1 U4027 ( .A(n3378), .B(n3379), .Y(n3342) );
  XOR2X1 U4028 ( .A(n3356), .B(n3372), .Y(n3379) );
  XNOR2X1 U4029 ( .A(n11233), .B(\U_0/PROCESSED_DATA [0]), .Y(n3372) );
  XOR2X1 U4031 ( .A(\U_0/U_3/TX_CRC [15]), .B(\U_0/PROCESSED_DATA [7]), .Y(
        n3356) );
  XNOR2X1 U4032 ( .A(n11209), .B(n3376), .Y(n3378) );
  XOR2X1 U4033 ( .A(n3369), .B(n3365), .Y(n3376) );
  XNOR2X1 U4034 ( .A(n3364), .B(n3368), .Y(n3365) );
  XNOR2X1 U4035 ( .A(n11224), .B(\U_0/PROCESSED_DATA [3]), .Y(n3368) );
  XNOR2X1 U4037 ( .A(\U_0/U_3/TX_CRC [12]), .B(n11213), .Y(n3364) );
  XOR2X1 U4039 ( .A(n3371), .B(n3367), .Y(n3369) );
  XOR2X1 U4040 ( .A(\U_0/U_3/TX_CRC [10]), .B(\U_0/PROCESSED_DATA [2]), .Y(
        n3367) );
  XNOR2X1 U4041 ( .A(\U_0/U_3/TX_CRC [9]), .B(\U_0/PROCESSED_DATA [1]), .Y(
        n3371) );
  XNOR2X1 U4043 ( .A(n3360), .B(n3363), .Y(n3361) );
  XOR2X1 U4044 ( .A(\U_0/U_3/TX_CRC [13]), .B(\U_0/PROCESSED_DATA [5]), .Y(
        n3363) );
  XNOR2X1 U4045 ( .A(\U_0/U_3/TX_CRC [14]), .B(n11210), .Y(n3360) );
  NAND3X1 U4048 ( .A(n3384), .B(n11114), .C(n3386), .Y(n3341) );
  NOR2X1 U4049 ( .A(n3387), .B(n11094), .Y(n3386) );
  AOI22X1 U4052 ( .A(\U_0/PROCESSED_DATA [6]), .B(n9239), .C(n10051), .D(
        \U_0/U_3/U_3/flop_data [6]), .Y(n3389) );
  AOI22X1 U4054 ( .A(\U_0/PROCESSED_DATA [5]), .B(n9239), .C(n10051), .D(
        \U_0/U_3/U_3/flop_data [5]), .Y(n3390) );
  AOI22X1 U4056 ( .A(\U_0/PROCESSED_DATA [4]), .B(n9239), .C(n10051), .D(
        \U_0/U_3/U_3/flop_data [4]), .Y(n3391) );
  AOI22X1 U4058 ( .A(\U_0/PROCESSED_DATA [3]), .B(n9239), .C(n10051), .D(
        \U_0/U_3/U_3/flop_data [3]), .Y(n3392) );
  AOI22X1 U4060 ( .A(\U_0/PROCESSED_DATA [2]), .B(n9239), .C(n10051), .D(
        \U_0/U_3/U_3/flop_data [2]), .Y(n3393) );
  AOI22X1 U4062 ( .A(\U_0/PROCESSED_DATA [1]), .B(n9239), .C(n10051), .D(
        \U_0/U_3/U_3/flop_data [1]), .Y(n3394) );
  AOI22X1 U4064 ( .A(\U_0/PROCESSED_DATA [0]), .B(n9239), .C(n10051), .D(
        \U_0/U_3/U_3/flop_data [0]), .Y(n3395) );
  NOR2X1 U4066 ( .A(n3396), .B(n3397), .Y(n776) );
  NAND3X1 U4067 ( .A(n10900), .B(n518), .C(n477), .Y(n3397) );
  NAND3X1 U4069 ( .A(n10898), .B(n9534), .C(n519), .Y(n3396) );
  OAI21X1 U4071 ( .A(n9335), .B(n3402), .C(n3403), .Y(n8495) );
  AOI22X1 U4072 ( .A(\U_0/U_3/U_3/N90 ), .B(n3404), .C(\U_0/U_3/U_3/N65 ), .D(
        n3405), .Y(n3403) );
  OAI21X1 U4073 ( .A(n11115), .B(n3402), .C(n3407), .Y(n8496) );
  AOI22X1 U4074 ( .A(\U_0/U_3/U_3/N89 ), .B(n3404), .C(\U_0/U_3/U_3/N64 ), .D(
        n3405), .Y(n3407) );
  OAI21X1 U4075 ( .A(n11120), .B(n3402), .C(n3409), .Y(n8497) );
  AOI22X1 U4076 ( .A(\U_0/U_3/U_3/N88 ), .B(n3404), .C(\U_0/U_3/U_3/N63 ), .D(
        n3405), .Y(n3409) );
  OAI21X1 U4077 ( .A(n11119), .B(n3402), .C(n3411), .Y(n8498) );
  AOI22X1 U4078 ( .A(\U_0/U_3/U_3/N87 ), .B(n3404), .C(\U_0/U_3/U_3/N62 ), .D(
        n3405), .Y(n3411) );
  OAI21X1 U4079 ( .A(n11118), .B(n3402), .C(n3413), .Y(n8499) );
  AOI22X1 U4080 ( .A(\U_0/U_3/U_3/N86 ), .B(n3404), .C(\U_0/U_3/U_3/N61 ), .D(
        n3405), .Y(n3413) );
  OAI21X1 U4081 ( .A(n11117), .B(n3402), .C(n3415), .Y(n8500) );
  AOI22X1 U4082 ( .A(\U_0/U_3/U_3/N85 ), .B(n3404), .C(\U_0/U_3/U_3/N60 ), .D(
        n3405), .Y(n3415) );
  OAI21X1 U4083 ( .A(n10012), .B(n11172), .C(n3418), .Y(n8501) );
  NAND2X1 U4084 ( .A(\U_0/U_0/U_0/N414 ), .B(n3419), .Y(n3418) );
  OAI21X1 U4085 ( .A(n10012), .B(n11180), .C(n3421), .Y(n8502) );
  NAND2X1 U4086 ( .A(\U_0/U_0/U_0/N413 ), .B(n3419), .Y(n3421) );
  OAI21X1 U4087 ( .A(n10012), .B(n11179), .C(n3423), .Y(n8503) );
  NAND2X1 U4088 ( .A(\U_0/U_0/U_0/N412 ), .B(n3419), .Y(n3423) );
  OAI21X1 U4089 ( .A(n10012), .B(n11178), .C(n3425), .Y(n8504) );
  NAND2X1 U4090 ( .A(\U_0/U_0/U_0/N411 ), .B(n3419), .Y(n3425) );
  OAI21X1 U4091 ( .A(n10012), .B(n11177), .C(n3427), .Y(n8505) );
  NAND2X1 U4092 ( .A(\U_0/U_0/U_0/N410 ), .B(n3419), .Y(n3427) );
  OAI21X1 U4093 ( .A(n10012), .B(n11176), .C(n3429), .Y(n8506) );
  NAND2X1 U4094 ( .A(\U_0/U_0/U_0/N409 ), .B(n3419), .Y(n3429) );
  OAI21X1 U4095 ( .A(n10012), .B(n11175), .C(n3431), .Y(n8507) );
  NAND2X1 U4096 ( .A(\U_0/U_0/U_0/N408 ), .B(n3419), .Y(n3431) );
  OAI21X1 U4097 ( .A(n10012), .B(n11174), .C(n3433), .Y(n8508) );
  NAND2X1 U4098 ( .A(\U_0/U_0/U_0/N407 ), .B(n3419), .Y(n3433) );
  NOR2X1 U4099 ( .A(n11155), .B(n3434), .Y(n3419) );
  OAI21X1 U4100 ( .A(n11148), .B(n3436), .C(n3437), .Y(n8509) );
  OAI21X1 U4101 ( .A(n3438), .B(n10042), .C(\U_0/U_0/U_0/permuteComplete ), 
        .Y(n3437) );
  NAND2X1 U4103 ( .A(n3441), .B(n3440), .Y(n3436) );
  NOR3X1 U4104 ( .A(n3442), .B(n3443), .C(n3444), .Y(n3440) );
  OAI21X1 U4105 ( .A(n11134), .B(n11241), .C(n3447), .Y(n8510) );
  NAND2X1 U4106 ( .A(\U_0/U_0/U_0/N431 ), .B(n3448), .Y(n3447) );
  OAI21X1 U4108 ( .A(n11134), .B(n11252), .C(n3450), .Y(n8511) );
  NAND2X1 U4109 ( .A(\U_0/U_0/U_0/N430 ), .B(n3448), .Y(n3450) );
  OAI21X1 U4111 ( .A(n11134), .B(n11251), .C(n3452), .Y(n8512) );
  NAND2X1 U4112 ( .A(\U_0/U_0/U_0/N429 ), .B(n3448), .Y(n3452) );
  OAI21X1 U4113 ( .A(n11134), .B(n11250), .C(n3454), .Y(n8513) );
  NAND2X1 U4114 ( .A(\U_0/U_0/U_0/N428 ), .B(n3448), .Y(n3454) );
  OAI21X1 U4115 ( .A(n11134), .B(n9543), .C(n3456), .Y(n8514) );
  NAND2X1 U4116 ( .A(\U_0/U_0/U_0/N427 ), .B(n3448), .Y(n3456) );
  OAI22X1 U4118 ( .A(n10043), .B(n11249), .C(n11248), .D(n3460), .Y(n8515) );
  OAI21X1 U4119 ( .A(n11134), .B(n11248), .C(n3461), .Y(n8516) );
  NAND2X1 U4120 ( .A(\U_0/U_0/U_0/N426 ), .B(n3448), .Y(n3461) );
  OAI22X1 U4122 ( .A(n10043), .B(n11245), .C(n9544), .D(n3460), .Y(n8517) );
  OAI21X1 U4123 ( .A(n11134), .B(n9544), .C(n3464), .Y(n8518) );
  NAND2X1 U4124 ( .A(\U_0/U_0/U_0/N425 ), .B(n3448), .Y(n3464) );
  OAI22X1 U4125 ( .A(n10043), .B(n11253), .C(n11242), .D(n3460), .Y(n8519) );
  NAND3X1 U4127 ( .A(n11158), .B(n9517), .C(n11134), .Y(n3460) );
  OAI21X1 U4128 ( .A(n11134), .B(n11242), .C(n3468), .Y(n8520) );
  NAND2X1 U4129 ( .A(\U_0/U_0/U_0/N424 ), .B(n3448), .Y(n3468) );
  NOR2X1 U4130 ( .A(n11148), .B(n3441), .Y(n3448) );
  NOR2X1 U4131 ( .A(n3469), .B(n3470), .Y(n3441) );
  NAND3X1 U4132 ( .A(\U_0/U_0/U_0/si[7] ), .B(\U_0/U_0/U_0/si[6] ), .C(n3471), 
        .Y(n3470) );
  NOR2X1 U4133 ( .A(n11250), .B(n11251), .Y(n3471) );
  NAND3X1 U4136 ( .A(\U_0/U_0/U_0/si[3] ), .B(\U_0/U_0/U_0/si[2] ), .C(n3472), 
        .Y(n3469) );
  NOR2X1 U4137 ( .A(n11242), .B(n9544), .Y(n3472) );
  NAND3X1 U4141 ( .A(n11138), .B(n11144), .C(n3475), .Y(n3473) );
  NOR2X1 U4142 ( .A(n3476), .B(n3477), .Y(n3475) );
  OAI21X1 U4143 ( .A(n11133), .B(n11197), .C(n3480), .Y(n8521) );
  NAND2X1 U4144 ( .A(\U_0/U_0/U_0/N480 ), .B(n3481), .Y(n3480) );
  OAI21X1 U4146 ( .A(n11133), .B(n11196), .C(n3483), .Y(n8522) );
  NAND2X1 U4147 ( .A(\U_0/U_0/U_0/N481 ), .B(n3481), .Y(n3483) );
  OAI21X1 U4149 ( .A(n11133), .B(n11195), .C(n3485), .Y(n8523) );
  NAND2X1 U4150 ( .A(\U_0/U_0/U_0/N482 ), .B(n3481), .Y(n3485) );
  OAI21X1 U4152 ( .A(n11133), .B(n11194), .C(n3487), .Y(n8524) );
  NAND2X1 U4153 ( .A(\U_0/U_0/U_0/N483 ), .B(n3481), .Y(n3487) );
  OAI21X1 U4155 ( .A(n11133), .B(n11193), .C(n3489), .Y(n8525) );
  NAND2X1 U4156 ( .A(\U_0/U_0/U_0/N484 ), .B(n3481), .Y(n3489) );
  OAI21X1 U4158 ( .A(n11133), .B(n11192), .C(n3491), .Y(n8526) );
  NAND2X1 U4159 ( .A(\U_0/U_0/U_0/N485 ), .B(n3481), .Y(n3491) );
  OAI21X1 U4161 ( .A(n11133), .B(n11191), .C(n3493), .Y(n8527) );
  NAND2X1 U4162 ( .A(\U_0/U_0/U_0/N486 ), .B(n3481), .Y(n3493) );
  OAI21X1 U4164 ( .A(n11133), .B(n11190), .C(n3495), .Y(n8528) );
  NAND2X1 U4165 ( .A(\U_0/U_0/U_0/N487 ), .B(n3481), .Y(n3495) );
  NAND3X1 U4168 ( .A(n11138), .B(n3497), .C(n3498), .Y(n3496) );
  NOR2X1 U4169 ( .A(n11143), .B(n3500), .Y(n3498) );
  NAND2X1 U4170 ( .A(n11141), .B(n11148), .Y(n3500) );
  NAND3X1 U4173 ( .A(n3503), .B(n3504), .C(n11139), .Y(n3502) );
  AOI22X1 U4175 ( .A(n3507), .B(\U_0/U_0/U_0/inti[7] ), .C(n3508), .D(
        \U_0/U_0/U_0/N503 ), .Y(n3506) );
  AOI22X1 U4177 ( .A(n3507), .B(\U_0/U_0/U_0/inti[6] ), .C(n3508), .D(
        \U_0/U_0/U_0/N502 ), .Y(n3509) );
  AOI22X1 U4179 ( .A(n3507), .B(\U_0/U_0/U_0/inti[5] ), .C(n3508), .D(
        \U_0/U_0/U_0/N501 ), .Y(n3510) );
  AOI22X1 U4181 ( .A(n3507), .B(\U_0/U_0/U_0/inti[4] ), .C(n3508), .D(
        \U_0/U_0/U_0/N500 ), .Y(n3511) );
  AOI22X1 U4183 ( .A(n3507), .B(\U_0/U_0/U_0/inti[3] ), .C(n3508), .D(
        \U_0/U_0/U_0/N499 ), .Y(n3512) );
  AOI22X1 U4185 ( .A(n3507), .B(\U_0/U_0/U_0/inti[2] ), .C(n3508), .D(
        \U_0/U_0/U_0/N498 ), .Y(n3513) );
  AOI22X1 U4187 ( .A(n3507), .B(\U_0/U_0/U_0/inti[1] ), .C(n3508), .D(
        \U_0/U_0/U_0/N497 ), .Y(n3514) );
  AOI22X1 U4189 ( .A(n3507), .B(\U_0/U_0/U_0/inti[0] ), .C(n3508), .D(
        \U_0/U_0/U_0/N496 ), .Y(n3515) );
  NOR2X1 U4190 ( .A(n9190), .B(n3507), .Y(n3508) );
  NAND3X1 U4191 ( .A(n11146), .B(n3518), .C(n10031), .Y(n3507) );
  OAI21X1 U4192 ( .A(n10021), .B(n11182), .C(n3522), .Y(n8537) );
  NAND2X1 U4193 ( .A(\U_0/U_0/U_0/N519 ), .B(n3523), .Y(n3522) );
  OAI21X1 U4195 ( .A(n10021), .B(n11189), .C(n3525), .Y(n8538) );
  NAND2X1 U4196 ( .A(\U_0/U_0/U_0/N518 ), .B(n3523), .Y(n3525) );
  OAI21X1 U4198 ( .A(n10021), .B(n11188), .C(n3527), .Y(n8539) );
  NAND2X1 U4199 ( .A(\U_0/U_0/U_0/N517 ), .B(n3523), .Y(n3527) );
  OAI21X1 U4201 ( .A(n10021), .B(n11187), .C(n3529), .Y(n8540) );
  NAND2X1 U4202 ( .A(\U_0/U_0/U_0/N516 ), .B(n3523), .Y(n3529) );
  OAI21X1 U4204 ( .A(n10021), .B(n11186), .C(n3531), .Y(n8541) );
  NAND2X1 U4205 ( .A(\U_0/U_0/U_0/N515 ), .B(n3523), .Y(n3531) );
  OAI21X1 U4207 ( .A(n10021), .B(n11185), .C(n3533), .Y(n8542) );
  NAND2X1 U4208 ( .A(\U_0/U_0/U_0/N514 ), .B(n3523), .Y(n3533) );
  OAI21X1 U4210 ( .A(n10021), .B(n11184), .C(n3535), .Y(n8543) );
  NAND2X1 U4211 ( .A(\U_0/U_0/U_0/N513 ), .B(n3523), .Y(n3535) );
  OAI21X1 U4213 ( .A(n10021), .B(n11183), .C(n3537), .Y(n8544) );
  NAND2X1 U4214 ( .A(\U_0/U_0/U_0/N512 ), .B(n3523), .Y(n3537) );
  NOR2X1 U4215 ( .A(n3518), .B(n3538), .Y(n3523) );
  OAI21X1 U4218 ( .A(n10041), .B(n11205), .C(n3541), .Y(n8545) );
  AOI22X1 U4219 ( .A(DATA_IN_H[7]), .B(n3542), .C(\U_0/U_0/U_0/N527 ), .D(
        n3543), .Y(n3541) );
  OAI21X1 U4220 ( .A(n10041), .B(n11204), .C(n3545), .Y(n8546) );
  AOI22X1 U4221 ( .A(DATA_IN_H[5]), .B(n3542), .C(\U_0/U_0/U_0/N525 ), .D(
        n3543), .Y(n3545) );
  OAI21X1 U4222 ( .A(n10041), .B(n11203), .C(n3547), .Y(n8547) );
  AOI22X1 U4223 ( .A(DATA_IN_H[4]), .B(n3542), .C(\U_0/U_0/U_0/N524 ), .D(
        n3543), .Y(n3547) );
  OAI21X1 U4224 ( .A(n10041), .B(n11202), .C(n3549), .Y(n8548) );
  AOI22X1 U4225 ( .A(DATA_IN_H[3]), .B(n3542), .C(\U_0/U_0/U_0/N523 ), .D(
        n3543), .Y(n3549) );
  OAI21X1 U4226 ( .A(n10041), .B(n11201), .C(n3551), .Y(n8549) );
  AOI22X1 U4227 ( .A(DATA_IN_H[2]), .B(n3542), .C(\U_0/U_0/U_0/N522 ), .D(
        n3543), .Y(n3551) );
  OAI21X1 U4228 ( .A(n10041), .B(n11200), .C(n3553), .Y(n8550) );
  AOI22X1 U4229 ( .A(DATA_IN_H[1]), .B(n3542), .C(\U_0/U_0/U_0/N521 ), .D(
        n3543), .Y(n3553) );
  OAI21X1 U4230 ( .A(n10041), .B(n11199), .C(n3555), .Y(n8551) );
  AOI22X1 U4231 ( .A(DATA_IN_H[0]), .B(n3542), .C(\U_0/U_0/U_0/N520 ), .D(
        n3543), .Y(n3555) );
  OAI21X1 U4232 ( .A(n10041), .B(n11198), .C(n3557), .Y(n8552) );
  AOI22X1 U4233 ( .A(DATA_IN_H[6]), .B(n3542), .C(\U_0/U_0/U_0/N526 ), .D(
        n3543), .Y(n3557) );
  NOR2X1 U4234 ( .A(n3558), .B(n3559), .Y(n3543) );
  AOI21X1 U4235 ( .A(n11131), .B(n3501), .C(n3559), .Y(n3542) );
  NAND3X1 U4237 ( .A(n3561), .B(n562), .C(n3562), .Y(n3559) );
  NOR2X1 U4238 ( .A(n3563), .B(n3442), .Y(n3562) );
  NAND3X1 U4239 ( .A(n11139), .B(n9189), .C(n3565), .Y(n3442) );
  NAND3X1 U4242 ( .A(n11159), .B(n11151), .C(n607), .Y(n3566) );
  NOR2X1 U4243 ( .A(n3569), .B(n3570), .Y(n607) );
  AOI22X1 U4247 ( .A(n3574), .B(\U_0/U_0/U_0/extratemp[0] ), .C(DATA_IN_H[0]), 
        .D(n9238), .Y(n3573) );
  AOI22X1 U4249 ( .A(n3574), .B(\U_0/U_0/U_0/extratemp[1] ), .C(DATA_IN_H[1]), 
        .D(n9238), .Y(n3576) );
  AOI22X1 U4251 ( .A(n3574), .B(\U_0/U_0/U_0/extratemp[2] ), .C(DATA_IN_H[2]), 
        .D(n9238), .Y(n3577) );
  AOI22X1 U4253 ( .A(n3574), .B(\U_0/U_0/U_0/extratemp[3] ), .C(DATA_IN_H[3]), 
        .D(n9238), .Y(n3578) );
  AOI22X1 U4255 ( .A(n3574), .B(\U_0/U_0/U_0/extratemp[4] ), .C(DATA_IN_H[4]), 
        .D(n9238), .Y(n3579) );
  AOI22X1 U4257 ( .A(n3574), .B(\U_0/U_0/U_0/extratemp[5] ), .C(DATA_IN_H[5]), 
        .D(n9238), .Y(n3580) );
  AOI22X1 U4259 ( .A(n3574), .B(\U_0/U_0/U_0/extratemp[6] ), .C(DATA_IN_H[6]), 
        .D(n9238), .Y(n3581) );
  AOI22X1 U4261 ( .A(n3574), .B(\U_0/U_0/U_0/extratemp[7] ), .C(DATA_IN_H[7]), 
        .D(n9238), .Y(n3582) );
  NAND3X1 U4263 ( .A(n11158), .B(n3583), .C(n3584), .Y(n3574) );
  NOR2X1 U4264 ( .A(n3585), .B(n3586), .Y(n3584) );
  AOI22X1 U4266 ( .A(\U_0/U_0/PLAINKEY [6]), .B(n9431), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[0][6] ), .Y(n3587) );
  AOI22X1 U4268 ( .A(\U_0/U_0/PLAINKEY [5]), .B(n9424), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[0][5] ), .Y(n3590) );
  AOI22X1 U4270 ( .A(\U_0/U_0/PLAINKEY [4]), .B(n9424), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[0][4] ), .Y(n3591) );
  OAI22X1 U4271 ( .A(n10789), .B(n9423), .C(n9436), .D(n11258), .Y(n8564) );
  OAI22X1 U4273 ( .A(n10787), .B(n9422), .C(n9436), .D(n11259), .Y(n8565) );
  OAI22X1 U4275 ( .A(n10785), .B(n9421), .C(n9436), .D(n11260), .Y(n8566) );
  OAI22X1 U4277 ( .A(n10783), .B(n9421), .C(n9436), .D(n11261), .Y(n8567) );
  AOI22X1 U4280 ( .A(\U_0/U_0/PLAINKEY [15]), .B(n9425), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[1][7] ), .Y(n3596) );
  AOI22X1 U4282 ( .A(\U_0/U_0/PLAINKEY [7]), .B(n9425), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[0][7] ), .Y(n3597) );
  AOI22X1 U4284 ( .A(\U_0/U_0/PLAINKEY [56]), .B(n9425), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[7][0] ), .Y(n3598) );
  AOI22X1 U4286 ( .A(\U_0/U_0/PLAINKEY [57]), .B(n9426), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[7][1] ), .Y(n3599) );
  AOI22X1 U4288 ( .A(\U_0/U_0/PLAINKEY [58]), .B(n9426), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[7][2] ), .Y(n3600) );
  AOI22X1 U4290 ( .A(\U_0/U_0/PLAINKEY [59]), .B(n9426), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[7][3] ), .Y(n3601) );
  AOI22X1 U4292 ( .A(\U_0/U_0/PLAINKEY [60]), .B(n9427), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[7][4] ), .Y(n3602) );
  AOI22X1 U4294 ( .A(\U_0/U_0/PLAINKEY [61]), .B(n9427), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[7][5] ), .Y(n3603) );
  AOI22X1 U4296 ( .A(\U_0/U_0/PLAINKEY [62]), .B(n9427), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[7][6] ), .Y(n3604) );
  AOI22X1 U4298 ( .A(\U_0/U_0/PLAINKEY [63]), .B(n9428), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[7][7] ), .Y(n3605) );
  AOI22X1 U4300 ( .A(\U_0/U_0/PLAINKEY [48]), .B(n9428), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[6][0] ), .Y(n3606) );
  AOI22X1 U4302 ( .A(\U_0/U_0/PLAINKEY [49]), .B(n9428), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[6][1] ), .Y(n3607) );
  AOI22X1 U4304 ( .A(\U_0/U_0/PLAINKEY [50]), .B(n9429), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[6][2] ), .Y(n3608) );
  AOI22X1 U4306 ( .A(\U_0/U_0/PLAINKEY [51]), .B(n9429), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[6][3] ), .Y(n3609) );
  AOI22X1 U4308 ( .A(\U_0/U_0/PLAINKEY [52]), .B(n9429), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[6][4] ), .Y(n3610) );
  AOI22X1 U4310 ( .A(\U_0/U_0/PLAINKEY [53]), .B(n9430), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[6][5] ), .Y(n3611) );
  AOI22X1 U4312 ( .A(\U_0/U_0/PLAINKEY [54]), .B(n9430), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[6][6] ), .Y(n3612) );
  AOI22X1 U4314 ( .A(\U_0/U_0/PLAINKEY [55]), .B(n9430), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[6][7] ), .Y(n3613) );
  AOI22X1 U4316 ( .A(\U_0/U_0/PLAINKEY [40]), .B(n9430), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[5][0] ), .Y(n3614) );
  AOI22X1 U4318 ( .A(\U_0/U_0/PLAINKEY [41]), .B(n9430), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[5][1] ), .Y(n3615) );
  AOI22X1 U4320 ( .A(\U_0/U_0/PLAINKEY [42]), .B(n9430), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[5][2] ), .Y(n3616) );
  AOI22X1 U4322 ( .A(\U_0/U_0/PLAINKEY [43]), .B(n9430), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[5][3] ), .Y(n3617) );
  AOI22X1 U4324 ( .A(\U_0/U_0/PLAINKEY [44]), .B(n9431), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[5][4] ), .Y(n3618) );
  AOI22X1 U4326 ( .A(\U_0/U_0/PLAINKEY [45]), .B(n9431), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[5][5] ), .Y(n3619) );
  AOI22X1 U4328 ( .A(\U_0/U_0/PLAINKEY [46]), .B(n9431), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[5][6] ), .Y(n3620) );
  AOI22X1 U4330 ( .A(\U_0/U_0/PLAINKEY [47]), .B(n9431), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[5][7] ), .Y(n3621) );
  AOI22X1 U4332 ( .A(\U_0/U_0/PLAINKEY [32]), .B(n9431), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[4][0] ), .Y(n3622) );
  AOI22X1 U4334 ( .A(\U_0/U_0/PLAINKEY [33]), .B(n9431), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[4][1] ), .Y(n3623) );
  AOI22X1 U4336 ( .A(\U_0/U_0/PLAINKEY [34]), .B(n9432), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[4][2] ), .Y(n3624) );
  AOI22X1 U4338 ( .A(\U_0/U_0/PLAINKEY [35]), .B(n9432), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[4][3] ), .Y(n3625) );
  AOI22X1 U4340 ( .A(\U_0/U_0/PLAINKEY [36]), .B(n9432), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[4][4] ), .Y(n3626) );
  AOI22X1 U4342 ( .A(\U_0/U_0/PLAINKEY [37]), .B(n9432), .C(n9421), .D(
        \U_0/U_0/U_0/keyTable[4][5] ), .Y(n3627) );
  AOI22X1 U4344 ( .A(\U_0/U_0/PLAINKEY [38]), .B(n9432), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[4][6] ), .Y(n3628) );
  AOI22X1 U4346 ( .A(\U_0/U_0/PLAINKEY [39]), .B(n9432), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[4][7] ), .Y(n3629) );
  AOI22X1 U4348 ( .A(\U_0/U_0/PLAINKEY [24]), .B(n9432), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[3][0] ), .Y(n3630) );
  AOI22X1 U4350 ( .A(\U_0/U_0/PLAINKEY [25]), .B(n9433), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[3][1] ), .Y(n3631) );
  AOI22X1 U4352 ( .A(\U_0/U_0/PLAINKEY [26]), .B(n9433), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[3][2] ), .Y(n3632) );
  AOI22X1 U4354 ( .A(\U_0/U_0/PLAINKEY [27]), .B(n9433), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[3][3] ), .Y(n3633) );
  AOI22X1 U4356 ( .A(\U_0/U_0/PLAINKEY [28]), .B(n9433), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[3][4] ), .Y(n3634) );
  AOI22X1 U4358 ( .A(\U_0/U_0/PLAINKEY [29]), .B(n9433), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[3][5] ), .Y(n3635) );
  AOI22X1 U4360 ( .A(\U_0/U_0/PLAINKEY [30]), .B(n9433), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[3][6] ), .Y(n3636) );
  AOI22X1 U4362 ( .A(\U_0/U_0/PLAINKEY [31]), .B(n9433), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[3][7] ), .Y(n3637) );
  AOI22X1 U4364 ( .A(\U_0/U_0/PLAINKEY [16]), .B(n9434), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[2][0] ), .Y(n3638) );
  AOI22X1 U4366 ( .A(\U_0/U_0/PLAINKEY [17]), .B(n9434), .C(n9422), .D(
        \U_0/U_0/U_0/keyTable[2][1] ), .Y(n3639) );
  AOI22X1 U4368 ( .A(\U_0/U_0/PLAINKEY [18]), .B(n9434), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[2][2] ), .Y(n3640) );
  AOI22X1 U4370 ( .A(\U_0/U_0/PLAINKEY [19]), .B(n9434), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[2][3] ), .Y(n3641) );
  AOI22X1 U4372 ( .A(\U_0/U_0/PLAINKEY [20]), .B(n9434), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[2][4] ), .Y(n3642) );
  AOI22X1 U4374 ( .A(\U_0/U_0/PLAINKEY [21]), .B(n9434), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[2][5] ), .Y(n3643) );
  AOI22X1 U4376 ( .A(\U_0/U_0/PLAINKEY [22]), .B(n9434), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[2][6] ), .Y(n3644) );
  AOI22X1 U4378 ( .A(\U_0/U_0/PLAINKEY [23]), .B(n9435), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[2][7] ), .Y(n3645) );
  AOI22X1 U4380 ( .A(\U_0/U_0/PLAINKEY [8]), .B(n9435), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[1][0] ), .Y(n3646) );
  AOI22X1 U4382 ( .A(\U_0/U_0/PLAINKEY [9]), .B(n9435), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[1][1] ), .Y(n3647) );
  AOI22X1 U4384 ( .A(\U_0/U_0/PLAINKEY [10]), .B(n9435), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[1][2] ), .Y(n3648) );
  AOI22X1 U4386 ( .A(\U_0/U_0/PLAINKEY [11]), .B(n9435), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[1][3] ), .Y(n3649) );
  AOI22X1 U4388 ( .A(\U_0/U_0/PLAINKEY [12]), .B(n9435), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[1][4] ), .Y(n3650) );
  AOI22X1 U4390 ( .A(\U_0/U_0/PLAINKEY [13]), .B(n9435), .C(n9423), .D(
        \U_0/U_0/U_0/keyTable[1][5] ), .Y(n3651) );
  AOI22X1 U4392 ( .A(\U_0/U_0/PLAINKEY [14]), .B(n9424), .C(n3589), .D(
        \U_0/U_0/U_0/keyTable[1][6] ), .Y(n3652) );
  NAND2X1 U4394 ( .A(n10012), .B(n3504), .Y(n3589) );
  NAND3X1 U4396 ( .A(n11146), .B(n10040), .C(n3654), .Y(n3434) );
  NOR2X1 U4397 ( .A(n3655), .B(n3585), .Y(n3654) );
  AOI22X1 U4399 ( .A(n10030), .B(\U_0/U_0/U_0/delaydata [6]), .C(
        \U_0/PRGA_IN [6]), .D(n3658), .Y(n3656) );
  AOI22X1 U4401 ( .A(n10030), .B(\U_0/U_0/U_0/delaydata [5]), .C(
        \U_0/PRGA_IN [5]), .D(n3658), .Y(n3659) );
  AOI22X1 U4403 ( .A(n10030), .B(\U_0/U_0/U_0/delaydata [4]), .C(
        \U_0/PRGA_IN [4]), .D(n3658), .Y(n3660) );
  AOI22X1 U4405 ( .A(n10030), .B(\U_0/U_0/U_0/delaydata [3]), .C(
        \U_0/PRGA_IN [3]), .D(n3658), .Y(n3661) );
  AOI22X1 U4407 ( .A(n10030), .B(\U_0/U_0/U_0/delaydata [2]), .C(
        \U_0/PRGA_IN [2]), .D(n3658), .Y(n3662) );
  AOI22X1 U4409 ( .A(n10030), .B(\U_0/U_0/U_0/delaydata [1]), .C(
        \U_0/PRGA_IN [1]), .D(n3658), .Y(n3663) );
  AOI22X1 U4411 ( .A(n10030), .B(\U_0/U_0/U_0/delaydata [0]), .C(
        \U_0/PRGA_IN [0]), .D(n3658), .Y(n3664) );
  AOI22X1 U4413 ( .A(n10030), .B(\U_0/U_0/U_0/delaydata [7]), .C(
        \U_0/PRGA_IN [7]), .D(n3658), .Y(n3665) );
  NOR2X1 U4415 ( .A(n3538), .B(n3655), .Y(n3658) );
  NAND3X1 U4416 ( .A(n11146), .B(n9190), .C(n10031), .Y(n3538) );
  NAND3X1 U4418 ( .A(n11155), .B(n3504), .C(n10040), .Y(n3586) );
  NAND3X1 U4420 ( .A(n3497), .B(n3667), .C(n3668), .Y(n3666) );
  AOI21X1 U4421 ( .A(n3669), .B(n3670), .C(n3671), .Y(n3668) );
  NAND2X1 U4422 ( .A(n3672), .B(n9496), .Y(n3671) );
  NOR3X1 U4423 ( .A(n3476), .B(n3673), .C(n3477), .Y(n3497) );
  OAI21X1 U4425 ( .A(n9951), .B(n11088), .C(n3676), .Y(n8633) );
  OAI21X1 U4426 ( .A(n3677), .B(n3678), .C(n9951), .Y(n3676) );
  NAND3X1 U4428 ( .A(n3681), .B(n3682), .C(n3683), .Y(n3680) );
  NOR2X1 U4429 ( .A(n3684), .B(n3685), .Y(n3683) );
  OAI22X1 U4430 ( .A(n3686), .B(n11019), .C(n3688), .D(n11029), .Y(n3685) );
  OAI22X1 U4431 ( .A(n3690), .B(n10999), .C(n3692), .D(n11009), .Y(n3684) );
  AOI22X1 U4432 ( .A(\U_0/U_1/U_1/opcode[26][1] ), .B(n3694), .C(
        \U_0/U_1/U_1/opcode[27][1] ), .D(n3695), .Y(n3682) );
  AOI22X1 U4433 ( .A(\U_0/U_1/U_1/opcode[24][1] ), .B(n3696), .C(
        \U_0/U_1/U_1/opcode[25][1] ), .D(n3697), .Y(n3681) );
  NAND3X1 U4434 ( .A(n3698), .B(n3699), .C(n3700), .Y(n3679) );
  NOR2X1 U4435 ( .A(n3701), .B(n3702), .Y(n3700) );
  OAI22X1 U4436 ( .A(n3703), .B(n11059), .C(n3705), .D(n11069), .Y(n3702) );
  OAI22X1 U4437 ( .A(n3707), .B(n11039), .C(n3709), .D(n11049), .Y(n3701) );
  AOI22X1 U4438 ( .A(\U_0/U_1/U_1/opcode[22][1] ), .B(n3711), .C(
        \U_0/U_1/U_1/opcode[23][1] ), .D(n3712), .Y(n3699) );
  AOI22X1 U4439 ( .A(\U_0/U_1/U_1/opcode[20][1] ), .B(n3713), .C(
        \U_0/U_1/U_1/opcode[21][1] ), .D(n3714), .Y(n3698) );
  NAND3X1 U4441 ( .A(n3717), .B(n3718), .C(n3719), .Y(n3716) );
  NOR2X1 U4442 ( .A(n3720), .B(n3721), .Y(n3719) );
  OAI22X1 U4443 ( .A(n3722), .B(n10989), .C(n3724), .D(n10954), .Y(n3721) );
  OAI22X1 U4444 ( .A(n3726), .B(n10969), .C(n3728), .D(n10979), .Y(n3720) );
  AOI22X1 U4445 ( .A(\U_0/U_1/U_1/opcode[14][1] ), .B(n3730), .C(
        \U_0/U_1/U_1/opcode[15][1] ), .D(n3731), .Y(n3718) );
  AOI22X1 U4446 ( .A(\U_0/U_1/U_1/opcode[12][1] ), .B(n3732), .C(
        \U_0/U_1/U_1/opcode[13][1] ), .D(n3733), .Y(n3717) );
  NAND3X1 U4447 ( .A(n3734), .B(n3735), .C(n3736), .Y(n3715) );
  NOR2X1 U4448 ( .A(n3737), .B(n3738), .Y(n3736) );
  OAI22X1 U4449 ( .A(n3739), .B(n10929), .C(n3741), .D(n10919), .Y(n3738) );
  OAI22X1 U4450 ( .A(n3743), .B(n10959), .C(n3745), .D(n10957), .Y(n3737) );
  AOI22X1 U4451 ( .A(\U_0/U_1/U_1/opcode[1][1] ), .B(n3747), .C(
        \U_0/U_1/U_1/opcode[0][1] ), .D(n3748), .Y(n3735) );
  AOI22X1 U4452 ( .A(\U_0/U_1/U_1/opcode[3][1] ), .B(n3749), .C(
        \U_0/U_1/U_1/opcode[2][1] ), .D(n3750), .Y(n3734) );
  OAI21X1 U4454 ( .A(n9951), .B(n11087), .C(n3751), .Y(n8634) );
  OAI21X1 U4455 ( .A(n3752), .B(n3753), .C(n9951), .Y(n3751) );
  NAND3X1 U4457 ( .A(n3756), .B(n3757), .C(n3758), .Y(n3755) );
  NOR2X1 U4458 ( .A(n3759), .B(n3760), .Y(n3758) );
  OAI22X1 U4459 ( .A(n3686), .B(n11018), .C(n3688), .D(n11028), .Y(n3760) );
  OAI22X1 U4460 ( .A(n3690), .B(n10998), .C(n3692), .D(n11008), .Y(n3759) );
  AOI22X1 U4461 ( .A(\U_0/U_1/U_1/opcode[26][0] ), .B(n3694), .C(
        \U_0/U_1/U_1/opcode[27][0] ), .D(n3695), .Y(n3757) );
  AOI22X1 U4462 ( .A(\U_0/U_1/U_1/opcode[24][0] ), .B(n3696), .C(
        \U_0/U_1/U_1/opcode[25][0] ), .D(n3697), .Y(n3756) );
  NAND3X1 U4463 ( .A(n3765), .B(n3766), .C(n3767), .Y(n3754) );
  NOR2X1 U4464 ( .A(n3768), .B(n3769), .Y(n3767) );
  OAI22X1 U4465 ( .A(n3703), .B(n11058), .C(n3705), .D(n11068), .Y(n3769) );
  OAI22X1 U4466 ( .A(n3707), .B(n11038), .C(n3709), .D(n11048), .Y(n3768) );
  AOI22X1 U4467 ( .A(\U_0/U_1/U_1/opcode[22][0] ), .B(n3711), .C(
        \U_0/U_1/U_1/opcode[23][0] ), .D(n3712), .Y(n3766) );
  AOI22X1 U4468 ( .A(\U_0/U_1/U_1/opcode[20][0] ), .B(n3713), .C(
        \U_0/U_1/U_1/opcode[21][0] ), .D(n3714), .Y(n3765) );
  NAND3X1 U4470 ( .A(n3776), .B(n3777), .C(n3778), .Y(n3775) );
  NOR2X1 U4471 ( .A(n3779), .B(n3780), .Y(n3778) );
  OAI22X1 U4472 ( .A(n3722), .B(n10988), .C(n3724), .D(n10955), .Y(n3780) );
  OAI22X1 U4473 ( .A(n3726), .B(n10968), .C(n3728), .D(n10978), .Y(n3779) );
  AOI22X1 U4474 ( .A(\U_0/U_1/U_1/opcode[14][0] ), .B(n3730), .C(
        \U_0/U_1/U_1/opcode[15][0] ), .D(n3731), .Y(n3777) );
  AOI22X1 U4475 ( .A(\U_0/U_1/U_1/opcode[12][0] ), .B(n3732), .C(
        \U_0/U_1/U_1/opcode[13][0] ), .D(n3733), .Y(n3776) );
  NAND3X1 U4476 ( .A(n3785), .B(n3786), .C(n3787), .Y(n3774) );
  NOR2X1 U4477 ( .A(n3788), .B(n3789), .Y(n3787) );
  OAI22X1 U4478 ( .A(n3739), .B(n10928), .C(n3741), .D(n10918), .Y(n3789) );
  OAI22X1 U4479 ( .A(n3743), .B(n10958), .C(n3745), .D(n10956), .Y(n3788) );
  AOI22X1 U4480 ( .A(\U_0/U_1/U_1/opcode[1][0] ), .B(n3747), .C(
        \U_0/U_1/U_1/opcode[0][0] ), .D(n3748), .Y(n3786) );
  AOI22X1 U4481 ( .A(\U_0/U_1/U_1/opcode[3][0] ), .B(n3749), .C(
        \U_0/U_1/U_1/opcode[2][0] ), .D(n3750), .Y(n3785) );
  OAI21X1 U4483 ( .A(n9951), .B(n11086), .C(n3794), .Y(n8635) );
  OAI21X1 U4484 ( .A(n3795), .B(n3796), .C(n9951), .Y(n3794) );
  NAND3X1 U4486 ( .A(n3799), .B(n3800), .C(n3801), .Y(n3798) );
  NOR2X1 U4487 ( .A(n3802), .B(n3803), .Y(n3801) );
  OAI22X1 U4488 ( .A(n3686), .B(n11027), .C(n3688), .D(n11037), .Y(n3803) );
  OAI22X1 U4489 ( .A(n3690), .B(n11007), .C(n3692), .D(n11017), .Y(n3802) );
  AOI22X1 U4490 ( .A(\U_0/U_1/U_1/memory[26][7] ), .B(n3694), .C(
        \U_0/U_1/U_1/memory[27][7] ), .D(n3695), .Y(n3800) );
  AOI22X1 U4491 ( .A(\U_0/U_1/U_1/memory[24][7] ), .B(n3696), .C(
        \U_0/U_1/U_1/memory[25][7] ), .D(n3697), .Y(n3799) );
  NAND3X1 U4492 ( .A(n3808), .B(n3809), .C(n3810), .Y(n3797) );
  NOR2X1 U4493 ( .A(n3811), .B(n3812), .Y(n3810) );
  OAI22X1 U4494 ( .A(n3703), .B(n11067), .C(n3705), .D(n11074), .Y(n3812) );
  OAI22X1 U4495 ( .A(n3707), .B(n11047), .C(n3709), .D(n11057), .Y(n3811) );
  AOI22X1 U4496 ( .A(\U_0/U_1/U_1/memory[22][7] ), .B(n3711), .C(
        \U_0/U_1/U_1/memory[23][7] ), .D(n3712), .Y(n3809) );
  AOI22X1 U4497 ( .A(\U_0/U_1/U_1/memory[20][7] ), .B(n3713), .C(
        \U_0/U_1/U_1/memory[21][7] ), .D(n3714), .Y(n3808) );
  NAND3X1 U4499 ( .A(n3819), .B(n3820), .C(n3821), .Y(n3818) );
  NOR2X1 U4500 ( .A(n3822), .B(n3823), .Y(n3821) );
  OAI22X1 U4501 ( .A(n3722), .B(n10997), .C(n3724), .D(n10967), .Y(n3823) );
  OAI22X1 U4502 ( .A(n3726), .B(n10977), .C(n3728), .D(n10987), .Y(n3822) );
  AOI22X1 U4503 ( .A(\U_0/U_1/U_1/memory[14][7] ), .B(n3730), .C(
        \U_0/U_1/U_1/memory[15][7] ), .D(n3731), .Y(n3820) );
  AOI22X1 U4504 ( .A(\U_0/U_1/U_1/memory[12][7] ), .B(n3732), .C(
        \U_0/U_1/U_1/memory[13][7] ), .D(n3733), .Y(n3819) );
  NAND3X1 U4505 ( .A(n3828), .B(n3829), .C(n3830), .Y(n3817) );
  NOR2X1 U4506 ( .A(n3831), .B(n3832), .Y(n3830) );
  OAI22X1 U4507 ( .A(n3739), .B(n10937), .C(n3741), .D(n10927), .Y(n3832) );
  OAI22X1 U4508 ( .A(n3743), .B(n10947), .C(n3745), .D(n10945), .Y(n3831) );
  AOI22X1 U4509 ( .A(\U_0/U_1/U_1/memory[1][7] ), .B(n3747), .C(
        \U_0/U_1/U_1/memory[0][7] ), .D(n3748), .Y(n3829) );
  AOI22X1 U4510 ( .A(\U_0/U_1/U_1/memory[3][7] ), .B(n3749), .C(
        \U_0/U_1/U_1/memory[2][7] ), .D(n3750), .Y(n3828) );
  OAI21X1 U4512 ( .A(n9951), .B(n11085), .C(n3837), .Y(n8636) );
  OAI21X1 U4513 ( .A(n3838), .B(n3839), .C(n9951), .Y(n3837) );
  NAND3X1 U4515 ( .A(n3842), .B(n3843), .C(n3844), .Y(n3841) );
  NOR2X1 U4516 ( .A(n3845), .B(n3846), .Y(n3844) );
  OAI22X1 U4517 ( .A(n3686), .B(n11026), .C(n3688), .D(n11036), .Y(n3846) );
  OAI22X1 U4518 ( .A(n3690), .B(n11006), .C(n3692), .D(n11016), .Y(n3845) );
  AOI22X1 U4519 ( .A(\U_0/U_1/U_1/memory[26][6] ), .B(n3694), .C(
        \U_0/U_1/U_1/memory[27][6] ), .D(n3695), .Y(n3843) );
  AOI22X1 U4520 ( .A(\U_0/U_1/U_1/memory[24][6] ), .B(n3696), .C(
        \U_0/U_1/U_1/memory[25][6] ), .D(n3697), .Y(n3842) );
  NAND3X1 U4521 ( .A(n3851), .B(n3852), .C(n3853), .Y(n3840) );
  NOR2X1 U4522 ( .A(n3854), .B(n3855), .Y(n3853) );
  OAI22X1 U4523 ( .A(n3703), .B(n11066), .C(n3705), .D(n11073), .Y(n3855) );
  OAI22X1 U4524 ( .A(n3707), .B(n11046), .C(n3709), .D(n11056), .Y(n3854) );
  AOI22X1 U4525 ( .A(\U_0/U_1/U_1/memory[22][6] ), .B(n3711), .C(
        \U_0/U_1/U_1/memory[23][6] ), .D(n3712), .Y(n3852) );
  AOI22X1 U4526 ( .A(\U_0/U_1/U_1/memory[20][6] ), .B(n3713), .C(
        \U_0/U_1/U_1/memory[21][6] ), .D(n3714), .Y(n3851) );
  NAND3X1 U4528 ( .A(n3862), .B(n3863), .C(n3864), .Y(n3861) );
  NOR2X1 U4529 ( .A(n3865), .B(n3866), .Y(n3864) );
  OAI22X1 U4530 ( .A(n3722), .B(n10996), .C(n3724), .D(n10966), .Y(n3866) );
  OAI22X1 U4531 ( .A(n3726), .B(n10976), .C(n3728), .D(n10986), .Y(n3865) );
  AOI22X1 U4532 ( .A(\U_0/U_1/U_1/memory[14][6] ), .B(n3730), .C(
        \U_0/U_1/U_1/memory[15][6] ), .D(n3731), .Y(n3863) );
  AOI22X1 U4533 ( .A(\U_0/U_1/U_1/memory[12][6] ), .B(n3732), .C(
        \U_0/U_1/U_1/memory[13][6] ), .D(n3733), .Y(n3862) );
  NAND3X1 U4534 ( .A(n3871), .B(n3872), .C(n3873), .Y(n3860) );
  NOR2X1 U4535 ( .A(n3874), .B(n3875), .Y(n3873) );
  OAI22X1 U4536 ( .A(n3739), .B(n10936), .C(n3741), .D(n10926), .Y(n3875) );
  OAI22X1 U4537 ( .A(n3743), .B(n10946), .C(n3745), .D(n10944), .Y(n3874) );
  AOI22X1 U4538 ( .A(\U_0/U_1/U_1/memory[1][6] ), .B(n3747), .C(
        \U_0/U_1/U_1/memory[0][6] ), .D(n3748), .Y(n3872) );
  AOI22X1 U4539 ( .A(\U_0/U_1/U_1/memory[3][6] ), .B(n3749), .C(
        \U_0/U_1/U_1/memory[2][6] ), .D(n3750), .Y(n3871) );
  OAI21X1 U4541 ( .A(n9951), .B(n11084), .C(n3880), .Y(n8637) );
  OAI21X1 U4542 ( .A(n3881), .B(n3882), .C(n9951), .Y(n3880) );
  NAND3X1 U4544 ( .A(n3885), .B(n3886), .C(n3887), .Y(n3884) );
  NOR2X1 U4545 ( .A(n3888), .B(n3889), .Y(n3887) );
  OAI22X1 U4546 ( .A(n3686), .B(n11025), .C(n3688), .D(n11035), .Y(n3889) );
  OAI22X1 U4547 ( .A(n3690), .B(n11005), .C(n3692), .D(n11015), .Y(n3888) );
  AOI22X1 U4548 ( .A(\U_0/U_1/U_1/memory[26][5] ), .B(n3694), .C(
        \U_0/U_1/U_1/memory[27][5] ), .D(n3695), .Y(n3886) );
  AOI22X1 U4549 ( .A(\U_0/U_1/U_1/memory[24][5] ), .B(n3696), .C(
        \U_0/U_1/U_1/memory[25][5] ), .D(n3697), .Y(n3885) );
  NAND3X1 U4550 ( .A(n3894), .B(n3895), .C(n3896), .Y(n3883) );
  NOR2X1 U4551 ( .A(n3897), .B(n3898), .Y(n3896) );
  OAI22X1 U4552 ( .A(n3703), .B(n11065), .C(n3705), .D(n11072), .Y(n3898) );
  OAI22X1 U4553 ( .A(n3707), .B(n11045), .C(n3709), .D(n11055), .Y(n3897) );
  AOI22X1 U4554 ( .A(\U_0/U_1/U_1/memory[22][5] ), .B(n3711), .C(
        \U_0/U_1/U_1/memory[23][5] ), .D(n3712), .Y(n3895) );
  AOI22X1 U4555 ( .A(\U_0/U_1/U_1/memory[20][5] ), .B(n3713), .C(
        \U_0/U_1/U_1/memory[21][5] ), .D(n3714), .Y(n3894) );
  NAND3X1 U4557 ( .A(n3905), .B(n3906), .C(n3907), .Y(n3904) );
  NOR2X1 U4558 ( .A(n3908), .B(n3909), .Y(n3907) );
  OAI22X1 U4559 ( .A(n3722), .B(n10995), .C(n3724), .D(n10965), .Y(n3909) );
  OAI22X1 U4560 ( .A(n3726), .B(n10975), .C(n3728), .D(n10985), .Y(n3908) );
  AOI22X1 U4561 ( .A(\U_0/U_1/U_1/memory[14][5] ), .B(n3730), .C(
        \U_0/U_1/U_1/memory[15][5] ), .D(n3731), .Y(n3906) );
  AOI22X1 U4562 ( .A(\U_0/U_1/U_1/memory[12][5] ), .B(n3732), .C(
        \U_0/U_1/U_1/memory[13][5] ), .D(n3733), .Y(n3905) );
  NAND3X1 U4563 ( .A(n3914), .B(n3915), .C(n3916), .Y(n3903) );
  NOR2X1 U4564 ( .A(n3917), .B(n3918), .Y(n3916) );
  OAI22X1 U4565 ( .A(n3739), .B(n10935), .C(n3741), .D(n10925), .Y(n3918) );
  OAI22X1 U4566 ( .A(n3743), .B(n10953), .C(n3745), .D(n10943), .Y(n3917) );
  AOI22X1 U4567 ( .A(\U_0/U_1/U_1/memory[1][5] ), .B(n3747), .C(
        \U_0/U_1/U_1/memory[0][5] ), .D(n3748), .Y(n3915) );
  AOI22X1 U4568 ( .A(\U_0/U_1/U_1/memory[3][5] ), .B(n3749), .C(
        \U_0/U_1/U_1/memory[2][5] ), .D(n3750), .Y(n3914) );
  OAI21X1 U4570 ( .A(n9951), .B(n11083), .C(n3923), .Y(n8638) );
  OAI21X1 U4571 ( .A(n3924), .B(n3925), .C(n9951), .Y(n3923) );
  NAND3X1 U4573 ( .A(n3928), .B(n3929), .C(n3930), .Y(n3927) );
  NOR2X1 U4574 ( .A(n3931), .B(n3932), .Y(n3930) );
  OAI22X1 U4575 ( .A(n3686), .B(n11024), .C(n3688), .D(n11034), .Y(n3932) );
  OAI22X1 U4576 ( .A(n3690), .B(n11004), .C(n3692), .D(n11014), .Y(n3931) );
  AOI22X1 U4577 ( .A(\U_0/U_1/U_1/memory[26][4] ), .B(n3694), .C(
        \U_0/U_1/U_1/memory[27][4] ), .D(n3695), .Y(n3929) );
  AOI22X1 U4578 ( .A(\U_0/U_1/U_1/memory[24][4] ), .B(n3696), .C(
        \U_0/U_1/U_1/memory[25][4] ), .D(n3697), .Y(n3928) );
  NAND3X1 U4579 ( .A(n3937), .B(n3938), .C(n3939), .Y(n3926) );
  NOR2X1 U4580 ( .A(n3940), .B(n3941), .Y(n3939) );
  OAI22X1 U4581 ( .A(n3703), .B(n11064), .C(n3705), .D(n11071), .Y(n3941) );
  OAI22X1 U4582 ( .A(n3707), .B(n11044), .C(n3709), .D(n11054), .Y(n3940) );
  AOI22X1 U4583 ( .A(\U_0/U_1/U_1/memory[22][4] ), .B(n3711), .C(
        \U_0/U_1/U_1/memory[23][4] ), .D(n3712), .Y(n3938) );
  AOI22X1 U4584 ( .A(\U_0/U_1/U_1/memory[20][4] ), .B(n3713), .C(
        \U_0/U_1/U_1/memory[21][4] ), .D(n3714), .Y(n3937) );
  NAND3X1 U4586 ( .A(n3948), .B(n3949), .C(n3950), .Y(n3947) );
  NOR2X1 U4587 ( .A(n3951), .B(n3952), .Y(n3950) );
  OAI22X1 U4588 ( .A(n3722), .B(n10994), .C(n3724), .D(n10964), .Y(n3952) );
  OAI22X1 U4589 ( .A(n3726), .B(n10974), .C(n3728), .D(n10984), .Y(n3951) );
  AOI22X1 U4590 ( .A(\U_0/U_1/U_1/memory[14][4] ), .B(n3730), .C(
        \U_0/U_1/U_1/memory[15][4] ), .D(n3731), .Y(n3949) );
  AOI22X1 U4591 ( .A(\U_0/U_1/U_1/memory[12][4] ), .B(n3732), .C(
        \U_0/U_1/U_1/memory[13][4] ), .D(n3733), .Y(n3948) );
  NAND3X1 U4592 ( .A(n3957), .B(n3958), .C(n3959), .Y(n3946) );
  NOR2X1 U4593 ( .A(n3960), .B(n3961), .Y(n3959) );
  OAI22X1 U4594 ( .A(n3739), .B(n10934), .C(n3741), .D(n10924), .Y(n3961) );
  OAI22X1 U4595 ( .A(n3743), .B(n10952), .C(n3745), .D(n10942), .Y(n3960) );
  AOI22X1 U4596 ( .A(\U_0/U_1/U_1/memory[1][4] ), .B(n3747), .C(
        \U_0/U_1/U_1/memory[0][4] ), .D(n3748), .Y(n3958) );
  AOI22X1 U4597 ( .A(\U_0/U_1/U_1/memory[3][4] ), .B(n3749), .C(
        \U_0/U_1/U_1/memory[2][4] ), .D(n3750), .Y(n3957) );
  OAI21X1 U4599 ( .A(n9951), .B(n11082), .C(n3966), .Y(n8639) );
  OAI21X1 U4600 ( .A(n3967), .B(n3968), .C(n9951), .Y(n3966) );
  NAND3X1 U4602 ( .A(n3971), .B(n3972), .C(n3973), .Y(n3970) );
  NOR2X1 U4603 ( .A(n3974), .B(n3975), .Y(n3973) );
  OAI22X1 U4604 ( .A(n3686), .B(n11023), .C(n3688), .D(n11033), .Y(n3975) );
  OAI22X1 U4605 ( .A(n3690), .B(n11003), .C(n3692), .D(n11013), .Y(n3974) );
  AOI22X1 U4606 ( .A(\U_0/U_1/U_1/memory[26][3] ), .B(n3694), .C(
        \U_0/U_1/U_1/memory[27][3] ), .D(n3695), .Y(n3972) );
  AOI22X1 U4607 ( .A(\U_0/U_1/U_1/memory[24][3] ), .B(n3696), .C(
        \U_0/U_1/U_1/memory[25][3] ), .D(n3697), .Y(n3971) );
  NAND3X1 U4608 ( .A(n3980), .B(n3981), .C(n3982), .Y(n3969) );
  NOR2X1 U4609 ( .A(n3983), .B(n3984), .Y(n3982) );
  OAI22X1 U4610 ( .A(n3703), .B(n11063), .C(n3705), .D(n11070), .Y(n3984) );
  OAI22X1 U4611 ( .A(n3707), .B(n11043), .C(n3709), .D(n11053), .Y(n3983) );
  AOI22X1 U4612 ( .A(\U_0/U_1/U_1/memory[22][3] ), .B(n3711), .C(
        \U_0/U_1/U_1/memory[23][3] ), .D(n3712), .Y(n3981) );
  AOI22X1 U4613 ( .A(\U_0/U_1/U_1/memory[20][3] ), .B(n3713), .C(
        \U_0/U_1/U_1/memory[21][3] ), .D(n3714), .Y(n3980) );
  NAND3X1 U4615 ( .A(n3991), .B(n3992), .C(n3993), .Y(n3990) );
  NOR2X1 U4616 ( .A(n3994), .B(n3995), .Y(n3993) );
  OAI22X1 U4617 ( .A(n3722), .B(n10993), .C(n3724), .D(n10963), .Y(n3995) );
  OAI22X1 U4618 ( .A(n3726), .B(n10973), .C(n3728), .D(n10983), .Y(n3994) );
  AOI22X1 U4619 ( .A(\U_0/U_1/U_1/memory[14][3] ), .B(n3730), .C(
        \U_0/U_1/U_1/memory[15][3] ), .D(n3731), .Y(n3992) );
  AOI22X1 U4620 ( .A(\U_0/U_1/U_1/memory[12][3] ), .B(n3732), .C(
        \U_0/U_1/U_1/memory[13][3] ), .D(n3733), .Y(n3991) );
  NAND3X1 U4621 ( .A(n4000), .B(n4001), .C(n4002), .Y(n3989) );
  NOR2X1 U4622 ( .A(n4003), .B(n4004), .Y(n4002) );
  OAI22X1 U4623 ( .A(n3739), .B(n10933), .C(n3741), .D(n10923), .Y(n4004) );
  OAI22X1 U4624 ( .A(n3743), .B(n10951), .C(n3745), .D(n10941), .Y(n4003) );
  AOI22X1 U4625 ( .A(\U_0/U_1/U_1/memory[1][3] ), .B(n3747), .C(
        \U_0/U_1/U_1/memory[0][3] ), .D(n3748), .Y(n4001) );
  AOI22X1 U4626 ( .A(\U_0/U_1/U_1/memory[3][3] ), .B(n3749), .C(
        \U_0/U_1/U_1/memory[2][3] ), .D(n3750), .Y(n4000) );
  OAI21X1 U4628 ( .A(n9951), .B(n11081), .C(n4009), .Y(n8640) );
  OAI21X1 U4629 ( .A(n4010), .B(n4011), .C(n9951), .Y(n4009) );
  NAND3X1 U4631 ( .A(n4014), .B(n4015), .C(n4016), .Y(n4013) );
  NOR2X1 U4632 ( .A(n4017), .B(n4018), .Y(n4016) );
  OAI22X1 U4633 ( .A(n3686), .B(n11022), .C(n3688), .D(n11032), .Y(n4018) );
  OAI22X1 U4634 ( .A(n3690), .B(n11002), .C(n3692), .D(n11012), .Y(n4017) );
  AOI22X1 U4635 ( .A(\U_0/U_1/U_1/memory[26][2] ), .B(n3694), .C(
        \U_0/U_1/U_1/memory[27][2] ), .D(n3695), .Y(n4015) );
  AOI22X1 U4636 ( .A(\U_0/U_1/U_1/memory[24][2] ), .B(n3696), .C(
        \U_0/U_1/U_1/memory[25][2] ), .D(n3697), .Y(n4014) );
  NAND3X1 U4637 ( .A(n4023), .B(n4024), .C(n4025), .Y(n4012) );
  NOR2X1 U4638 ( .A(n4026), .B(n4027), .Y(n4025) );
  OAI22X1 U4639 ( .A(n3703), .B(n11062), .C(n3705), .D(n11077), .Y(n4027) );
  OAI22X1 U4640 ( .A(n3707), .B(n11042), .C(n3709), .D(n11052), .Y(n4026) );
  AOI22X1 U4641 ( .A(\U_0/U_1/U_1/memory[22][2] ), .B(n3711), .C(
        \U_0/U_1/U_1/memory[23][2] ), .D(n3712), .Y(n4024) );
  AOI22X1 U4642 ( .A(\U_0/U_1/U_1/memory[20][2] ), .B(n3713), .C(
        \U_0/U_1/U_1/memory[21][2] ), .D(n3714), .Y(n4023) );
  NAND3X1 U4644 ( .A(n4034), .B(n4035), .C(n4036), .Y(n4033) );
  NOR2X1 U4645 ( .A(n4037), .B(n4038), .Y(n4036) );
  OAI22X1 U4646 ( .A(n3722), .B(n10992), .C(n3724), .D(n10962), .Y(n4038) );
  OAI22X1 U4647 ( .A(n3726), .B(n10972), .C(n3728), .D(n10982), .Y(n4037) );
  AOI22X1 U4648 ( .A(\U_0/U_1/U_1/memory[14][2] ), .B(n3730), .C(
        \U_0/U_1/U_1/memory[15][2] ), .D(n3731), .Y(n4035) );
  AOI22X1 U4649 ( .A(\U_0/U_1/U_1/memory[12][2] ), .B(n3732), .C(
        \U_0/U_1/U_1/memory[13][2] ), .D(n3733), .Y(n4034) );
  NAND3X1 U4650 ( .A(n4043), .B(n4044), .C(n4045), .Y(n4032) );
  NOR2X1 U4651 ( .A(n4046), .B(n4047), .Y(n4045) );
  OAI22X1 U4652 ( .A(n3739), .B(n10932), .C(n3741), .D(n10922), .Y(n4047) );
  OAI22X1 U4653 ( .A(n3743), .B(n10950), .C(n3745), .D(n10940), .Y(n4046) );
  AOI22X1 U4654 ( .A(\U_0/U_1/U_1/memory[1][2] ), .B(n3747), .C(
        \U_0/U_1/U_1/memory[0][2] ), .D(n3748), .Y(n4044) );
  AOI22X1 U4655 ( .A(\U_0/U_1/U_1/memory[3][2] ), .B(n3749), .C(
        \U_0/U_1/U_1/memory[2][2] ), .D(n3750), .Y(n4043) );
  OAI21X1 U4657 ( .A(n9951), .B(n11080), .C(n4052), .Y(n8641) );
  OAI21X1 U4658 ( .A(n4053), .B(n4054), .C(n9951), .Y(n4052) );
  NAND3X1 U4660 ( .A(n4057), .B(n4058), .C(n4059), .Y(n4056) );
  NOR2X1 U4661 ( .A(n4060), .B(n4061), .Y(n4059) );
  OAI22X1 U4662 ( .A(n3686), .B(n11021), .C(n3688), .D(n11031), .Y(n4061) );
  OAI22X1 U4663 ( .A(n3690), .B(n11001), .C(n3692), .D(n11011), .Y(n4060) );
  AOI22X1 U4664 ( .A(\U_0/U_1/U_1/memory[26][1] ), .B(n3694), .C(
        \U_0/U_1/U_1/memory[27][1] ), .D(n3695), .Y(n4058) );
  AOI22X1 U4665 ( .A(\U_0/U_1/U_1/memory[24][1] ), .B(n3696), .C(
        \U_0/U_1/U_1/memory[25][1] ), .D(n3697), .Y(n4057) );
  NAND3X1 U4666 ( .A(n4066), .B(n4067), .C(n4068), .Y(n4055) );
  NOR2X1 U4667 ( .A(n4069), .B(n4070), .Y(n4068) );
  OAI22X1 U4668 ( .A(n3703), .B(n11061), .C(n3705), .D(n11076), .Y(n4070) );
  OAI22X1 U4669 ( .A(n3707), .B(n11041), .C(n3709), .D(n11051), .Y(n4069) );
  AOI22X1 U4670 ( .A(\U_0/U_1/U_1/memory[22][1] ), .B(n3711), .C(
        \U_0/U_1/U_1/memory[23][1] ), .D(n3712), .Y(n4067) );
  AOI22X1 U4671 ( .A(\U_0/U_1/U_1/memory[20][1] ), .B(n3713), .C(
        \U_0/U_1/U_1/memory[21][1] ), .D(n3714), .Y(n4066) );
  NAND3X1 U4673 ( .A(n4077), .B(n4078), .C(n4079), .Y(n4076) );
  NOR2X1 U4674 ( .A(n4080), .B(n4081), .Y(n4079) );
  OAI22X1 U4675 ( .A(n3722), .B(n10991), .C(n3724), .D(n10961), .Y(n4081) );
  OAI22X1 U4676 ( .A(n3726), .B(n10971), .C(n3728), .D(n10981), .Y(n4080) );
  AOI22X1 U4677 ( .A(\U_0/U_1/U_1/memory[14][1] ), .B(n3730), .C(
        \U_0/U_1/U_1/memory[15][1] ), .D(n3731), .Y(n4078) );
  AOI22X1 U4678 ( .A(\U_0/U_1/U_1/memory[12][1] ), .B(n3732), .C(
        \U_0/U_1/U_1/memory[13][1] ), .D(n3733), .Y(n4077) );
  NAND3X1 U4679 ( .A(n4086), .B(n4087), .C(n4088), .Y(n4075) );
  NOR2X1 U4680 ( .A(n4089), .B(n4090), .Y(n4088) );
  OAI22X1 U4681 ( .A(n3739), .B(n10931), .C(n3741), .D(n10921), .Y(n4090) );
  OAI22X1 U4682 ( .A(n3743), .B(n10949), .C(n3745), .D(n10939), .Y(n4089) );
  AOI22X1 U4683 ( .A(\U_0/U_1/U_1/memory[1][1] ), .B(n3747), .C(
        \U_0/U_1/U_1/memory[0][1] ), .D(n3748), .Y(n4087) );
  AOI22X1 U4684 ( .A(\U_0/U_1/U_1/memory[3][1] ), .B(n3749), .C(
        \U_0/U_1/U_1/memory[2][1] ), .D(n3750), .Y(n4086) );
  OAI21X1 U4686 ( .A(n9951), .B(n11079), .C(n4095), .Y(n8642) );
  OAI21X1 U4687 ( .A(n4096), .B(n4097), .C(n9951), .Y(n4095) );
  NAND3X1 U4689 ( .A(n4100), .B(n4101), .C(n4102), .Y(n4099) );
  NOR2X1 U4690 ( .A(n4103), .B(n4104), .Y(n4102) );
  OAI22X1 U4691 ( .A(n3686), .B(n11020), .C(n3688), .D(n11030), .Y(n4104) );
  NAND2X1 U4692 ( .A(n10913), .B(n4108), .Y(n3688) );
  NAND2X1 U4693 ( .A(n10909), .B(n4108), .Y(n3686) );
  OAI22X1 U4694 ( .A(n3690), .B(n11000), .C(n3692), .D(n11010), .Y(n4103) );
  NAND2X1 U4695 ( .A(n10913), .B(n4112), .Y(n3692) );
  NAND2X1 U4696 ( .A(n10909), .B(n4112), .Y(n3690) );
  AOI22X1 U4697 ( .A(\U_0/U_1/U_1/memory[26][0] ), .B(n3694), .C(
        \U_0/U_1/U_1/memory[27][0] ), .D(n3695), .Y(n4101) );
  AOI22X1 U4700 ( .A(\U_0/U_1/U_1/memory[24][0] ), .B(n3696), .C(
        \U_0/U_1/U_1/memory[25][0] ), .D(n3697), .Y(n4100) );
  NAND3X1 U4703 ( .A(n9331), .B(\U_0/U_1/U_1/readptr[0] ), .C(
        \U_0/U_1/U_1/readptr[4] ), .Y(n4115) );
  NAND3X1 U4706 ( .A(n9331), .B(n9334), .C(\U_0/U_1/U_1/readptr[4] ), .Y(n4116) );
  NAND3X1 U4707 ( .A(n4118), .B(n4119), .C(n4120), .Y(n4098) );
  NOR2X1 U4708 ( .A(n4121), .B(n4122), .Y(n4120) );
  OAI22X1 U4709 ( .A(n3703), .B(n11060), .C(n3705), .D(n11075), .Y(n4122) );
  NAND2X1 U4710 ( .A(n10914), .B(n4113), .Y(n3705) );
  NAND2X1 U4711 ( .A(n10910), .B(n4113), .Y(n3703) );
  OAI22X1 U4712 ( .A(n3707), .B(n11040), .C(n3709), .D(n11050), .Y(n4121) );
  NAND2X1 U4713 ( .A(n10914), .B(n4114), .Y(n3709) );
  NAND2X1 U4714 ( .A(n10910), .B(n4114), .Y(n3707) );
  AOI22X1 U4715 ( .A(\U_0/U_1/U_1/memory[22][0] ), .B(n3711), .C(
        \U_0/U_1/U_1/memory[23][0] ), .D(n3712), .Y(n4119) );
  AOI22X1 U4718 ( .A(\U_0/U_1/U_1/memory[20][0] ), .B(n3713), .C(
        \U_0/U_1/U_1/memory[21][0] ), .D(n3714), .Y(n4118) );
  NAND3X1 U4721 ( .A(\U_0/U_1/U_1/readptr[0] ), .B(n9330), .C(
        \U_0/U_1/U_1/readptr[4] ), .Y(n4129) );
  NAND3X1 U4724 ( .A(n9334), .B(n9330), .C(\U_0/U_1/U_1/readptr[4] ), .Y(n4131) );
  NAND3X1 U4726 ( .A(n4134), .B(n4135), .C(n4136), .Y(n4133) );
  NOR2X1 U4727 ( .A(n4137), .B(n4138), .Y(n4136) );
  OAI22X1 U4728 ( .A(n3722), .B(n10990), .C(n3724), .D(n10960), .Y(n4138) );
  NAND2X1 U4729 ( .A(n10915), .B(n4113), .Y(n3724) );
  NAND2X1 U4730 ( .A(n10911), .B(n4113), .Y(n3722) );
  OAI22X1 U4731 ( .A(n3726), .B(n10970), .C(n3728), .D(n10980), .Y(n4137) );
  NAND2X1 U4732 ( .A(n10915), .B(n4114), .Y(n3728) );
  NAND2X1 U4733 ( .A(n10911), .B(n4114), .Y(n3726) );
  AOI22X1 U4734 ( .A(\U_0/U_1/U_1/memory[14][0] ), .B(n3730), .C(
        \U_0/U_1/U_1/memory[15][0] ), .D(n3731), .Y(n4135) );
  AOI22X1 U4737 ( .A(\U_0/U_1/U_1/memory[12][0] ), .B(n3732), .C(
        \U_0/U_1/U_1/memory[13][0] ), .D(n3733), .Y(n4134) );
  NAND3X1 U4740 ( .A(\U_0/U_1/U_1/readptr[0] ), .B(n9329), .C(n9331), .Y(n4145) );
  NAND3X1 U4743 ( .A(n9334), .B(n9329), .C(n9331), .Y(n4147) );
  NAND3X1 U4744 ( .A(n4148), .B(n4149), .C(n4150), .Y(n4132) );
  NOR2X1 U4745 ( .A(n4151), .B(n4152), .Y(n4150) );
  OAI22X1 U4746 ( .A(n3739), .B(n10930), .C(n3741), .D(n10920), .Y(n4152) );
  NAND2X1 U4747 ( .A(n4112), .B(n10912), .Y(n3741) );
  NAND2X1 U4748 ( .A(n4112), .B(n10916), .Y(n3739) );
  OAI22X1 U4750 ( .A(n3743), .B(n10948), .C(n3745), .D(n10938), .Y(n4151) );
  NAND2X1 U4751 ( .A(n4108), .B(n10912), .Y(n3745) );
  NAND2X1 U4752 ( .A(n4108), .B(n10916), .Y(n3743) );
  AOI22X1 U4754 ( .A(\U_0/U_1/U_1/memory[1][0] ), .B(n3747), .C(
        \U_0/U_1/U_1/memory[0][0] ), .D(n3748), .Y(n4149) );
  NOR2X1 U4757 ( .A(\U_0/U_1/U_1/readptr[1] ), .B(\U_0/U_1/U_1/readptr[2] ), 
        .Y(n4114) );
  AOI22X1 U4758 ( .A(\U_0/U_1/U_1/memory[3][0] ), .B(n3749), .C(
        \U_0/U_1/U_1/memory[2][0] ), .D(n3750), .Y(n4148) );
  NAND3X1 U4761 ( .A(n9330), .B(n9329), .C(n9334), .Y(n4160) );
  NAND3X1 U4765 ( .A(n9330), .B(n9329), .C(\U_0/U_1/U_1/readptr[0] ), .Y(n4161) );
  NOR2X1 U4768 ( .A(n9333), .B(\U_0/U_1/U_1/readptr[2] ), .Y(n4113) );
  NAND3X1 U4772 ( .A(\U_0/U_1/U_1/N195 ), .B(n9519), .C(n9353), .Y(n4162) );
  AOI22X1 U4774 ( .A(n9949), .B(\U_0/U_1/U_1/memory[0][7] ), .C(n9352), .D(
        n4165), .Y(n4163) );
  AOI22X1 U4776 ( .A(n9949), .B(\U_0/U_1/U_1/memory[0][6] ), .C(n4165), .D(
        \U_0/RCV_DATA [6]), .Y(n4166) );
  AOI22X1 U4778 ( .A(n9949), .B(\U_0/U_1/U_1/memory[0][5] ), .C(n4165), .D(
        n9348), .Y(n4167) );
  AOI22X1 U4780 ( .A(n9949), .B(\U_0/U_1/U_1/memory[0][4] ), .C(n4165), .D(
        n9346), .Y(n4168) );
  AOI22X1 U4782 ( .A(n9949), .B(\U_0/U_1/U_1/memory[0][3] ), .C(n4165), .D(
        n9344), .Y(n4169) );
  AOI22X1 U4784 ( .A(n9949), .B(\U_0/U_1/U_1/memory[0][2] ), .C(n4165), .D(
        n9342), .Y(n4170) );
  AOI22X1 U4786 ( .A(n9949), .B(\U_0/U_1/U_1/memory[0][1] ), .C(n4165), .D(
        n9340), .Y(n4171) );
  AOI22X1 U4788 ( .A(n9949), .B(\U_0/U_1/U_1/memory[0][0] ), .C(n4165), .D(
        n9338), .Y(n4172) );
  AOI22X1 U4790 ( .A(n9940), .B(\U_0/U_1/U_1/memory[1][7] ), .C(
        \U_0/RCV_DATA [7]), .D(n4175), .Y(n4173) );
  AOI22X1 U4792 ( .A(n9940), .B(\U_0/U_1/U_1/memory[1][6] ), .C(
        \U_0/RCV_DATA [6]), .D(n4175), .Y(n4176) );
  AOI22X1 U4794 ( .A(n9940), .B(\U_0/U_1/U_1/memory[1][5] ), .C(
        \U_0/RCV_DATA [5]), .D(n4175), .Y(n4177) );
  AOI22X1 U4796 ( .A(n9940), .B(\U_0/U_1/U_1/memory[1][4] ), .C(n9346), .D(
        n4175), .Y(n4178) );
  AOI22X1 U4798 ( .A(n9940), .B(\U_0/U_1/U_1/memory[1][3] ), .C(n9344), .D(
        n4175), .Y(n4179) );
  AOI22X1 U4800 ( .A(n9940), .B(\U_0/U_1/U_1/memory[1][2] ), .C(
        \U_0/RCV_DATA [2]), .D(n4175), .Y(n4180) );
  AOI22X1 U4802 ( .A(n9940), .B(\U_0/U_1/U_1/memory[1][1] ), .C(
        \U_0/RCV_DATA [1]), .D(n4175), .Y(n4181) );
  AOI22X1 U4804 ( .A(n9940), .B(\U_0/U_1/U_1/memory[1][0] ), .C(n9338), .D(
        n4175), .Y(n4182) );
  AOI22X1 U4806 ( .A(n9931), .B(\U_0/U_1/U_1/memory[2][7] ), .C(n9352), .D(
        n4185), .Y(n4183) );
  AOI22X1 U4808 ( .A(n9931), .B(\U_0/U_1/U_1/memory[2][6] ), .C(
        \U_0/RCV_DATA [6]), .D(n4185), .Y(n4186) );
  AOI22X1 U4810 ( .A(n9931), .B(\U_0/U_1/U_1/memory[2][5] ), .C(n9348), .D(
        n4185), .Y(n4187) );
  AOI22X1 U4812 ( .A(n9931), .B(\U_0/U_1/U_1/memory[2][4] ), .C(n9346), .D(
        n4185), .Y(n4188) );
  AOI22X1 U4814 ( .A(n9931), .B(\U_0/U_1/U_1/memory[2][3] ), .C(n9344), .D(
        n4185), .Y(n4189) );
  AOI22X1 U4816 ( .A(n9931), .B(\U_0/U_1/U_1/memory[2][2] ), .C(n9342), .D(
        n4185), .Y(n4190) );
  AOI22X1 U4818 ( .A(n9931), .B(\U_0/U_1/U_1/memory[2][1] ), .C(n9340), .D(
        n4185), .Y(n4191) );
  AOI22X1 U4820 ( .A(n9931), .B(\U_0/U_1/U_1/memory[2][0] ), .C(n9338), .D(
        n4185), .Y(n4192) );
  AOI22X1 U4822 ( .A(n9922), .B(\U_0/U_1/U_1/memory[3][7] ), .C(
        \U_0/RCV_DATA [7]), .D(n4195), .Y(n4193) );
  AOI22X1 U4824 ( .A(n9922), .B(\U_0/U_1/U_1/memory[3][6] ), .C(
        \U_0/RCV_DATA [6]), .D(n4195), .Y(n4196) );
  AOI22X1 U4826 ( .A(n9922), .B(\U_0/U_1/U_1/memory[3][5] ), .C(
        \U_0/RCV_DATA [5]), .D(n4195), .Y(n4197) );
  AOI22X1 U4828 ( .A(n9922), .B(\U_0/U_1/U_1/memory[3][4] ), .C(n9346), .D(
        n4195), .Y(n4198) );
  AOI22X1 U4830 ( .A(n9922), .B(\U_0/U_1/U_1/memory[3][3] ), .C(n9344), .D(
        n4195), .Y(n4199) );
  AOI22X1 U4832 ( .A(n9922), .B(\U_0/U_1/U_1/memory[3][2] ), .C(
        \U_0/RCV_DATA [2]), .D(n4195), .Y(n4200) );
  AOI22X1 U4834 ( .A(n9922), .B(\U_0/U_1/U_1/memory[3][1] ), .C(
        \U_0/RCV_DATA [1]), .D(n4195), .Y(n4201) );
  AOI22X1 U4836 ( .A(n9922), .B(\U_0/U_1/U_1/memory[3][0] ), .C(n9338), .D(
        n4195), .Y(n4202) );
  OAI22X1 U4837 ( .A(n4203), .B(n10927), .C(n9351), .D(n9913), .Y(n8675) );
  OAI22X1 U4839 ( .A(n4203), .B(n10926), .C(n9349), .D(n9913), .Y(n8676) );
  OAI22X1 U4841 ( .A(n4203), .B(n10925), .C(n9347), .D(n9913), .Y(n8677) );
  OAI22X1 U4843 ( .A(n4203), .B(n10924), .C(n9345), .D(n9913), .Y(n8678) );
  OAI22X1 U4845 ( .A(n4203), .B(n10923), .C(n9343), .D(n9913), .Y(n8679) );
  OAI22X1 U4847 ( .A(n4203), .B(n10922), .C(n9341), .D(n9913), .Y(n8680) );
  OAI22X1 U4849 ( .A(n4203), .B(n10921), .C(n9339), .D(n9913), .Y(n8681) );
  OAI22X1 U4851 ( .A(n4203), .B(n10920), .C(n9337), .D(n9913), .Y(n8682) );
  OAI22X1 U4853 ( .A(n4213), .B(n10937), .C(n9351), .D(n9912), .Y(n8683) );
  OAI22X1 U4855 ( .A(n4213), .B(n10936), .C(n9349), .D(n9912), .Y(n8684) );
  OAI22X1 U4857 ( .A(n4213), .B(n10935), .C(n9347), .D(n9912), .Y(n8685) );
  OAI22X1 U4859 ( .A(n4213), .B(n10934), .C(n9345), .D(n9912), .Y(n8686) );
  OAI22X1 U4861 ( .A(n4213), .B(n10933), .C(n9343), .D(n9912), .Y(n8687) );
  OAI22X1 U4863 ( .A(n4213), .B(n10932), .C(n9341), .D(n9912), .Y(n8688) );
  OAI22X1 U4865 ( .A(n4213), .B(n10931), .C(n9339), .D(n9912), .Y(n8689) );
  OAI22X1 U4867 ( .A(n4213), .B(n10930), .C(n9337), .D(n9912), .Y(n8690) );
  OAI22X1 U4869 ( .A(n4215), .B(n10945), .C(n9351), .D(n9911), .Y(n8691) );
  OAI22X1 U4871 ( .A(n4215), .B(n10944), .C(n9349), .D(n9911), .Y(n8692) );
  OAI22X1 U4873 ( .A(n4215), .B(n10943), .C(n9347), .D(n9911), .Y(n8693) );
  OAI22X1 U4875 ( .A(n4215), .B(n10942), .C(n9345), .D(n9911), .Y(n8694) );
  OAI22X1 U4877 ( .A(n4215), .B(n10941), .C(n9343), .D(n9911), .Y(n8695) );
  OAI22X1 U4879 ( .A(n4215), .B(n10940), .C(n9341), .D(n9911), .Y(n8696) );
  OAI22X1 U4881 ( .A(n4215), .B(n10939), .C(n9339), .D(n9911), .Y(n8697) );
  OAI22X1 U4883 ( .A(n4215), .B(n10938), .C(n9337), .D(n9911), .Y(n8698) );
  OAI22X1 U4885 ( .A(n4217), .B(n10953), .C(n9347), .D(n9910), .Y(n8699) );
  OAI22X1 U4887 ( .A(n4217), .B(n10952), .C(n9345), .D(n9910), .Y(n8700) );
  OAI22X1 U4889 ( .A(n4217), .B(n10951), .C(n9343), .D(n9910), .Y(n8701) );
  OAI22X1 U4891 ( .A(n4217), .B(n10950), .C(n9341), .D(n9910), .Y(n8702) );
  OAI22X1 U4893 ( .A(n4217), .B(n10949), .C(n9339), .D(n9910), .Y(n8703) );
  OAI22X1 U4895 ( .A(n4217), .B(n10948), .C(n9337), .D(n9910), .Y(n8704) );
  OAI22X1 U4897 ( .A(n4217), .B(n10947), .C(n9351), .D(n9910), .Y(n8705) );
  OAI22X1 U4899 ( .A(n4217), .B(n10946), .C(n9349), .D(n9910), .Y(n8706) );
  OAI22X1 U4901 ( .A(n9236), .B(n10977), .C(n9351), .D(n9908), .Y(n8707) );
  OAI22X1 U4903 ( .A(n9236), .B(n10976), .C(n9349), .D(n9908), .Y(n8708) );
  OAI22X1 U4905 ( .A(n9236), .B(n10975), .C(n9347), .D(n9908), .Y(n8709) );
  OAI22X1 U4907 ( .A(n9236), .B(n10974), .C(n9345), .D(n9908), .Y(n8710) );
  OAI22X1 U4909 ( .A(n9236), .B(n10973), .C(n9343), .D(n9908), .Y(n8711) );
  OAI22X1 U4911 ( .A(n9236), .B(n10972), .C(n9341), .D(n9908), .Y(n8712) );
  OAI22X1 U4913 ( .A(n9236), .B(n10971), .C(n9339), .D(n9908), .Y(n8713) );
  OAI22X1 U4915 ( .A(n9236), .B(n10970), .C(n9337), .D(n9908), .Y(n8714) );
  OAI22X1 U4917 ( .A(n9235), .B(n10987), .C(n9351), .D(n9907), .Y(n8715) );
  OAI22X1 U4919 ( .A(n9235), .B(n10986), .C(n9349), .D(n9907), .Y(n8716) );
  OAI22X1 U4921 ( .A(n9235), .B(n10985), .C(n9347), .D(n9907), .Y(n8717) );
  OAI22X1 U4923 ( .A(n9235), .B(n10984), .C(n9345), .D(n9907), .Y(n8718) );
  OAI22X1 U4925 ( .A(n9235), .B(n10983), .C(n9343), .D(n9907), .Y(n8719) );
  OAI22X1 U4927 ( .A(n9235), .B(n10982), .C(n9341), .D(n9907), .Y(n8720) );
  OAI22X1 U4929 ( .A(n9235), .B(n10981), .C(n9339), .D(n9907), .Y(n8721) );
  OAI22X1 U4931 ( .A(n9235), .B(n10980), .C(n9337), .D(n9907), .Y(n8722) );
  OAI22X1 U4933 ( .A(n9234), .B(n10997), .C(n9351), .D(n9906), .Y(n8723) );
  OAI22X1 U4935 ( .A(n9234), .B(n10996), .C(n9349), .D(n9906), .Y(n8724) );
  OAI22X1 U4937 ( .A(n9234), .B(n10995), .C(n9347), .D(n9906), .Y(n8725) );
  OAI22X1 U4939 ( .A(n9234), .B(n10994), .C(n9345), .D(n9906), .Y(n8726) );
  OAI22X1 U4941 ( .A(n9234), .B(n10993), .C(n9343), .D(n9906), .Y(n8727) );
  OAI22X1 U4943 ( .A(n9234), .B(n10992), .C(n9341), .D(n9906), .Y(n8728) );
  OAI22X1 U4945 ( .A(n9234), .B(n10991), .C(n9339), .D(n9906), .Y(n8729) );
  OAI22X1 U4947 ( .A(n9234), .B(n10990), .C(n9337), .D(n9906), .Y(n8730) );
  OAI22X1 U4949 ( .A(n9237), .B(n10967), .C(n9351), .D(n9909), .Y(n8731) );
  OAI22X1 U4951 ( .A(n9237), .B(n10966), .C(n9349), .D(n9909), .Y(n8732) );
  OAI22X1 U4953 ( .A(n9237), .B(n10965), .C(n9347), .D(n9909), .Y(n8733) );
  OAI22X1 U4955 ( .A(n9237), .B(n10964), .C(n9345), .D(n9909), .Y(n8734) );
  OAI22X1 U4957 ( .A(n9237), .B(n10963), .C(n9343), .D(n9909), .Y(n8735) );
  OAI22X1 U4959 ( .A(n9237), .B(n10962), .C(n9341), .D(n9909), .Y(n8736) );
  OAI22X1 U4961 ( .A(n9237), .B(n10961), .C(n9339), .D(n9909), .Y(n8737) );
  OAI22X1 U4963 ( .A(n9237), .B(n10960), .C(n9337), .D(n9909), .Y(n8738) );
  NOR2X1 U4966 ( .A(n4227), .B(n4228), .Y(n4225) );
  AOI22X1 U4968 ( .A(n9905), .B(\U_0/U_1/U_1/memory[12][7] ), .C(n9352), .D(
        n9233), .Y(n4229) );
  AOI22X1 U4970 ( .A(n9905), .B(\U_0/U_1/U_1/memory[12][6] ), .C(
        \U_0/RCV_DATA [6]), .D(n9233), .Y(n4232) );
  AOI22X1 U4972 ( .A(n9905), .B(\U_0/U_1/U_1/memory[12][5] ), .C(n9348), .D(
        n9233), .Y(n4233) );
  AOI22X1 U4974 ( .A(n9905), .B(\U_0/U_1/U_1/memory[12][4] ), .C(n9346), .D(
        n9233), .Y(n4234) );
  AOI22X1 U4976 ( .A(n9905), .B(\U_0/U_1/U_1/memory[12][3] ), .C(n9344), .D(
        n9233), .Y(n4235) );
  AOI22X1 U4978 ( .A(n9905), .B(\U_0/U_1/U_1/memory[12][2] ), .C(n9342), .D(
        n9233), .Y(n4236) );
  AOI22X1 U4980 ( .A(n9905), .B(\U_0/U_1/U_1/memory[12][1] ), .C(n9340), .D(
        n9233), .Y(n4237) );
  AOI22X1 U4982 ( .A(n9905), .B(\U_0/U_1/U_1/memory[12][0] ), .C(n9338), .D(
        n9233), .Y(n4238) );
  AOI22X1 U4984 ( .A(n9896), .B(\U_0/U_1/U_1/memory[13][7] ), .C(
        \U_0/RCV_DATA [7]), .D(n9232), .Y(n4239) );
  AOI22X1 U4986 ( .A(n9896), .B(\U_0/U_1/U_1/memory[13][6] ), .C(
        \U_0/RCV_DATA [6]), .D(n9232), .Y(n4242) );
  AOI22X1 U4988 ( .A(n9896), .B(\U_0/U_1/U_1/memory[13][5] ), .C(
        \U_0/RCV_DATA [5]), .D(n9232), .Y(n4243) );
  AOI22X1 U4990 ( .A(n9896), .B(\U_0/U_1/U_1/memory[13][4] ), .C(n9346), .D(
        n9232), .Y(n4244) );
  AOI22X1 U4992 ( .A(n9896), .B(\U_0/U_1/U_1/memory[13][3] ), .C(n9344), .D(
        n9232), .Y(n4245) );
  AOI22X1 U4994 ( .A(n9896), .B(\U_0/U_1/U_1/memory[13][2] ), .C(
        \U_0/RCV_DATA [2]), .D(n9232), .Y(n4246) );
  AOI22X1 U4996 ( .A(n9896), .B(\U_0/U_1/U_1/memory[13][1] ), .C(
        \U_0/RCV_DATA [1]), .D(n9232), .Y(n4247) );
  AOI22X1 U4998 ( .A(n9896), .B(\U_0/U_1/U_1/memory[13][0] ), .C(n9338), .D(
        n9232), .Y(n4248) );
  AOI22X1 U5000 ( .A(n9887), .B(\U_0/U_1/U_1/memory[14][7] ), .C(n9352), .D(
        n9231), .Y(n4249) );
  AOI22X1 U5002 ( .A(n9887), .B(\U_0/U_1/U_1/memory[14][6] ), .C(
        \U_0/RCV_DATA [6]), .D(n9231), .Y(n4252) );
  AOI22X1 U5004 ( .A(n9887), .B(\U_0/U_1/U_1/memory[14][5] ), .C(n9348), .D(
        n9231), .Y(n4253) );
  AOI22X1 U5006 ( .A(n9887), .B(\U_0/U_1/U_1/memory[14][4] ), .C(n9346), .D(
        n9231), .Y(n4254) );
  AOI22X1 U5008 ( .A(n9887), .B(\U_0/U_1/U_1/memory[14][3] ), .C(n9344), .D(
        n9231), .Y(n4255) );
  AOI22X1 U5010 ( .A(n9887), .B(\U_0/U_1/U_1/memory[14][2] ), .C(n9342), .D(
        n9231), .Y(n4256) );
  AOI22X1 U5012 ( .A(n9887), .B(\U_0/U_1/U_1/memory[14][1] ), .C(n9340), .D(
        n9231), .Y(n4257) );
  AOI22X1 U5014 ( .A(n9887), .B(\U_0/U_1/U_1/memory[14][0] ), .C(n9338), .D(
        n9231), .Y(n4258) );
  AOI22X1 U5016 ( .A(n9878), .B(\U_0/U_1/U_1/memory[15][7] ), .C(
        \U_0/RCV_DATA [7]), .D(n9230), .Y(n4259) );
  AOI22X1 U5018 ( .A(n9878), .B(\U_0/U_1/U_1/memory[15][6] ), .C(n9350), .D(
        n9230), .Y(n4262) );
  AOI22X1 U5020 ( .A(n9878), .B(\U_0/U_1/U_1/memory[15][5] ), .C(
        \U_0/RCV_DATA [5]), .D(n9230), .Y(n4263) );
  AOI22X1 U5022 ( .A(n9878), .B(\U_0/U_1/U_1/memory[15][4] ), .C(
        \U_0/RCV_DATA [4]), .D(n9230), .Y(n4264) );
  AOI22X1 U5024 ( .A(n9878), .B(\U_0/U_1/U_1/memory[15][3] ), .C(
        \U_0/RCV_DATA [3]), .D(n9230), .Y(n4265) );
  AOI22X1 U5026 ( .A(n9878), .B(\U_0/U_1/U_1/memory[15][2] ), .C(
        \U_0/RCV_DATA [2]), .D(n9230), .Y(n4266) );
  AOI22X1 U5028 ( .A(n9878), .B(\U_0/U_1/U_1/memory[15][1] ), .C(
        \U_0/RCV_DATA [1]), .D(n9230), .Y(n4267) );
  AOI22X1 U5030 ( .A(n9878), .B(\U_0/U_1/U_1/memory[15][0] ), .C(
        \U_0/RCV_DATA [0]), .D(n9230), .Y(n4268) );
  OAI22X1 U5031 ( .A(n9229), .B(n11047), .C(n9351), .D(n9869), .Y(n8771) );
  OAI22X1 U5033 ( .A(n9229), .B(n11046), .C(n9349), .D(n9869), .Y(n8772) );
  OAI22X1 U5035 ( .A(n9229), .B(n11045), .C(n9347), .D(n9869), .Y(n8773) );
  OAI22X1 U5037 ( .A(n9229), .B(n11044), .C(n9345), .D(n9869), .Y(n8774) );
  OAI22X1 U5039 ( .A(n9229), .B(n11043), .C(n9343), .D(n9869), .Y(n8775) );
  OAI22X1 U5041 ( .A(n9229), .B(n11042), .C(n9341), .D(n9869), .Y(n8776) );
  OAI22X1 U5043 ( .A(n9229), .B(n11041), .C(n9339), .D(n9869), .Y(n8777) );
  OAI22X1 U5045 ( .A(n9229), .B(n11040), .C(n9337), .D(n9869), .Y(n8778) );
  OAI22X1 U5047 ( .A(n9228), .B(n11057), .C(n9351), .D(n9868), .Y(n8779) );
  OAI22X1 U5049 ( .A(n9228), .B(n11056), .C(n9349), .D(n9868), .Y(n8780) );
  OAI22X1 U5051 ( .A(n9228), .B(n11055), .C(n9347), .D(n9868), .Y(n8781) );
  OAI22X1 U5053 ( .A(n9228), .B(n11054), .C(n9345), .D(n9868), .Y(n8782) );
  OAI22X1 U5055 ( .A(n9228), .B(n11053), .C(n9343), .D(n9868), .Y(n8783) );
  OAI22X1 U5057 ( .A(n9228), .B(n11052), .C(n9341), .D(n9868), .Y(n8784) );
  OAI22X1 U5059 ( .A(n9228), .B(n11051), .C(n9339), .D(n9868), .Y(n8785) );
  OAI22X1 U5061 ( .A(n9228), .B(n11050), .C(n9337), .D(n9868), .Y(n8786) );
  OAI22X1 U5063 ( .A(n9227), .B(n11067), .C(n9351), .D(n9867), .Y(n8787) );
  OAI22X1 U5065 ( .A(n9227), .B(n11066), .C(n9349), .D(n9867), .Y(n8788) );
  OAI22X1 U5067 ( .A(n9227), .B(n11065), .C(n9347), .D(n9867), .Y(n8789) );
  OAI22X1 U5069 ( .A(n9227), .B(n11064), .C(n9345), .D(n9867), .Y(n8790) );
  OAI22X1 U5071 ( .A(n9227), .B(n11063), .C(n9343), .D(n9867), .Y(n8791) );
  OAI22X1 U5073 ( .A(n9227), .B(n11062), .C(n9341), .D(n9867), .Y(n8792) );
  OAI22X1 U5075 ( .A(n9227), .B(n11061), .C(n9339), .D(n9867), .Y(n8793) );
  OAI22X1 U5077 ( .A(n9227), .B(n11060), .C(n9337), .D(n9867), .Y(n8794) );
  OAI22X1 U5079 ( .A(n9226), .B(n11077), .C(n9341), .D(n9866), .Y(n8795) );
  OAI22X1 U5081 ( .A(n9226), .B(n11076), .C(n9339), .D(n9866), .Y(n8796) );
  OAI22X1 U5083 ( .A(n9226), .B(n11075), .C(n9337), .D(n9866), .Y(n8797) );
  OAI22X1 U5085 ( .A(n9226), .B(n11074), .C(n9351), .D(n9866), .Y(n8798) );
  OAI22X1 U5087 ( .A(n9226), .B(n11073), .C(n9349), .D(n9866), .Y(n8799) );
  OAI22X1 U5089 ( .A(n9226), .B(n11072), .C(n9347), .D(n9866), .Y(n8800) );
  OAI22X1 U5091 ( .A(n9226), .B(n11071), .C(n9345), .D(n9866), .Y(n8801) );
  OAI22X1 U5093 ( .A(n9226), .B(n11070), .C(n9343), .D(n9866), .Y(n8802) );
  AOI22X1 U5096 ( .A(n9865), .B(\U_0/U_1/U_1/memory[20][7] ), .C(n9352), .D(
        n9225), .Y(n4277) );
  AOI22X1 U5098 ( .A(n9865), .B(\U_0/U_1/U_1/memory[20][6] ), .C(n9350), .D(
        n9225), .Y(n4280) );
  AOI22X1 U5100 ( .A(n9865), .B(\U_0/U_1/U_1/memory[20][5] ), .C(n9348), .D(
        n9225), .Y(n4281) );
  AOI22X1 U5102 ( .A(n9865), .B(\U_0/U_1/U_1/memory[20][4] ), .C(
        \U_0/RCV_DATA [4]), .D(n9225), .Y(n4282) );
  AOI22X1 U5104 ( .A(n9865), .B(\U_0/U_1/U_1/memory[20][3] ), .C(
        \U_0/RCV_DATA [3]), .D(n9225), .Y(n4283) );
  AOI22X1 U5106 ( .A(n9865), .B(\U_0/U_1/U_1/memory[20][2] ), .C(n9342), .D(
        n9225), .Y(n4284) );
  AOI22X1 U5108 ( .A(n9865), .B(\U_0/U_1/U_1/memory[20][1] ), .C(n9340), .D(
        n9225), .Y(n4285) );
  AOI22X1 U5110 ( .A(n9865), .B(\U_0/U_1/U_1/memory[20][0] ), .C(
        \U_0/RCV_DATA [0]), .D(n9225), .Y(n4286) );
  AOI22X1 U5112 ( .A(n9856), .B(\U_0/U_1/U_1/memory[21][7] ), .C(
        \U_0/RCV_DATA [7]), .D(n9224), .Y(n4287) );
  AOI22X1 U5114 ( .A(n9856), .B(\U_0/U_1/U_1/memory[21][6] ), .C(n9350), .D(
        n9224), .Y(n4290) );
  AOI22X1 U5116 ( .A(n9856), .B(\U_0/U_1/U_1/memory[21][5] ), .C(
        \U_0/RCV_DATA [5]), .D(n9224), .Y(n4291) );
  AOI22X1 U5118 ( .A(n9856), .B(\U_0/U_1/U_1/memory[21][4] ), .C(
        \U_0/RCV_DATA [4]), .D(n9224), .Y(n4292) );
  AOI22X1 U5120 ( .A(n9856), .B(\U_0/U_1/U_1/memory[21][3] ), .C(
        \U_0/RCV_DATA [3]), .D(n9224), .Y(n4293) );
  AOI22X1 U5122 ( .A(n9856), .B(\U_0/U_1/U_1/memory[21][2] ), .C(
        \U_0/RCV_DATA [2]), .D(n9224), .Y(n4294) );
  AOI22X1 U5124 ( .A(n9856), .B(\U_0/U_1/U_1/memory[21][1] ), .C(
        \U_0/RCV_DATA [1]), .D(n9224), .Y(n4295) );
  AOI22X1 U5126 ( .A(n9856), .B(\U_0/U_1/U_1/memory[21][0] ), .C(
        \U_0/RCV_DATA [0]), .D(n9224), .Y(n4296) );
  AOI22X1 U5128 ( .A(n9847), .B(\U_0/U_1/U_1/memory[22][7] ), .C(n9352), .D(
        n9223), .Y(n4297) );
  AOI22X1 U5130 ( .A(n9847), .B(\U_0/U_1/U_1/memory[22][6] ), .C(n9350), .D(
        n9223), .Y(n4300) );
  AOI22X1 U5132 ( .A(n9847), .B(\U_0/U_1/U_1/memory[22][5] ), .C(n9348), .D(
        n9223), .Y(n4301) );
  AOI22X1 U5134 ( .A(n9847), .B(\U_0/U_1/U_1/memory[22][4] ), .C(
        \U_0/RCV_DATA [4]), .D(n9223), .Y(n4302) );
  AOI22X1 U5136 ( .A(n9847), .B(\U_0/U_1/U_1/memory[22][3] ), .C(
        \U_0/RCV_DATA [3]), .D(n9223), .Y(n4303) );
  AOI22X1 U5138 ( .A(n9847), .B(\U_0/U_1/U_1/memory[22][2] ), .C(n9342), .D(
        n9223), .Y(n4304) );
  AOI22X1 U5140 ( .A(n9847), .B(\U_0/U_1/U_1/memory[22][1] ), .C(n9340), .D(
        n9223), .Y(n4305) );
  AOI22X1 U5142 ( .A(n9847), .B(\U_0/U_1/U_1/memory[22][0] ), .C(
        \U_0/RCV_DATA [0]), .D(n9223), .Y(n4306) );
  AOI22X1 U5144 ( .A(n9838), .B(\U_0/U_1/U_1/memory[23][7] ), .C(
        \U_0/RCV_DATA [7]), .D(n9222), .Y(n4307) );
  AOI22X1 U5146 ( .A(n9838), .B(\U_0/U_1/U_1/memory[23][6] ), .C(n9350), .D(
        n9222), .Y(n4310) );
  AOI22X1 U5148 ( .A(n9838), .B(\U_0/U_1/U_1/memory[23][5] ), .C(
        \U_0/RCV_DATA [5]), .D(n9222), .Y(n4311) );
  AOI22X1 U5150 ( .A(n9838), .B(\U_0/U_1/U_1/memory[23][4] ), .C(
        \U_0/RCV_DATA [4]), .D(n9222), .Y(n4312) );
  AOI22X1 U5152 ( .A(n9838), .B(\U_0/U_1/U_1/memory[23][3] ), .C(
        \U_0/RCV_DATA [3]), .D(n9222), .Y(n4313) );
  AOI22X1 U5154 ( .A(n9838), .B(\U_0/U_1/U_1/memory[23][2] ), .C(
        \U_0/RCV_DATA [2]), .D(n9222), .Y(n4314) );
  AOI22X1 U5156 ( .A(n9838), .B(\U_0/U_1/U_1/memory[23][1] ), .C(
        \U_0/RCV_DATA [1]), .D(n9222), .Y(n4315) );
  AOI22X1 U5158 ( .A(n9838), .B(\U_0/U_1/U_1/memory[23][0] ), .C(
        \U_0/RCV_DATA [0]), .D(n9222), .Y(n4316) );
  AOI22X1 U5160 ( .A(n9829), .B(\U_0/U_1/U_1/memory[24][7] ), .C(n9352), .D(
        n9221), .Y(n4317) );
  AOI22X1 U5162 ( .A(n9829), .B(\U_0/U_1/U_1/memory[24][6] ), .C(n9350), .D(
        n9221), .Y(n4320) );
  AOI22X1 U5164 ( .A(n9829), .B(\U_0/U_1/U_1/memory[24][5] ), .C(n9348), .D(
        n9221), .Y(n4321) );
  AOI22X1 U5166 ( .A(n9829), .B(\U_0/U_1/U_1/memory[24][4] ), .C(
        \U_0/RCV_DATA [4]), .D(n9221), .Y(n4322) );
  AOI22X1 U5168 ( .A(n9829), .B(\U_0/U_1/U_1/memory[24][3] ), .C(
        \U_0/RCV_DATA [3]), .D(n9221), .Y(n4323) );
  AOI22X1 U5170 ( .A(n9829), .B(\U_0/U_1/U_1/memory[24][2] ), .C(n9342), .D(
        n9221), .Y(n4324) );
  AOI22X1 U5172 ( .A(n9829), .B(\U_0/U_1/U_1/memory[24][1] ), .C(n9340), .D(
        n9221), .Y(n4325) );
  AOI22X1 U5174 ( .A(n9829), .B(\U_0/U_1/U_1/memory[24][0] ), .C(
        \U_0/RCV_DATA [0]), .D(n9221), .Y(n4326) );
  AOI22X1 U5176 ( .A(n9820), .B(\U_0/U_1/U_1/memory[25][7] ), .C(
        \U_0/RCV_DATA [7]), .D(n9220), .Y(n4327) );
  AOI22X1 U5178 ( .A(n9820), .B(\U_0/U_1/U_1/memory[25][6] ), .C(n9350), .D(
        n9220), .Y(n4330) );
  AOI22X1 U5180 ( .A(n9820), .B(\U_0/U_1/U_1/memory[25][5] ), .C(
        \U_0/RCV_DATA [5]), .D(n9220), .Y(n4331) );
  AOI22X1 U5182 ( .A(n9820), .B(\U_0/U_1/U_1/memory[25][4] ), .C(
        \U_0/RCV_DATA [4]), .D(n9220), .Y(n4332) );
  AOI22X1 U5184 ( .A(n9820), .B(\U_0/U_1/U_1/memory[25][3] ), .C(
        \U_0/RCV_DATA [3]), .D(n9220), .Y(n4333) );
  AOI22X1 U5186 ( .A(n9820), .B(\U_0/U_1/U_1/memory[25][2] ), .C(
        \U_0/RCV_DATA [2]), .D(n9220), .Y(n4334) );
  AOI22X1 U5188 ( .A(n9820), .B(\U_0/U_1/U_1/memory[25][1] ), .C(
        \U_0/RCV_DATA [1]), .D(n9220), .Y(n4335) );
  AOI22X1 U5190 ( .A(n9820), .B(\U_0/U_1/U_1/memory[25][0] ), .C(
        \U_0/RCV_DATA [0]), .D(n9220), .Y(n4336) );
  AOI22X1 U5192 ( .A(n9811), .B(\U_0/U_1/U_1/memory[26][7] ), .C(n9352), .D(
        n9219), .Y(n4337) );
  AOI22X1 U5194 ( .A(n9811), .B(\U_0/U_1/U_1/memory[26][6] ), .C(n9350), .D(
        n9219), .Y(n4340) );
  AOI22X1 U5196 ( .A(n9811), .B(\U_0/U_1/U_1/memory[26][5] ), .C(n9348), .D(
        n9219), .Y(n4341) );
  AOI22X1 U5198 ( .A(n9811), .B(\U_0/U_1/U_1/memory[26][4] ), .C(n9346), .D(
        n9219), .Y(n4342) );
  AOI22X1 U5200 ( .A(n9811), .B(\U_0/U_1/U_1/memory[26][3] ), .C(n9344), .D(
        n9219), .Y(n4343) );
  AOI22X1 U5202 ( .A(n9811), .B(\U_0/U_1/U_1/memory[26][2] ), .C(n9342), .D(
        n9219), .Y(n4344) );
  AOI22X1 U5204 ( .A(n9811), .B(\U_0/U_1/U_1/memory[26][1] ), .C(n9340), .D(
        n9219), .Y(n4345) );
  AOI22X1 U5206 ( .A(n9811), .B(\U_0/U_1/U_1/memory[26][0] ), .C(n9338), .D(
        n9219), .Y(n4346) );
  AOI22X1 U5208 ( .A(n9802), .B(\U_0/U_1/U_1/memory[27][7] ), .C(n9352), .D(
        n9218), .Y(n4347) );
  AOI22X1 U5210 ( .A(n9802), .B(\U_0/U_1/U_1/memory[27][6] ), .C(n9350), .D(
        n9218), .Y(n4350) );
  AOI22X1 U5212 ( .A(n9802), .B(\U_0/U_1/U_1/memory[27][5] ), .C(n9348), .D(
        n9218), .Y(n4351) );
  AOI22X1 U5214 ( .A(n9802), .B(\U_0/U_1/U_1/memory[27][4] ), .C(n9346), .D(
        n9218), .Y(n4352) );
  AOI22X1 U5216 ( .A(n9802), .B(\U_0/U_1/U_1/memory[27][3] ), .C(n9344), .D(
        n9218), .Y(n4353) );
  AOI22X1 U5218 ( .A(n9802), .B(\U_0/U_1/U_1/memory[27][2] ), .C(n9342), .D(
        n9218), .Y(n4354) );
  AOI22X1 U5220 ( .A(n9802), .B(\U_0/U_1/U_1/memory[27][1] ), .C(n9340), .D(
        n9218), .Y(n4355) );
  AOI22X1 U5222 ( .A(n9802), .B(\U_0/U_1/U_1/memory[27][0] ), .C(n9338), .D(
        n9218), .Y(n4356) );
  OAI22X1 U5223 ( .A(n9217), .B(n11007), .C(n9351), .D(n9793), .Y(n8867) );
  OAI22X1 U5225 ( .A(n9217), .B(n11006), .C(n9349), .D(n9793), .Y(n8868) );
  OAI22X1 U5227 ( .A(n9217), .B(n11005), .C(n9347), .D(n9793), .Y(n8869) );
  OAI22X1 U5229 ( .A(n9217), .B(n11004), .C(n9345), .D(n9793), .Y(n8870) );
  OAI22X1 U5231 ( .A(n9217), .B(n11003), .C(n9343), .D(n9793), .Y(n8871) );
  OAI22X1 U5233 ( .A(n9217), .B(n11002), .C(n9341), .D(n9793), .Y(n8872) );
  OAI22X1 U5235 ( .A(n9217), .B(n11001), .C(n9339), .D(n9793), .Y(n8873) );
  OAI22X1 U5237 ( .A(n9217), .B(n11000), .C(n9337), .D(n9793), .Y(n8874) );
  OAI22X1 U5239 ( .A(n9216), .B(n11017), .C(n9351), .D(n9792), .Y(n8875) );
  OAI22X1 U5241 ( .A(n9216), .B(n11016), .C(n9349), .D(n9792), .Y(n8876) );
  OAI22X1 U5243 ( .A(n9216), .B(n11015), .C(n9347), .D(n9792), .Y(n8877) );
  OAI22X1 U5245 ( .A(n9216), .B(n11014), .C(n9345), .D(n9792), .Y(n8878) );
  OAI22X1 U5247 ( .A(n9216), .B(n11013), .C(n9343), .D(n9792), .Y(n8879) );
  OAI22X1 U5249 ( .A(n9216), .B(n11012), .C(n9341), .D(n9792), .Y(n8880) );
  OAI22X1 U5251 ( .A(n9216), .B(n11011), .C(n9339), .D(n9792), .Y(n8881) );
  OAI22X1 U5253 ( .A(n9216), .B(n11010), .C(n9337), .D(n9792), .Y(n8882) );
  OAI22X1 U5255 ( .A(n9215), .B(n11027), .C(n9351), .D(n9791), .Y(n8883) );
  OAI22X1 U5257 ( .A(n9215), .B(n11026), .C(n9349), .D(n9791), .Y(n8884) );
  OAI22X1 U5259 ( .A(n9215), .B(n11025), .C(n9347), .D(n9791), .Y(n8885) );
  OAI22X1 U5261 ( .A(n9215), .B(n11024), .C(n9345), .D(n9791), .Y(n8886) );
  OAI22X1 U5263 ( .A(n9215), .B(n11023), .C(n9343), .D(n9791), .Y(n8887) );
  OAI22X1 U5265 ( .A(n9215), .B(n11022), .C(n9341), .D(n9791), .Y(n8888) );
  OAI22X1 U5267 ( .A(n9215), .B(n11021), .C(n9339), .D(n9791), .Y(n8889) );
  OAI22X1 U5269 ( .A(n9215), .B(n11020), .C(n9337), .D(n9791), .Y(n8890) );
  OAI22X1 U5271 ( .A(n9214), .B(n11037), .C(n9351), .D(n9790), .Y(n8891) );
  OAI22X1 U5273 ( .A(n9214), .B(n11036), .C(n9349), .D(n9790), .Y(n8892) );
  OAI22X1 U5275 ( .A(n9214), .B(n11035), .C(n9347), .D(n9790), .Y(n8893) );
  OAI22X1 U5277 ( .A(n9214), .B(n11034), .C(n9345), .D(n9790), .Y(n8894) );
  OAI22X1 U5279 ( .A(n9214), .B(n11033), .C(n9343), .D(n9790), .Y(n8895) );
  OAI22X1 U5281 ( .A(n9214), .B(n11032), .C(n9341), .D(n9790), .Y(n8896) );
  OAI22X1 U5283 ( .A(n9214), .B(n11031), .C(n9339), .D(n9790), .Y(n8897) );
  OAI22X1 U5285 ( .A(n9214), .B(n11030), .C(n9337), .D(n9790), .Y(n8898) );
  AOI22X1 U5288 ( .A(n4366), .B(n10805), .C(\U_0/U_1/U_1/opcode[0][1] ), .D(
        n9742), .Y(n4365) );
  AOI22X1 U5290 ( .A(n9181), .B(n4366), .C(\U_0/U_1/U_1/opcode[0][0] ), .D(
        n9742), .Y(n4369) );
  OAI21X1 U5292 ( .A(n4371), .B(n4372), .C(n9949), .Y(n4366) );
  NOR2X1 U5294 ( .A(n4373), .B(n4374), .Y(n4165) );
  AOI22X1 U5296 ( .A(n4376), .B(n10805), .C(\U_0/U_1/U_1/opcode[1][1] ), .D(
        n9739), .Y(n4375) );
  AOI22X1 U5298 ( .A(n9181), .B(n4376), .C(\U_0/U_1/U_1/opcode[1][0] ), .D(
        n9739), .Y(n4378) );
  OAI21X1 U5300 ( .A(n4228), .B(n4372), .C(n9940), .Y(n4376) );
  NOR2X1 U5302 ( .A(n4379), .B(n4373), .Y(n4175) );
  AOI22X1 U5304 ( .A(n4381), .B(n10805), .C(\U_0/U_1/U_1/opcode[2][1] ), .D(
        n9736), .Y(n4380) );
  AOI22X1 U5306 ( .A(n9181), .B(n4381), .C(\U_0/U_1/U_1/opcode[2][0] ), .D(
        n9736), .Y(n4383) );
  OAI21X1 U5308 ( .A(n4384), .B(n4372), .C(n9931), .Y(n4381) );
  NOR2X1 U5310 ( .A(n4371), .B(n4373), .Y(n4185) );
  AOI22X1 U5312 ( .A(n4386), .B(n10805), .C(\U_0/U_1/U_1/opcode[3][1] ), .D(
        n9733), .Y(n4385) );
  AOI22X1 U5314 ( .A(n9181), .B(n4386), .C(\U_0/U_1/U_1/opcode[3][0] ), .D(
        n9733), .Y(n4388) );
  OAI21X1 U5316 ( .A(n4389), .B(n4372), .C(n9922), .Y(n4386) );
  NOR2X1 U5318 ( .A(n4228), .B(n4373), .Y(n4195) );
  OAI22X1 U5319 ( .A(n9730), .B(n9193), .C(n10919), .D(n4392), .Y(n8907) );
  OAI22X1 U5321 ( .A(n9210), .B(n9730), .C(n10918), .D(n4392), .Y(n8908) );
  OAI21X1 U5324 ( .A(n4394), .B(n4372), .C(n9913), .Y(n4392) );
  NOR2X1 U5326 ( .A(n4384), .B(n4373), .Y(n4203) );
  OAI22X1 U5327 ( .A(n9729), .B(n9194), .C(n10929), .D(n4396), .Y(n8909) );
  OAI22X1 U5329 ( .A(n9210), .B(n9729), .C(n10928), .D(n4396), .Y(n8910) );
  OAI21X1 U5332 ( .A(n4397), .B(n4372), .C(n9912), .Y(n4396) );
  NOR2X1 U5334 ( .A(n4389), .B(n4373), .Y(n4213) );
  OAI22X1 U5335 ( .A(n9789), .B(n9193), .C(n10957), .D(n4399), .Y(n8911) );
  OAI22X1 U5337 ( .A(n9210), .B(n9789), .C(n10956), .D(n4399), .Y(n8912) );
  OAI21X1 U5340 ( .A(n4374), .B(n4400), .C(n9911), .Y(n4399) );
  NOR2X1 U5342 ( .A(n4394), .B(n4373), .Y(n4215) );
  OAI22X1 U5343 ( .A(n9788), .B(n9195), .C(n10959), .D(n4402), .Y(n8913) );
  OAI22X1 U5345 ( .A(n9210), .B(n9788), .C(n10958), .D(n4402), .Y(n8914) );
  OAI21X1 U5348 ( .A(n4379), .B(n4400), .C(n9910), .Y(n4402) );
  NOR2X1 U5350 ( .A(n4397), .B(n4373), .Y(n4217) );
  NAND3X1 U5351 ( .A(n9325), .B(n9327), .C(n4405), .Y(n4373) );
  OAI22X1 U5352 ( .A(n9787), .B(n9193), .C(n10969), .D(n4407), .Y(n8915) );
  OAI22X1 U5354 ( .A(n9210), .B(n9787), .C(n10968), .D(n4407), .Y(n8916) );
  OAI21X1 U5357 ( .A(n4371), .B(n4400), .C(n9908), .Y(n4407) );
  NOR2X1 U5359 ( .A(n4227), .B(n4374), .Y(n4219) );
  OAI22X1 U5360 ( .A(n9786), .B(n9195), .C(n10979), .D(n4409), .Y(n8917) );
  OAI22X1 U5362 ( .A(n9210), .B(n9786), .C(n10978), .D(n4409), .Y(n8918) );
  OAI21X1 U5365 ( .A(n4228), .B(n4400), .C(n9907), .Y(n4409) );
  NOR2X1 U5367 ( .A(n4227), .B(n4379), .Y(n4221) );
  OAI22X1 U5368 ( .A(n9785), .B(n9194), .C(n10989), .D(n4411), .Y(n8919) );
  OAI22X1 U5370 ( .A(n9210), .B(n9785), .C(n10988), .D(n4411), .Y(n8920) );
  OAI21X1 U5373 ( .A(n4384), .B(n4400), .C(n9906), .Y(n4411) );
  NOR2X1 U5375 ( .A(n4227), .B(n4371), .Y(n4223) );
  OAI22X1 U5376 ( .A(n9950), .B(n10955), .C(n9210), .D(n4413), .Y(n8921) );
  OAI22X1 U5378 ( .A(n9950), .B(n10954), .C(n9194), .D(n4413), .Y(n8922) );
  NAND3X1 U5381 ( .A(n4414), .B(n9326), .C(n4415), .Y(n4413) );
  AOI21X1 U5382 ( .A(n4228), .B(n9195), .C(n4416), .Y(n4415) );
  NAND2X1 U5383 ( .A(n9510), .B(n9327), .Y(n4416) );
  AOI21X1 U5384 ( .A(n10805), .B(n4389), .C(n4417), .Y(n4414) );
  AOI22X1 U5386 ( .A(n4419), .B(n10805), .C(\U_0/U_1/U_1/opcode[12][1] ), .D(
        n9784), .Y(n4418) );
  AOI22X1 U5388 ( .A(n9181), .B(n4419), .C(\U_0/U_1/U_1/opcode[12][0] ), .D(
        n9784), .Y(n4421) );
  OAI21X1 U5390 ( .A(n4394), .B(n4400), .C(n9905), .Y(n4419) );
  NOR2X1 U5392 ( .A(n4227), .B(n4384), .Y(n4231) );
  AOI22X1 U5394 ( .A(n4423), .B(n10805), .C(\U_0/U_1/U_1/opcode[13][1] ), .D(
        n9781), .Y(n4422) );
  AOI22X1 U5396 ( .A(n9181), .B(n4423), .C(\U_0/U_1/U_1/opcode[13][0] ), .D(
        n9781), .Y(n4425) );
  OAI21X1 U5398 ( .A(n4397), .B(n4400), .C(n9896), .Y(n4423) );
  NOR2X1 U5400 ( .A(n4227), .B(n4389), .Y(n4241) );
  NAND3X1 U5401 ( .A(n9326), .B(n9327), .C(n4426), .Y(n4400) );
  AOI22X1 U5403 ( .A(n4428), .B(n10805), .C(\U_0/U_1/U_1/opcode[14][1] ), .D(
        n9778), .Y(n4427) );
  AOI22X1 U5405 ( .A(n9181), .B(n4428), .C(\U_0/U_1/U_1/opcode[14][0] ), .D(
        n9778), .Y(n4430) );
  OAI21X1 U5407 ( .A(n4374), .B(n4431), .C(n9887), .Y(n4428) );
  NOR2X1 U5409 ( .A(n4227), .B(n4394), .Y(n4251) );
  AOI22X1 U5411 ( .A(n4433), .B(n10805), .C(\U_0/U_1/U_1/opcode[15][1] ), .D(
        n9775), .Y(n4432) );
  AOI22X1 U5413 ( .A(n9181), .B(n4433), .C(\U_0/U_1/U_1/opcode[15][0] ), .D(
        n9775), .Y(n4435) );
  OAI21X1 U5415 ( .A(n4379), .B(n4431), .C(n9878), .Y(n4433) );
  NOR2X1 U5417 ( .A(n4227), .B(n4397), .Y(n4261) );
  NAND3X1 U5418 ( .A(n4405), .B(n9327), .C(n9326), .Y(n4227) );
  OAI22X1 U5419 ( .A(n9772), .B(n9195), .C(n11039), .D(n4437), .Y(n8931) );
  OAI22X1 U5421 ( .A(n9210), .B(n9772), .C(n11038), .D(n4437), .Y(n8932) );
  OAI21X1 U5424 ( .A(n4371), .B(n4431), .C(n9869), .Y(n4437) );
  NOR2X1 U5426 ( .A(n4438), .B(n4374), .Y(n4269) );
  OAI22X1 U5427 ( .A(n9771), .B(n9194), .C(n11049), .D(n4440), .Y(n8933) );
  OAI22X1 U5429 ( .A(n9210), .B(n9771), .C(n11048), .D(n4440), .Y(n8934) );
  OAI21X1 U5432 ( .A(n4228), .B(n4431), .C(n9868), .Y(n4440) );
  NOR2X1 U5434 ( .A(n4438), .B(n4379), .Y(n4271) );
  OAI22X1 U5435 ( .A(n9770), .B(n9193), .C(n11059), .D(n4442), .Y(n8935) );
  OAI22X1 U5437 ( .A(n9210), .B(n9770), .C(n11058), .D(n4442), .Y(n8936) );
  OAI21X1 U5440 ( .A(n4384), .B(n4431), .C(n9867), .Y(n4442) );
  NOR2X1 U5442 ( .A(n4438), .B(n4371), .Y(n4273) );
  OAI22X1 U5443 ( .A(n9769), .B(n9194), .C(n11069), .D(n4444), .Y(n8937) );
  OAI22X1 U5445 ( .A(n9210), .B(n9769), .C(n11068), .D(n4444), .Y(n8938) );
  OAI21X1 U5448 ( .A(n4389), .B(n4431), .C(n9866), .Y(n4444) );
  NOR2X1 U5450 ( .A(n4438), .B(n4228), .Y(n4275) );
  AOI22X1 U5452 ( .A(n4446), .B(n10805), .C(\U_0/U_1/U_1/opcode[20][1] ), .D(
        n9768), .Y(n4445) );
  AOI22X1 U5454 ( .A(n9181), .B(n4446), .C(\U_0/U_1/U_1/opcode[20][0] ), .D(
        n9768), .Y(n4448) );
  OAI21X1 U5456 ( .A(n4394), .B(n4431), .C(n9865), .Y(n4446) );
  NOR2X1 U5458 ( .A(n4438), .B(n4384), .Y(n4279) );
  AOI22X1 U5460 ( .A(n4450), .B(n10805), .C(\U_0/U_1/U_1/opcode[21][1] ), .D(
        n9765), .Y(n4449) );
  AOI22X1 U5462 ( .A(n9181), .B(n4450), .C(\U_0/U_1/U_1/opcode[21][0] ), .D(
        n9765), .Y(n4452) );
  OAI21X1 U5464 ( .A(n4397), .B(n4431), .C(n9856), .Y(n4450) );
  NOR2X1 U5466 ( .A(n4438), .B(n4389), .Y(n4289) );
  NAND3X1 U5467 ( .A(\U_0/U_1/U_1/writeptr[4] ), .B(n9325), .C(n4426), .Y(
        n4431) );
  AOI22X1 U5469 ( .A(n4454), .B(n10805), .C(\U_0/U_1/U_1/opcode[22][1] ), .D(
        n9762), .Y(n4453) );
  AOI22X1 U5471 ( .A(n9181), .B(n4454), .C(\U_0/U_1/U_1/opcode[22][0] ), .D(
        n9762), .Y(n4456) );
  OAI21X1 U5473 ( .A(n4374), .B(n4457), .C(n9847), .Y(n4454) );
  NOR2X1 U5475 ( .A(n4438), .B(n4394), .Y(n4299) );
  AOI22X1 U5477 ( .A(n4459), .B(n10805), .C(\U_0/U_1/U_1/opcode[23][1] ), .D(
        n9759), .Y(n4458) );
  AOI22X1 U5479 ( .A(n9181), .B(n4459), .C(\U_0/U_1/U_1/opcode[23][0] ), .D(
        n9759), .Y(n4461) );
  OAI21X1 U5481 ( .A(n4379), .B(n4457), .C(n9838), .Y(n4459) );
  NOR2X1 U5483 ( .A(n4438), .B(n4397), .Y(n4309) );
  NAND3X1 U5484 ( .A(n4405), .B(n9325), .C(n9328), .Y(n4438) );
  AOI22X1 U5486 ( .A(n4463), .B(n10805), .C(\U_0/U_1/U_1/opcode[24][1] ), .D(
        n9756), .Y(n4462) );
  AOI22X1 U5488 ( .A(n9181), .B(n4463), .C(\U_0/U_1/U_1/opcode[24][0] ), .D(
        n9756), .Y(n4465) );
  OAI21X1 U5490 ( .A(n4371), .B(n4457), .C(n9829), .Y(n4463) );
  NOR2X1 U5492 ( .A(n4466), .B(n4374), .Y(n4319) );
  AOI22X1 U5494 ( .A(n4468), .B(n10805), .C(\U_0/U_1/U_1/opcode[25][1] ), .D(
        n9753), .Y(n4467) );
  AOI22X1 U5496 ( .A(n9181), .B(n4468), .C(\U_0/U_1/U_1/opcode[25][0] ), .D(
        n9753), .Y(n4470) );
  OAI21X1 U5498 ( .A(n4228), .B(n4457), .C(n9820), .Y(n4468) );
  NOR2X1 U5500 ( .A(n4466), .B(n4379), .Y(n4329) );
  AOI22X1 U5502 ( .A(n4472), .B(n10805), .C(\U_0/U_1/U_1/opcode[26][1] ), .D(
        n9750), .Y(n4471) );
  AOI22X1 U5504 ( .A(n9181), .B(n4472), .C(\U_0/U_1/U_1/opcode[26][0] ), .D(
        n9750), .Y(n4474) );
  OAI21X1 U5506 ( .A(n4384), .B(n4457), .C(n9811), .Y(n4472) );
  NOR2X1 U5508 ( .A(n4466), .B(n4371), .Y(n4339) );
  NAND3X1 U5509 ( .A(n10917), .B(n9321), .C(n9324), .Y(n4371) );
  AOI22X1 U5511 ( .A(n4478), .B(n10805), .C(\U_0/U_1/U_1/opcode[27][1] ), .D(
        n9747), .Y(n4477) );
  AOI22X1 U5513 ( .A(n9181), .B(n4478), .C(\U_0/U_1/U_1/opcode[27][0] ), .D(
        n9747), .Y(n4480) );
  OAI21X1 U5515 ( .A(n4389), .B(n4457), .C(n9802), .Y(n4478) );
  NOR2X1 U5517 ( .A(n4466), .B(n4228), .Y(n4349) );
  NAND3X1 U5518 ( .A(\U_0/U_1/U_1/writeptr[0] ), .B(n9321), .C(n9324), .Y(
        n4228) );
  OAI22X1 U5519 ( .A(n9744), .B(n9193), .C(n10999), .D(n4482), .Y(n8955) );
  OAI22X1 U5521 ( .A(n9210), .B(n9744), .C(n10998), .D(n4482), .Y(n8956) );
  OAI21X1 U5524 ( .A(n4394), .B(n4457), .C(n9793), .Y(n4482) );
  NOR2X1 U5526 ( .A(n4466), .B(n4384), .Y(n4357) );
  NAND3X1 U5527 ( .A(n10917), .B(n9323), .C(\U_0/U_1/U_1/writeptr[2] ), .Y(
        n4384) );
  OAI22X1 U5528 ( .A(n9743), .B(n9195), .C(n11009), .D(n4485), .Y(n8957) );
  OAI22X1 U5530 ( .A(n9210), .B(n9743), .C(n11008), .D(n4485), .Y(n8958) );
  OAI21X1 U5533 ( .A(n4397), .B(n4457), .C(n9792), .Y(n4485) );
  NOR2X1 U5535 ( .A(n4466), .B(n4389), .Y(n4359) );
  NAND3X1 U5536 ( .A(\U_0/U_1/U_1/writeptr[0] ), .B(n9323), .C(n9322), .Y(
        n4389) );
  NAND3X1 U5537 ( .A(\U_0/U_1/U_1/writeptr[4] ), .B(n9326), .C(n4426), .Y(
        n4457) );
  OAI22X1 U5538 ( .A(n9728), .B(n9193), .C(n11019), .D(n4487), .Y(n8959) );
  OAI22X1 U5540 ( .A(n9210), .B(n9728), .C(n11018), .D(n4487), .Y(n8960) );
  OAI21X1 U5543 ( .A(n4374), .B(n4372), .C(n9791), .Y(n4487) );
  NOR2X1 U5545 ( .A(n4466), .B(n4394), .Y(n4361) );
  NAND3X1 U5546 ( .A(n9324), .B(n10917), .C(\U_0/U_1/U_1/writeptr[2] ), .Y(
        n4394) );
  NAND3X1 U5547 ( .A(n9323), .B(n9321), .C(n10917), .Y(n4374) );
  OAI22X1 U5548 ( .A(n9727), .B(n9195), .C(n11029), .D(n4489), .Y(n8961) );
  OAI22X1 U5550 ( .A(n9210), .B(n9727), .C(n11028), .D(n4489), .Y(n8962) );
  OAI21X1 U5553 ( .A(n4379), .B(n4372), .C(n9790), .Y(n4489) );
  NOR2X1 U5555 ( .A(n4466), .B(n4397), .Y(n4363) );
  NAND3X1 U5556 ( .A(n9324), .B(\U_0/U_1/U_1/writeptr[0] ), .C(
        \U_0/U_1/U_1/writeptr[2] ), .Y(n4397) );
  NAND3X1 U5557 ( .A(n9326), .B(n4405), .C(n9328), .Y(n4466) );
  NAND3X1 U5559 ( .A(n9325), .B(n9327), .C(n4426), .Y(n4372) );
  NAND3X1 U5561 ( .A(n9323), .B(n9321), .C(\U_0/U_1/U_1/writeptr[0] ), .Y(
        n4379) );
  OAI21X1 U5562 ( .A(n10793), .B(n9325), .C(n4493), .Y(n8963) );
  AOI22X1 U5563 ( .A(\U_0/U_1/U_1/N50 ), .B(n4490), .C(\U_0/U_1/U_1/N45 ), .D(
        n4491), .Y(n4493) );
  OAI21X1 U5565 ( .A(n10793), .B(n9321), .C(n4494), .Y(n8964) );
  AOI22X1 U5566 ( .A(\U_0/U_1/U_1/N49 ), .B(n4490), .C(\U_0/U_1/U_1/N44 ), .D(
        n4491), .Y(n4494) );
  OAI21X1 U5568 ( .A(n10793), .B(n9323), .C(n4495), .Y(n8965) );
  AOI22X1 U5569 ( .A(\U_0/U_1/U_1/N48 ), .B(n4490), .C(\U_0/U_1/U_1/N43 ), .D(
        n4491), .Y(n4495) );
  OAI21X1 U5571 ( .A(n10793), .B(n10917), .C(n4496), .Y(n8966) );
  AOI22X1 U5572 ( .A(n10917), .B(n4490), .C(n10917), .D(n4491), .Y(n4496) );
  OAI21X1 U5574 ( .A(n10793), .B(n9327), .C(n4497), .Y(n8967) );
  AOI22X1 U5575 ( .A(\U_0/U_1/U_1/N51 ), .B(n4490), .C(\U_0/U_1/U_1/N46 ), .D(
        n4491), .Y(n4497) );
  NOR2X1 U5576 ( .A(n4417), .B(n9194), .Y(n4491) );
  NOR2X1 U5577 ( .A(n4417), .B(n10805), .Y(n4490) );
  NAND2X1 U5580 ( .A(\U_0/U_1/U_1/N36 ), .B(n9418), .Y(n4417) );
  OAI21X1 U5581 ( .A(n11114), .B(n3402), .C(n4499), .Y(n8968) );
  AOI22X1 U5582 ( .A(\U_0/U_3/U_3/N84 ), .B(n3404), .C(\U_0/U_3/U_3/N59 ), .D(
        n3405), .Y(n4499) );
  OAI21X1 U5584 ( .A(n4501), .B(n519), .C(n4502), .Y(n4500) );
  NOR2X1 U5585 ( .A(n10896), .B(n10892), .Y(n4502) );
  OAI21X1 U5586 ( .A(n4501), .B(n522), .C(n4505), .Y(n3404) );
  OAI21X1 U5587 ( .A(n10894), .B(n11093), .C(n10902), .Y(n4505) );
  NAND2X1 U5588 ( .A(n10896), .B(n10871), .Y(n3402) );
  OAI21X1 U5589 ( .A(RST), .B(n9713), .C(n4511), .Y(n8969) );
  NAND2X1 U5590 ( .A(CRCE_H), .B(RST), .Y(n4511) );
  OAI22X1 U5591 ( .A(n9531), .B(n10867), .C(RST), .D(n9713), .Y(n8970) );
  OAI21X1 U5593 ( .A(n9714), .B(n10867), .C(n4515), .Y(n4513) );
  NAND3X1 U5594 ( .A(n10805), .B(n10818), .C(n4517), .Y(n4515) );
  OAI21X1 U5596 ( .A(n9417), .B(n10819), .C(n4520), .Y(n8971) );
  NAND2X1 U5597 ( .A(\U_0/U_2/rx_CHECK_CRC [15]), .B(n9417), .Y(n4520) );
  OAI21X1 U5598 ( .A(n9417), .B(n10863), .C(n4522), .Y(n8972) );
  NAND2X1 U5599 ( .A(\U_0/U_2/rx_CHECK_CRC [14]), .B(n9417), .Y(n4522) );
  OAI21X1 U5600 ( .A(n9417), .B(n10862), .C(n4524), .Y(n8973) );
  NAND2X1 U5601 ( .A(\U_0/U_2/rx_CHECK_CRC [13]), .B(n9417), .Y(n4524) );
  OAI21X1 U5602 ( .A(n9417), .B(n10861), .C(n4526), .Y(n8974) );
  NAND2X1 U5603 ( .A(\U_0/U_2/rx_CHECK_CRC [12]), .B(n9417), .Y(n4526) );
  OAI21X1 U5604 ( .A(n9417), .B(n10860), .C(n4528), .Y(n8975) );
  NAND2X1 U5605 ( .A(\U_0/U_2/rx_CHECK_CRC [11]), .B(n9417), .Y(n4528) );
  OAI21X1 U5606 ( .A(n9417), .B(n10859), .C(n4530), .Y(n8976) );
  NAND2X1 U5607 ( .A(\U_0/U_2/rx_CHECK_CRC [10]), .B(n9417), .Y(n4530) );
  OAI21X1 U5608 ( .A(n9417), .B(n9599), .C(n4532), .Y(n8977) );
  NAND2X1 U5609 ( .A(\U_0/U_2/rx_CHECK_CRC [9]), .B(n9417), .Y(n4532) );
  OAI21X1 U5610 ( .A(n9417), .B(n10858), .C(n4534), .Y(n8978) );
  NAND2X1 U5611 ( .A(\U_0/U_2/rx_CHECK_CRC [8]), .B(n9417), .Y(n4534) );
  OAI22X1 U5612 ( .A(n10819), .B(n9418), .C(n9417), .D(n9351), .Y(n8979) );
  OAI22X1 U5614 ( .A(n9419), .B(n10863), .C(n9417), .D(n9349), .Y(n8980) );
  OAI22X1 U5616 ( .A(n9418), .B(n10862), .C(n9417), .D(n9347), .Y(n8981) );
  OAI22X1 U5618 ( .A(n9419), .B(n10861), .C(n9417), .D(n9345), .Y(n8982) );
  OAI22X1 U5620 ( .A(n9419), .B(n10860), .C(n9417), .D(n9343), .Y(n8983) );
  OAI22X1 U5622 ( .A(n9420), .B(n10859), .C(n9417), .D(n9341), .Y(n8984) );
  OAI22X1 U5624 ( .A(n9420), .B(n9599), .C(n9417), .D(n9339), .Y(n8985) );
  OAI22X1 U5626 ( .A(n9418), .B(n10858), .C(n9417), .D(n9337), .Y(n8986) );
  OAI21X1 U5630 ( .A(n9380), .B(n10846), .C(n4538), .Y(n8987) );
  NAND2X1 U5631 ( .A(\U_0/U_2/RX_CRC [14]), .B(n9382), .Y(n4538) );
  OAI22X1 U5632 ( .A(n9379), .B(n10845), .C(n9213), .D(n10846), .Y(n8988) );
  OAI22X1 U5634 ( .A(n9211), .B(n10843), .C(n10845), .D(n9212), .Y(n8989) );
  OAI21X1 U5635 ( .A(n9380), .B(n10849), .C(n4545), .Y(n8990) );
  NAND2X1 U5636 ( .A(\U_0/U_2/RX_CRC [13]), .B(n9382), .Y(n4545) );
  OAI22X1 U5637 ( .A(n9379), .B(n10842), .C(n9213), .D(n10849), .Y(n8991) );
  OAI22X1 U5639 ( .A(n9211), .B(n10840), .C(n9212), .D(n10842), .Y(n8992) );
  OAI21X1 U5641 ( .A(n9380), .B(n10839), .C(n4549), .Y(n8993) );
  NAND2X1 U5642 ( .A(\U_0/U_2/RX_CRC [12]), .B(n9382), .Y(n4549) );
  OAI22X1 U5643 ( .A(n9379), .B(n10838), .C(n9213), .D(n10839), .Y(n8994) );
  OAI22X1 U5645 ( .A(n9211), .B(n10836), .C(n9212), .D(n10838), .Y(n8995) );
  OAI21X1 U5647 ( .A(n9380), .B(n10850), .C(n4553), .Y(n8996) );
  NAND2X1 U5648 ( .A(\U_0/U_2/RX_CRC [11]), .B(n9381), .Y(n4553) );
  OAI22X1 U5649 ( .A(n9379), .B(n10835), .C(n9213), .D(n10850), .Y(n8997) );
  OAI22X1 U5651 ( .A(n9211), .B(n10833), .C(n9212), .D(n10835), .Y(n8998) );
  OAI21X1 U5653 ( .A(n9380), .B(n10855), .C(n4557), .Y(n8999) );
  NAND2X1 U5654 ( .A(\U_0/U_2/RX_CRC [10]), .B(n9381), .Y(n4557) );
  OAI22X1 U5655 ( .A(n9379), .B(n10832), .C(n9213), .D(n10855), .Y(n9000) );
  OAI22X1 U5657 ( .A(n9211), .B(n10830), .C(n9212), .D(n10832), .Y(n9001) );
  OAI21X1 U5659 ( .A(n9380), .B(n10854), .C(n4561), .Y(n9002) );
  NAND2X1 U5660 ( .A(\U_0/U_2/RX_CRC [9]), .B(n9381), .Y(n4561) );
  OAI22X1 U5661 ( .A(n9380), .B(n10853), .C(n9213), .D(n10854), .Y(n9003) );
  OAI22X1 U5663 ( .A(n9212), .B(n10853), .C(n4563), .D(n9211), .Y(n9004) );
  XNOR2X1 U5664 ( .A(\U_0/U_2/U_2/current_crc[1] ), .B(n4564), .Y(n4563) );
  OAI21X1 U5666 ( .A(n9380), .B(n10856), .C(n4566), .Y(n9005) );
  NAND2X1 U5667 ( .A(\U_0/U_2/RX_CRC [8]), .B(n9381), .Y(n4566) );
  OAI22X1 U5668 ( .A(n9380), .B(n10829), .C(n9213), .D(n10856), .Y(n9006) );
  OAI22X1 U5670 ( .A(n9212), .B(n10829), .C(n4568), .D(n9211), .Y(n9007) );
  XOR2X1 U5671 ( .A(n4569), .B(n4570), .Y(n4568) );
  XNOR2X1 U5672 ( .A(\U_0/U_2/U_2/current_crc[0] ), .B(n4564), .Y(n4569) );
  OAI21X1 U5674 ( .A(n9380), .B(n10848), .C(n4572), .Y(n9008) );
  NAND2X1 U5675 ( .A(\U_0/U_2/RX_CRC [7]), .B(n9381), .Y(n4572) );
  OAI22X1 U5676 ( .A(n9379), .B(n10847), .C(n9213), .D(n10848), .Y(n9009) );
  OAI22X1 U5678 ( .A(n9212), .B(n10847), .C(n4574), .D(n9211), .Y(n9010) );
  OAI21X1 U5679 ( .A(n9380), .B(n10844), .C(n4576), .Y(n9011) );
  NAND2X1 U5680 ( .A(\U_0/U_2/RX_CRC [6]), .B(n9381), .Y(n4576) );
  OAI22X1 U5681 ( .A(n9380), .B(n10843), .C(n9213), .D(n10844), .Y(n9012) );
  OAI22X1 U5683 ( .A(n9212), .B(n10843), .C(n4577), .D(n9211), .Y(n9013) );
  XNOR2X1 U5684 ( .A(n4578), .B(n4579), .Y(n4577) );
  OAI21X1 U5686 ( .A(n9381), .B(n10841), .C(n4581), .Y(n9014) );
  NAND2X1 U5687 ( .A(\U_0/U_2/RX_CRC [5]), .B(n9381), .Y(n4581) );
  OAI22X1 U5688 ( .A(n9379), .B(n10840), .C(n9213), .D(n10841), .Y(n9015) );
  OAI22X1 U5690 ( .A(n9212), .B(n10840), .C(n4582), .D(n9211), .Y(n9016) );
  OAI21X1 U5692 ( .A(n9381), .B(n10837), .C(n4584), .Y(n9017) );
  NAND2X1 U5693 ( .A(\U_0/U_2/RX_CRC [4]), .B(n9381), .Y(n4584) );
  OAI22X1 U5694 ( .A(n9380), .B(n10836), .C(n9213), .D(n10837), .Y(n9018) );
  OAI22X1 U5696 ( .A(n9212), .B(n10836), .C(n4585), .D(n9211), .Y(n9019) );
  XNOR2X1 U5697 ( .A(n4586), .B(n4587), .Y(n4585) );
  OAI21X1 U5699 ( .A(n9381), .B(n10834), .C(n4589), .Y(n9020) );
  NAND2X1 U5700 ( .A(\U_0/U_2/RX_CRC [3]), .B(n9382), .Y(n4589) );
  OAI22X1 U5701 ( .A(n9379), .B(n10833), .C(n9213), .D(n10834), .Y(n9021) );
  OAI22X1 U5703 ( .A(n9212), .B(n10833), .C(n4590), .D(n9211), .Y(n9022) );
  OAI21X1 U5705 ( .A(n9381), .B(n10831), .C(n4592), .Y(n9023) );
  NAND2X1 U5706 ( .A(\U_0/U_2/RX_CRC [2]), .B(n9382), .Y(n4592) );
  OAI22X1 U5707 ( .A(n9379), .B(n10830), .C(n9213), .D(n10831), .Y(n9024) );
  OAI22X1 U5709 ( .A(n9212), .B(n10830), .C(n4593), .D(n9211), .Y(n9025) );
  XNOR2X1 U5710 ( .A(n4594), .B(n4595), .Y(n4593) );
  OAI21X1 U5712 ( .A(n9381), .B(n10852), .C(n4597), .Y(n9026) );
  NAND2X1 U5713 ( .A(\U_0/U_2/RX_CRC [1]), .B(n9382), .Y(n4597) );
  OAI22X1 U5714 ( .A(n9379), .B(n10851), .C(n9213), .D(n10852), .Y(n9027) );
  OAI22X1 U5716 ( .A(n9212), .B(n10851), .C(n4599), .D(n9211), .Y(n9028) );
  XOR2X1 U5717 ( .A(n4600), .B(n4601), .Y(n4599) );
  OAI21X1 U5719 ( .A(n9381), .B(n10828), .C(n4603), .Y(n9029) );
  NAND2X1 U5720 ( .A(\U_0/U_2/RX_CRC [0]), .B(n9382), .Y(n4603) );
  OAI22X1 U5721 ( .A(n9379), .B(n10827), .C(n9213), .D(n10828), .Y(n9030) );
  OAI22X1 U5723 ( .A(n9212), .B(n10827), .C(n4605), .D(n9211), .Y(n9031) );
  OAI22X1 U5725 ( .A(n9531), .B(n10866), .C(RST), .D(n747), .Y(n9032) );
  NOR2X1 U5726 ( .A(n4607), .B(n4608), .Y(n747) );
  OAI21X1 U5727 ( .A(n4609), .B(n9690), .C(n4610), .Y(n4608) );
  OAI21X1 U5728 ( .A(n9714), .B(n10866), .C(n4611), .Y(n4607) );
  OAI21X1 U5730 ( .A(n4613), .B(n4614), .C(n4615), .Y(n4612) );
  NAND2X1 U5731 ( .A(n4616), .B(n10825), .Y(n4614) );
  OAI21X1 U5733 ( .A(n9693), .B(n10821), .C(n4620), .Y(n9033) );
  NAND3X1 U5734 ( .A(n9209), .B(n10821), .C(n9692), .Y(n4620) );
  OAI21X1 U5736 ( .A(n4624), .B(n10822), .C(n4626), .Y(n9034) );
  NAND3X1 U5737 ( .A(n9209), .B(n10822), .C(n4627), .Y(n4626) );
  NOR2X1 U5738 ( .A(n4628), .B(n10821), .Y(n4627) );
  AOI21X1 U5739 ( .A(n4629), .B(n10821), .C(n4623), .Y(n4624) );
  OAI21X1 U5740 ( .A(n9209), .B(n10796), .C(n4631), .Y(n4623) );
  OAI21X1 U5741 ( .A(n9691), .B(n10823), .C(n4634), .Y(n9035) );
  NAND3X1 U5742 ( .A(n9692), .B(n10823), .C(n9711), .Y(n4634) );
  OAI21X1 U5744 ( .A(n4637), .B(n10824), .C(n4639), .Y(n9036) );
  NAND3X1 U5745 ( .A(n9692), .B(n10824), .C(n4640), .Y(n4639) );
  NOR2X1 U5746 ( .A(n4641), .B(n10823), .Y(n4640) );
  NAND2X1 U5748 ( .A(n4629), .B(n4631), .Y(n4628) );
  AOI21X1 U5749 ( .A(n4629), .B(n10823), .C(n4636), .Y(n4637) );
  OAI21X1 U5750 ( .A(n9711), .B(n10796), .C(n4631), .Y(n4636) );
  NAND3X1 U5753 ( .A(\U_0/U_2/U_5/count[0] ), .B(n9209), .C(
        \U_0/U_2/U_5/count[1] ), .Y(n4641) );
  NOR2X1 U5754 ( .A(n10797), .B(n4643), .Y(n4629) );
  OAI21X1 U5755 ( .A(n9381), .B(n10857), .C(n4645), .Y(n9037) );
  NAND2X1 U5756 ( .A(\U_0/U_2/RX_CRC [15]), .B(n9382), .Y(n4645) );
  OAI22X1 U5757 ( .A(n9379), .B(n10826), .C(n9213), .D(n10857), .Y(n9038) );
  OAI22X1 U5761 ( .A(n9212), .B(n10826), .C(n4647), .D(n9211), .Y(n9039) );
  XNOR2X1 U5762 ( .A(n4605), .B(n10847), .Y(n4647) );
  XOR2X1 U5764 ( .A(n4648), .B(n4601), .Y(n4605) );
  XOR2X1 U5765 ( .A(n4590), .B(n4582), .Y(n4601) );
  XNOR2X1 U5766 ( .A(n4587), .B(n4578), .Y(n4582) );
  XNOR2X1 U5767 ( .A(\U_0/U_2/U_2/current_crc[12] ), .B(n9345), .Y(n4578) );
  XNOR2X1 U5768 ( .A(\U_0/U_2/U_2/current_crc[11] ), .B(n9343), .Y(n4587) );
  XNOR2X1 U5769 ( .A(n4595), .B(n4586), .Y(n4590) );
  XNOR2X1 U5770 ( .A(\U_0/U_2/U_2/current_crc[10] ), .B(n9341), .Y(n4586) );
  XNOR2X1 U5771 ( .A(\U_0/U_2/U_2/current_crc[9] ), .B(n9339), .Y(n4595) );
  XOR2X1 U5772 ( .A(n4600), .B(n4594), .Y(n4648) );
  XNOR2X1 U5773 ( .A(\U_0/U_2/U_2/current_crc[8] ), .B(n9337), .Y(n4594) );
  XOR2X1 U5774 ( .A(n4564), .B(n4574), .Y(n4600) );
  XNOR2X1 U5775 ( .A(n4579), .B(n4570), .Y(n4574) );
  XNOR2X1 U5776 ( .A(n10845), .B(n9350), .Y(n4570) );
  XNOR2X1 U5778 ( .A(\U_0/U_2/U_2/current_crc[13] ), .B(n9347), .Y(n4579) );
  XNOR2X1 U5779 ( .A(\U_0/U_2/U_2/current_crc[15] ), .B(n9351), .Y(n4564) );
  OAI22X1 U5785 ( .A(n9209), .B(n9337), .C(n9339), .D(n9183), .Y(n9040) );
  OAI22X1 U5786 ( .A(n9209), .B(n9339), .C(n9341), .D(n9183), .Y(n9041) );
  OAI22X1 U5788 ( .A(n9209), .B(n9341), .C(n9343), .D(n9183), .Y(n9042) );
  OAI22X1 U5790 ( .A(n9209), .B(n9343), .C(n9345), .D(n9183), .Y(n9043) );
  OAI22X1 U5791 ( .A(n9209), .B(n9345), .C(n9347), .D(n9183), .Y(n9044) );
  OAI22X1 U5792 ( .A(n9209), .B(n9347), .C(n9349), .D(n9183), .Y(n9045) );
  OAI22X1 U5794 ( .A(n9209), .B(n9349), .C(n9351), .D(n9183), .Y(n9046) );
  OAI22X1 U5796 ( .A(n9209), .B(n9351), .C(n9183), .D(n4651), .Y(n9047) );
  XNOR2X1 U5797 ( .A(n10814), .B(\U_0/U_2/U_1/DP_hold1 ), .Y(n4651) );
  NAND2X1 U5800 ( .A(n4653), .B(n4654), .Y(n9048) );
  AOI22X1 U5801 ( .A(DPRH), .B(n10811), .C(\U_0/U_2/U_1/DP_hold1 ), .D(n4656), 
        .Y(n4653) );
  OAI21X1 U5802 ( .A(n10814), .B(n4657), .C(n4658), .Y(n9049) );
  OAI21X1 U5803 ( .A(\U_0/U_2/U_1/DP_hold1 ), .B(n9694), .C(n4657), .Y(n4658)
         );
  NOR2X1 U5805 ( .A(\U_0/U_2/U_1/state[3] ), .B(n9192), .Y(n4654) );
  OAI21X1 U5806 ( .A(n4656), .B(n10811), .C(n4661), .Y(n4657) );
  NOR2X1 U5807 ( .A(n9192), .B(n9209), .Y(n4661) );
  NOR3X1 U5810 ( .A(n4664), .B(n4665), .C(n4666), .Y(n4663) );
  OAI21X1 U5811 ( .A(n9407), .B(n10790), .C(n4668), .Y(n9050) );
  AOI22X1 U5812 ( .A(n4669), .B(n4670), .C(n9412), .D(n10645), .Y(n4668) );
  OAI22X1 U5813 ( .A(n4673), .B(n4674), .C(n9208), .D(n4676), .Y(n4669) );
  OAI21X1 U5814 ( .A(\U_0/U_0/U_1/RCV_DATA [5]), .B(n4677), .C(n9411), .Y(
        n4674) );
  OAI21X1 U5815 ( .A(n10627), .B(n4680), .C(n9208), .Y(n4673) );
  AOI22X1 U5816 ( .A(n4681), .B(n4682), .C(n10749), .D(n10766), .Y(n4680) );
  OAI22X1 U5817 ( .A(\U_0/U_0/U_1/RCV_DATA [3]), .B(n4684), .C(n10680), .D(
        n4686), .Y(n4681) );
  AOI22X1 U5818 ( .A(n4687), .B(n4688), .C(n10731), .D(n9482), .Y(n4686) );
  OAI22X1 U5820 ( .A(n4690), .B(n10663), .C(\U_0/U_0/U_1/RCV_DATA [1]), .D(
        n4692), .Y(n4687) );
  NAND2X1 U5822 ( .A(n4693), .B(n4694), .Y(n4692) );
  AOI22X1 U5823 ( .A(n4695), .B(n9487), .C(n10714), .D(n10790), .Y(n4690) );
  NOR2X1 U5826 ( .A(n4697), .B(n4698), .Y(n4695) );
  NAND2X1 U5828 ( .A(n9726), .B(n4700), .Y(n9051) );
  AOI22X1 U5829 ( .A(n9408), .B(\U_0/U_0/U_1/U_8/currentPlainKey[62] ), .C(
        n9412), .D(n10698), .Y(n4700) );
  OAI22X1 U5831 ( .A(n4676), .B(n4670), .C(n4704), .D(n4705), .Y(n4703) );
  OAI21X1 U5832 ( .A(n4706), .B(n4707), .C(n9411), .Y(n4705) );
  OAI22X1 U5833 ( .A(n10764), .B(n9208), .C(n10766), .D(n4677), .Y(n4707) );
  OAI21X1 U5834 ( .A(n9383), .B(n4682), .C(n4708), .Y(n4706) );
  AOI22X1 U5835 ( .A(n10680), .B(n9481), .C(n10628), .D(n4710), .Y(n4708) );
  OAI21X1 U5836 ( .A(n9392), .B(n4688), .C(n4711), .Y(n4710) );
  NAND2X1 U5837 ( .A(n4712), .B(n4688), .Y(n4711) );
  OAI21X1 U5838 ( .A(n4713), .B(n4714), .C(n4715), .Y(n4712) );
  OAI21X1 U5839 ( .A(n4713), .B(n4697), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[62] ), .Y(n4715) );
  NAND2X1 U5840 ( .A(n4716), .B(n4694), .Y(n4688) );
  NAND2X1 U5842 ( .A(n4718), .B(n4670), .Y(n4704) );
  NAND2X1 U5843 ( .A(n4719), .B(n4720), .Y(n9052) );
  AOI22X1 U5844 ( .A(n4721), .B(n4722), .C(n10698), .D(n9360), .Y(n4720) );
  OAI21X1 U5845 ( .A(n10764), .B(n4670), .C(n4724), .Y(n4722) );
  OAI21X1 U5846 ( .A(n4725), .B(n4726), .C(n4670), .Y(n4724) );
  OAI22X1 U5847 ( .A(n10766), .B(n9208), .C(n9482), .D(n4682), .Y(n4726) );
  OAI21X1 U5848 ( .A(n4727), .B(n4717), .C(n4728), .Y(n4725) );
  AOI22X1 U5849 ( .A(n10680), .B(\U_0/U_0/U_1/RCV_DATA [1]), .C(n10627), .D(
        \U_0/U_0/U_1/RCV_DATA [3]), .Y(n4728) );
  NAND2X1 U5852 ( .A(n4729), .B(n4684), .Y(n4717) );
  NAND2X1 U5853 ( .A(n4730), .B(n4694), .Y(n4684) );
  AOI22X1 U5854 ( .A(n4731), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[61] ), .D(n10732), .Y(n4727) );
  NOR2X1 U5856 ( .A(n4697), .B(n4733), .Y(n4731) );
  AOI22X1 U5857 ( .A(n10647), .B(n9412), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[61] ), .D(n9406), .Y(n4719) );
  NAND2X1 U5858 ( .A(n4735), .B(n4736), .Y(n9053) );
  AOI22X1 U5859 ( .A(n4737), .B(n4738), .C(n10647), .D(n9360), .Y(n4736) );
  OAI21X1 U5860 ( .A(n9723), .B(n4740), .C(n4741), .Y(n4737) );
  AOI22X1 U5861 ( .A(n9405), .B(n10645), .C(n4743), .D(n10698), .Y(n4741) );
  OAI21X1 U5862 ( .A(n4744), .B(n4745), .C(n4670), .Y(n4740) );
  OAI22X1 U5863 ( .A(n9383), .B(n9208), .C(n9483), .D(n4677), .Y(n4745) );
  OAI21X1 U5864 ( .A(n9392), .B(n4682), .C(n4746), .Y(n4744) );
  NAND2X1 U5865 ( .A(n4729), .B(n4747), .Y(n4746) );
  OAI21X1 U5866 ( .A(n4748), .B(n4714), .C(n4749), .Y(n4747) );
  OAI21X1 U5867 ( .A(n4748), .B(n4697), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[60] ), .Y(n4749) );
  NOR2X1 U5868 ( .A(n4750), .B(n10749), .Y(n4729) );
  NAND2X1 U5870 ( .A(n4751), .B(n4694), .Y(n4682) );
  AOI22X1 U5872 ( .A(n10715), .B(n9412), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[60] ), .D(n9406), .Y(n4735) );
  NAND2X1 U5873 ( .A(n4753), .B(n4754), .Y(n9054) );
  AOI22X1 U5874 ( .A(n4755), .B(n4756), .C(n10715), .D(n9360), .Y(n4754) );
  OAI21X1 U5875 ( .A(n4757), .B(n9355), .C(n4759), .Y(n4756) );
  AOI22X1 U5876 ( .A(n4721), .B(n4760), .C(n9404), .D(n10698), .Y(n4759) );
  OAI21X1 U5877 ( .A(n9383), .B(n4670), .C(n4761), .Y(n4760) );
  OAI21X1 U5878 ( .A(n4762), .B(n4763), .C(n4670), .Y(n4761) );
  OAI22X1 U5879 ( .A(n9388), .B(n4677), .C(n4764), .D(n4750), .Y(n4763) );
  NAND2X1 U5880 ( .A(n4677), .B(n9208), .Y(n4750) );
  AOI22X1 U5881 ( .A(n4765), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[59] ), .D(n10750), .Y(n4764) );
  NOR2X1 U5883 ( .A(n4697), .B(n4767), .Y(n4765) );
  NAND2X1 U5884 ( .A(n4768), .B(n4694), .Y(n4677) );
  NOR2X1 U5885 ( .A(n9484), .B(n9208), .Y(n4762) );
  NOR2X1 U5886 ( .A(n10646), .B(n9409), .Y(n4721) );
  AOI22X1 U5887 ( .A(n10664), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[59] ), .D(n9406), .Y(n4753) );
  NAND2X1 U5888 ( .A(n4772), .B(n4773), .Y(n9055) );
  AOI22X1 U5889 ( .A(n4774), .B(n4775), .C(n10664), .D(n9360), .Y(n4773) );
  OAI21X1 U5890 ( .A(n9355), .B(n4738), .C(n4776), .Y(n4775) );
  AOI22X1 U5891 ( .A(n4777), .B(n4778), .C(n9403), .D(n10647), .Y(n4776) );
  NOR2X1 U5892 ( .A(n10647), .B(n10715), .Y(n4778) );
  NOR2X1 U5893 ( .A(n4779), .B(n9409), .Y(n4777) );
  AOI21X1 U5894 ( .A(n10698), .B(\U_0/U_0/U_1/RCV_DATA [3]), .C(n4780), .Y(
        n4779) );
  OAI21X1 U5895 ( .A(n9484), .B(n4670), .C(n4781), .Y(n4780) );
  NAND3X1 U5896 ( .A(n4718), .B(n4670), .C(n4782), .Y(n4781) );
  OAI22X1 U5897 ( .A(n9388), .B(n9208), .C(n9169), .D(n4784), .Y(n4782) );
  AOI22X1 U5898 ( .A(n4785), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[58] ), .D(n10629), .Y(n4784) );
  NOR2X1 U5900 ( .A(n4697), .B(n4787), .Y(n4785) );
  AOI22X1 U5903 ( .A(n10733), .B(n9412), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[58] ), .D(n9406), .Y(n4772) );
  NAND2X1 U5904 ( .A(n4790), .B(n4791), .Y(n9056) );
  AOI22X1 U5905 ( .A(n4792), .B(n4793), .C(n10733), .D(n9360), .Y(n4791) );
  OAI21X1 U5906 ( .A(n9355), .B(n4794), .C(n4795), .Y(n4793) );
  AOI22X1 U5907 ( .A(n4796), .B(n4755), .C(n10715), .D(n9405), .Y(n4795) );
  NOR2X1 U5908 ( .A(n4797), .B(n9409), .Y(n4796) );
  AOI21X1 U5909 ( .A(n10647), .B(\U_0/U_0/U_1/RCV_DATA [3]), .C(n4798), .Y(
        n4797) );
  OAI22X1 U5910 ( .A(n9483), .B(n4718), .C(n4799), .D(n10646), .Y(n4798) );
  AOI22X1 U5912 ( .A(n4801), .B(n4670), .C(n10645), .D(
        \U_0/U_0/U_1/RCV_DATA [1]), .Y(n4799) );
  NAND2X1 U5914 ( .A(n4694), .B(n4802), .Y(n4670) );
  OAI21X1 U5915 ( .A(n4803), .B(n4714), .C(n4804), .Y(n4801) );
  OAI21X1 U5916 ( .A(n4803), .B(n4697), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[57] ), .Y(n4804) );
  AOI22X1 U5917 ( .A(n10611), .B(n9412), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[57] ), .D(n9406), .Y(n4790) );
  NAND2X1 U5918 ( .A(n4806), .B(n4807), .Y(n9057) );
  AOI22X1 U5919 ( .A(n4808), .B(n4809), .C(n10611), .D(n9360), .Y(n4807) );
  OAI21X1 U5920 ( .A(n9355), .B(n4810), .C(n4811), .Y(n4809) );
  AOI22X1 U5921 ( .A(n4812), .B(n4774), .C(n10664), .D(n9404), .Y(n4811) );
  NOR2X1 U5922 ( .A(n4813), .B(n9409), .Y(n4812) );
  AOI21X1 U5923 ( .A(n10715), .B(\U_0/U_0/U_1/RCV_DATA [3]), .C(n4814), .Y(
        n4813) );
  OAI22X1 U5924 ( .A(n9483), .B(n4757), .C(n10715), .D(n4815), .Y(n4814) );
  AOI22X1 U5925 ( .A(n10698), .B(\U_0/U_0/U_1/RCV_DATA [1]), .C(n4800), .D(
        n4816), .Y(n4815) );
  OAI21X1 U5926 ( .A(n4817), .B(n4714), .C(n4818), .Y(n4816) );
  OAI21X1 U5927 ( .A(n4817), .B(n4697), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[56] ), .Y(n4818) );
  NAND2X1 U5928 ( .A(n10757), .B(n9486), .Y(n4714) );
  NAND2X1 U5930 ( .A(\U_0/U_0/U_1/U_8/address[3] ), .B(n4820), .Y(n4697) );
  NOR2X1 U5931 ( .A(n10647), .B(n10698), .Y(n4800) );
  NAND2X1 U5933 ( .A(n4821), .B(n10709), .Y(n4718) );
  AOI22X1 U5935 ( .A(n10682), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[56] ), .D(n4701), .Y(n4806) );
  NAND2X1 U5936 ( .A(n4824), .B(n4825), .Y(n9058) );
  AOI22X1 U5937 ( .A(n4826), .B(n4827), .C(n10682), .D(n9360), .Y(n4825) );
  OAI21X1 U5938 ( .A(n9355), .B(n4828), .C(n4829), .Y(n4827) );
  AOI22X1 U5939 ( .A(n4830), .B(n4792), .C(n10733), .D(n9405), .Y(n4829) );
  OAI21X1 U5941 ( .A(n9383), .B(n4794), .C(n4832), .Y(n4831) );
  AOI22X1 U5942 ( .A(n4755), .B(n4833), .C(n10715), .D(n9481), .Y(n4832) );
  OAI22X1 U5943 ( .A(n9388), .B(n4757), .C(n10647), .D(n4834), .Y(n4833) );
  AOI22X1 U5944 ( .A(n10699), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[55] ), .D(n4836), .Y(n4834) );
  NAND2X1 U5946 ( .A(n4837), .B(n10709), .Y(n4836) );
  NAND2X1 U5948 ( .A(n4821), .B(n10658), .Y(n4757) );
  NOR2X1 U5949 ( .A(n10664), .B(n10715), .Y(n4755) );
  AOI22X1 U5950 ( .A(n10630), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[55] ), .D(n9408), .Y(n4824) );
  NAND2X1 U5951 ( .A(n4840), .B(n4841), .Y(n9059) );
  AOI22X1 U5952 ( .A(n4842), .B(n4843), .C(n10630), .D(n9360), .Y(n4841) );
  OAI21X1 U5953 ( .A(n9355), .B(n4844), .C(n4845), .Y(n4843) );
  AOI22X1 U5954 ( .A(n4846), .B(n4808), .C(n10611), .D(n9405), .Y(n4845) );
  OAI21X1 U5956 ( .A(n9383), .B(n4810), .C(n4848), .Y(n4847) );
  AOI22X1 U5957 ( .A(n4774), .B(n4849), .C(n10664), .D(n9481), .Y(n4848) );
  OAI22X1 U5958 ( .A(n9388), .B(n4738), .C(n10715), .D(n4850), .Y(n4849) );
  AOI22X1 U5959 ( .A(n10648), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[54] ), .D(n4852), .Y(n4850) );
  NAND2X1 U5961 ( .A(n4837), .B(n10658), .Y(n4852) );
  NAND2X1 U5963 ( .A(n4821), .B(n10726), .Y(n4738) );
  NOR2X1 U5964 ( .A(n10733), .B(n10664), .Y(n4774) );
  AOI22X1 U5965 ( .A(n10713), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[54] ), .D(n9406), .Y(n4840) );
  NAND2X1 U5966 ( .A(n4855), .B(n4856), .Y(n9060) );
  AOI22X1 U5967 ( .A(n4857), .B(n4858), .C(n10713), .D(n9360), .Y(n4856) );
  OAI21X1 U5968 ( .A(n9355), .B(n4859), .C(n4860), .Y(n4858) );
  AOI22X1 U5969 ( .A(n4861), .B(n4826), .C(n10682), .D(n9405), .Y(n4860) );
  OAI21X1 U5971 ( .A(n9383), .B(n4828), .C(n4863), .Y(n4862) );
  AOI22X1 U5972 ( .A(n4792), .B(n4864), .C(n10733), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n4863) );
  OAI22X1 U5973 ( .A(n9388), .B(n4794), .C(n10664), .D(n4865), .Y(n4864) );
  AOI22X1 U5974 ( .A(n10716), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[53] ), .D(n4867), .Y(n4865) );
  NAND2X1 U5976 ( .A(n4837), .B(n10726), .Y(n4867) );
  NAND2X1 U5978 ( .A(n4821), .B(n10675), .Y(n4794) );
  NOR2X1 U5979 ( .A(n10611), .B(n10733), .Y(n4792) );
  AOI22X1 U5980 ( .A(n10662), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[53] ), .D(n9406), .Y(n4855) );
  NAND2X1 U5981 ( .A(n4870), .B(n4871), .Y(n9061) );
  AOI22X1 U5982 ( .A(n4872), .B(n4873), .C(n10662), .D(n9360), .Y(n4871) );
  OAI21X1 U5983 ( .A(n9355), .B(n4874), .C(n4875), .Y(n4873) );
  AOI22X1 U5984 ( .A(n4876), .B(n4842), .C(n10630), .D(n9405), .Y(n4875) );
  OAI21X1 U5986 ( .A(n9383), .B(n4844), .C(n4878), .Y(n4877) );
  AOI22X1 U5987 ( .A(n4808), .B(n4879), .C(n10611), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n4878) );
  OAI22X1 U5988 ( .A(n9388), .B(n4810), .C(n10733), .D(n4880), .Y(n4879) );
  AOI22X1 U5989 ( .A(n10665), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[52] ), .D(n4882), .Y(n4880) );
  NAND2X1 U5991 ( .A(n4837), .B(n10675), .Y(n4882) );
  NAND2X1 U5993 ( .A(n4821), .B(n10744), .Y(n4810) );
  NOR2X1 U5994 ( .A(n10682), .B(n10611), .Y(n4808) );
  AOI22X1 U5995 ( .A(n10730), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[52] ), .D(n9406), .Y(n4870) );
  NAND2X1 U5996 ( .A(n4885), .B(n4886), .Y(n9062) );
  AOI22X1 U5997 ( .A(n4887), .B(n4888), .C(n10730), .D(n9360), .Y(n4886) );
  OAI21X1 U5998 ( .A(n9355), .B(n4889), .C(n4890), .Y(n4888) );
  AOI22X1 U5999 ( .A(n4891), .B(n4857), .C(n10713), .D(n9405), .Y(n4890) );
  OAI21X1 U6001 ( .A(n9383), .B(n4859), .C(n4893), .Y(n4892) );
  AOI22X1 U6002 ( .A(n4826), .B(n4894), .C(n10682), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n4893) );
  OAI22X1 U6003 ( .A(n9388), .B(n4828), .C(n10611), .D(n4895), .Y(n4894) );
  AOI22X1 U6004 ( .A(n10734), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[51] ), .D(n4897), .Y(n4895) );
  NAND2X1 U6006 ( .A(n4837), .B(n10744), .Y(n4897) );
  NAND2X1 U6008 ( .A(n4821), .B(n10622), .Y(n4828) );
  NOR2X1 U6009 ( .A(n10630), .B(n10682), .Y(n4826) );
  AOI22X1 U6010 ( .A(n10679), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[51] ), .D(n9406), .Y(n4885) );
  NAND2X1 U6011 ( .A(n4900), .B(n4901), .Y(n9063) );
  AOI22X1 U6012 ( .A(n4902), .B(n4903), .C(n10679), .D(n9360), .Y(n4901) );
  OAI21X1 U6013 ( .A(n9355), .B(n4904), .C(n4905), .Y(n4903) );
  AOI22X1 U6014 ( .A(n4906), .B(n4872), .C(n10662), .D(n9405), .Y(n4905) );
  OAI21X1 U6016 ( .A(n9383), .B(n4874), .C(n4908), .Y(n4907) );
  AOI22X1 U6017 ( .A(n4842), .B(n4909), .C(n10630), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n4908) );
  OAI22X1 U6018 ( .A(n9388), .B(n4844), .C(n10682), .D(n4910), .Y(n4909) );
  AOI22X1 U6019 ( .A(n10612), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[50] ), .D(n4912), .Y(n4910) );
  NAND2X1 U6021 ( .A(n4837), .B(n10622), .Y(n4912) );
  NAND2X1 U6023 ( .A(n4821), .B(n10693), .Y(n4844) );
  NOR2X1 U6024 ( .A(n10713), .B(n10630), .Y(n4842) );
  AOI22X1 U6025 ( .A(n10748), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[50] ), .D(n9406), .Y(n4900) );
  NAND2X1 U6026 ( .A(n4915), .B(n4916), .Y(n9064) );
  AOI22X1 U6027 ( .A(n4917), .B(n4918), .C(n10748), .D(n9360), .Y(n4916) );
  OAI21X1 U6028 ( .A(n9355), .B(n4919), .C(n4920), .Y(n4918) );
  AOI22X1 U6029 ( .A(n4921), .B(n4887), .C(n10730), .D(n9405), .Y(n4920) );
  OAI21X1 U6031 ( .A(n9383), .B(n4889), .C(n4923), .Y(n4922) );
  AOI22X1 U6032 ( .A(n4857), .B(n4924), .C(n10713), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n4923) );
  OAI22X1 U6033 ( .A(n9388), .B(n4859), .C(n10630), .D(n4925), .Y(n4924) );
  AOI22X1 U6034 ( .A(n10683), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[49] ), .D(n4927), .Y(n4925) );
  NAND2X1 U6036 ( .A(n4837), .B(n10693), .Y(n4927) );
  NAND2X1 U6038 ( .A(n4821), .B(n10641), .Y(n4859) );
  NOR2X1 U6041 ( .A(n10662), .B(n10713), .Y(n4857) );
  AOI22X1 U6042 ( .A(n10626), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[49] ), .D(n9406), .Y(n4915) );
  NAND2X1 U6043 ( .A(n4932), .B(n4933), .Y(n9065) );
  AOI22X1 U6044 ( .A(n4934), .B(n4935), .C(n10626), .D(n9361), .Y(n4933) );
  OAI21X1 U6045 ( .A(n9355), .B(n4936), .C(n4937), .Y(n4935) );
  AOI22X1 U6046 ( .A(n4938), .B(n4902), .C(n10679), .D(n9405), .Y(n4937) );
  OAI21X1 U6048 ( .A(n9383), .B(n4904), .C(n4940), .Y(n4939) );
  AOI22X1 U6049 ( .A(n4872), .B(n4941), .C(n10662), .D(n9481), .Y(n4940) );
  OAI22X1 U6050 ( .A(n9388), .B(n4874), .C(n10713), .D(n4942), .Y(n4941) );
  AOI22X1 U6051 ( .A(n10631), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[48] ), .D(n4944), .Y(n4942) );
  NAND2X1 U6053 ( .A(n4837), .B(n10641), .Y(n4944) );
  NAND2X1 U6056 ( .A(n4945), .B(n4946), .Y(n4874) );
  NOR2X1 U6057 ( .A(n10730), .B(n10662), .Y(n4872) );
  AOI22X1 U6058 ( .A(n10697), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[48] ), .D(n4701), .Y(n4932) );
  NAND2X1 U6059 ( .A(n4948), .B(n4949), .Y(n9066) );
  AOI22X1 U6060 ( .A(n4950), .B(n4951), .C(n10697), .D(n9361), .Y(n4949) );
  OAI21X1 U6061 ( .A(n9355), .B(n4952), .C(n4953), .Y(n4951) );
  AOI22X1 U6062 ( .A(n4954), .B(n4917), .C(n10748), .D(n9405), .Y(n4953) );
  OAI21X1 U6064 ( .A(n9384), .B(n4919), .C(n4956), .Y(n4955) );
  AOI22X1 U6065 ( .A(n4887), .B(n4957), .C(n10730), .D(n9481), .Y(n4956) );
  OAI22X1 U6066 ( .A(n9388), .B(n4889), .C(n10662), .D(n4958), .Y(n4957) );
  AOI22X1 U6067 ( .A(n10700), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[47] ), .D(n4960), .Y(n4958) );
  NAND2X1 U6069 ( .A(n4961), .B(n10709), .Y(n4960) );
  NAND2X1 U6071 ( .A(n4945), .B(n4693), .Y(n4889) );
  NOR2X1 U6072 ( .A(n10679), .B(n10730), .Y(n4887) );
  AOI22X1 U6073 ( .A(n10644), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[47] ), .D(n9408), .Y(n4948) );
  NAND2X1 U6074 ( .A(n4963), .B(n4964), .Y(n9067) );
  AOI22X1 U6075 ( .A(n4965), .B(n4966), .C(n10644), .D(n9361), .Y(n4964) );
  OAI21X1 U6076 ( .A(n9356), .B(n4967), .C(n4968), .Y(n4966) );
  AOI22X1 U6077 ( .A(n4969), .B(n4934), .C(n10626), .D(n9405), .Y(n4968) );
  OAI21X1 U6079 ( .A(n9384), .B(n4936), .C(n4971), .Y(n4970) );
  AOI22X1 U6080 ( .A(n4902), .B(n4972), .C(n10679), .D(n9481), .Y(n4971) );
  OAI22X1 U6081 ( .A(n9390), .B(n4904), .C(n10730), .D(n4973), .Y(n4972) );
  AOI22X1 U6082 ( .A(n10649), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[46] ), .D(n4975), .Y(n4973) );
  NAND2X1 U6084 ( .A(n4961), .B(n10658), .Y(n4975) );
  NAND2X1 U6086 ( .A(n4945), .B(n4716), .Y(n4904) );
  NOR2X1 U6087 ( .A(n10748), .B(n10679), .Y(n4902) );
  AOI22X1 U6088 ( .A(n10701), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[46] ), .D(n9408), .Y(n4963) );
  NAND2X1 U6089 ( .A(n4977), .B(n4978), .Y(n9068) );
  AOI22X1 U6090 ( .A(n4979), .B(n4980), .C(n10701), .D(n9361), .Y(n4978) );
  OAI21X1 U6091 ( .A(n9356), .B(n4981), .C(n4982), .Y(n4980) );
  AOI22X1 U6092 ( .A(n4983), .B(n4950), .C(n10697), .D(n9405), .Y(n4982) );
  OAI21X1 U6094 ( .A(n9385), .B(n4952), .C(n4985), .Y(n4984) );
  AOI22X1 U6095 ( .A(n4917), .B(n4986), .C(n10748), .D(n9481), .Y(n4985) );
  OAI22X1 U6096 ( .A(n9389), .B(n4919), .C(n10679), .D(n4987), .Y(n4986) );
  AOI22X1 U6097 ( .A(n10717), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[45] ), .D(n4989), .Y(n4987) );
  NAND2X1 U6099 ( .A(n4961), .B(n10726), .Y(n4989) );
  NAND2X1 U6101 ( .A(n4945), .B(n4730), .Y(n4919) );
  NOR2X1 U6102 ( .A(n10626), .B(n10748), .Y(n4917) );
  AOI22X1 U6103 ( .A(n10650), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[45] ), .D(n9408), .Y(n4977) );
  NAND2X1 U6104 ( .A(n4991), .B(n4992), .Y(n9069) );
  AOI22X1 U6105 ( .A(n4993), .B(n4994), .C(n10650), .D(n9361), .Y(n4992) );
  OAI21X1 U6106 ( .A(n9356), .B(n4995), .C(n4996), .Y(n4994) );
  AOI22X1 U6107 ( .A(n4997), .B(n4965), .C(n10644), .D(n9405), .Y(n4996) );
  OAI21X1 U6109 ( .A(n9384), .B(n4967), .C(n4999), .Y(n4998) );
  AOI22X1 U6110 ( .A(n4934), .B(n5000), .C(n10626), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n4999) );
  OAI22X1 U6111 ( .A(n9389), .B(n4936), .C(n10748), .D(n5001), .Y(n5000) );
  AOI22X1 U6112 ( .A(n10666), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[44] ), .D(n5003), .Y(n5001) );
  NAND2X1 U6114 ( .A(n4961), .B(n10675), .Y(n5003) );
  NAND2X1 U6116 ( .A(n4945), .B(n4751), .Y(n4936) );
  NOR2X1 U6117 ( .A(n10697), .B(n10626), .Y(n4934) );
  AOI22X1 U6118 ( .A(n10718), .B(n9413), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[44] ), .D(n9408), .Y(n4991) );
  NAND2X1 U6119 ( .A(n5005), .B(n5006), .Y(n9070) );
  AOI22X1 U6120 ( .A(n5007), .B(n5008), .C(n10718), .D(n9361), .Y(n5006) );
  OAI21X1 U6121 ( .A(n9356), .B(n5009), .C(n5010), .Y(n5008) );
  AOI22X1 U6122 ( .A(n5011), .B(n4979), .C(n10701), .D(n9405), .Y(n5010) );
  OAI21X1 U6124 ( .A(n9384), .B(n4981), .C(n5013), .Y(n5012) );
  AOI22X1 U6125 ( .A(n4950), .B(n5014), .C(n10697), .D(n9481), .Y(n5013) );
  OAI22X1 U6126 ( .A(n9389), .B(n4952), .C(n10626), .D(n5015), .Y(n5014) );
  AOI22X1 U6127 ( .A(n10735), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[43] ), .D(n5017), .Y(n5015) );
  NAND2X1 U6129 ( .A(n4961), .B(n10744), .Y(n5017) );
  NAND2X1 U6131 ( .A(n4945), .B(n4768), .Y(n4952) );
  NOR2X1 U6132 ( .A(n10644), .B(n10697), .Y(n4950) );
  AOI22X1 U6133 ( .A(n10667), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[43] ), .D(n9408), .Y(n5005) );
  NAND2X1 U6134 ( .A(n5019), .B(n5020), .Y(n9071) );
  AOI22X1 U6135 ( .A(n5021), .B(n5022), .C(n10667), .D(n9361), .Y(n5020) );
  OAI21X1 U6136 ( .A(n9356), .B(n5023), .C(n5024), .Y(n5022) );
  AOI22X1 U6137 ( .A(n5025), .B(n4993), .C(n10650), .D(n9404), .Y(n5024) );
  OAI21X1 U6139 ( .A(n9384), .B(n4995), .C(n5027), .Y(n5026) );
  AOI22X1 U6140 ( .A(n4965), .B(n5028), .C(n10644), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n5027) );
  OAI22X1 U6141 ( .A(n9389), .B(n4967), .C(n10697), .D(n5029), .Y(n5028) );
  AOI22X1 U6142 ( .A(n10613), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[42] ), .D(n5031), .Y(n5029) );
  NAND2X1 U6144 ( .A(n4961), .B(n10622), .Y(n5031) );
  NAND2X1 U6146 ( .A(n4945), .B(n4788), .Y(n4967) );
  NOR2X1 U6147 ( .A(n10701), .B(n10644), .Y(n4965) );
  AOI22X1 U6148 ( .A(n10736), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[42] ), .D(n9408), .Y(n5019) );
  NAND2X1 U6149 ( .A(n5033), .B(n5034), .Y(n9072) );
  AOI22X1 U6150 ( .A(n5035), .B(n5036), .C(n10736), .D(n9361), .Y(n5034) );
  OAI21X1 U6151 ( .A(n9356), .B(n5037), .C(n5038), .Y(n5036) );
  AOI22X1 U6152 ( .A(n5039), .B(n5007), .C(n10718), .D(n9404), .Y(n5038) );
  OAI21X1 U6154 ( .A(n9384), .B(n5009), .C(n5041), .Y(n5040) );
  AOI22X1 U6155 ( .A(n4979), .B(n5042), .C(n10701), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n5041) );
  OAI22X1 U6156 ( .A(n9389), .B(n4981), .C(n10644), .D(n5043), .Y(n5042) );
  AOI22X1 U6157 ( .A(n10684), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[41] ), .D(n5045), .Y(n5043) );
  NAND2X1 U6159 ( .A(n4961), .B(n10693), .Y(n5045) );
  NAND2X1 U6161 ( .A(n4945), .B(n4802), .Y(n4981) );
  NOR2X1 U6162 ( .A(n10650), .B(n10701), .Y(n4979) );
  AOI22X1 U6163 ( .A(n10614), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[41] ), .D(n9408), .Y(n5033) );
  NAND2X1 U6164 ( .A(n5047), .B(n5048), .Y(n9073) );
  AOI22X1 U6165 ( .A(n5049), .B(n5050), .C(n10614), .D(n9361), .Y(n5048) );
  OAI21X1 U6166 ( .A(n9356), .B(n5051), .C(n5052), .Y(n5050) );
  AOI22X1 U6167 ( .A(n5053), .B(n5021), .C(n10667), .D(n9404), .Y(n5052) );
  OAI21X1 U6169 ( .A(n9384), .B(n5023), .C(n5055), .Y(n5054) );
  AOI22X1 U6170 ( .A(n4993), .B(n5056), .C(n10650), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n5055) );
  OAI22X1 U6171 ( .A(n9389), .B(n4995), .C(n10701), .D(n5057), .Y(n5056) );
  AOI22X1 U6172 ( .A(n10632), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[40] ), .D(n5059), .Y(n5057) );
  NAND2X1 U6174 ( .A(n4961), .B(n10641), .Y(n5059) );
  NAND2X1 U6177 ( .A(n5061), .B(n10709), .Y(n4995) );
  NOR2X1 U6178 ( .A(n10718), .B(n10650), .Y(n4993) );
  AOI22X1 U6179 ( .A(n10685), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[40] ), .D(n9408), .Y(n5047) );
  NAND2X1 U6180 ( .A(n5063), .B(n5064), .Y(n9074) );
  AOI22X1 U6181 ( .A(n5065), .B(n5066), .C(n10685), .D(n9361), .Y(n5064) );
  OAI21X1 U6182 ( .A(n9356), .B(n5067), .C(n5068), .Y(n5066) );
  AOI22X1 U6183 ( .A(n5069), .B(n5035), .C(n10736), .D(n9404), .Y(n5068) );
  OAI21X1 U6185 ( .A(n9384), .B(n5037), .C(n5071), .Y(n5070) );
  AOI22X1 U6186 ( .A(n5007), .B(n5072), .C(n10718), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n5071) );
  OAI22X1 U6187 ( .A(n9389), .B(n5009), .C(n10650), .D(n5073), .Y(n5072) );
  AOI22X1 U6188 ( .A(n10702), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[39] ), .D(n5075), .Y(n5073) );
  NAND2X1 U6190 ( .A(n5076), .B(n10709), .Y(n5075) );
  NAND2X1 U6192 ( .A(n5061), .B(n10658), .Y(n5009) );
  NOR2X1 U6193 ( .A(n10667), .B(n10718), .Y(n5007) );
  AOI22X1 U6194 ( .A(n10633), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[39] ), .D(n9408), .Y(n5063) );
  NAND2X1 U6195 ( .A(n5078), .B(n5079), .Y(n9075) );
  AOI22X1 U6196 ( .A(n5080), .B(n5081), .C(n10633), .D(n9361), .Y(n5079) );
  OAI21X1 U6197 ( .A(n9356), .B(n5082), .C(n5083), .Y(n5081) );
  AOI22X1 U6198 ( .A(n5084), .B(n5049), .C(n10614), .D(n9404), .Y(n5083) );
  OAI21X1 U6200 ( .A(n9384), .B(n5051), .C(n5086), .Y(n5085) );
  AOI22X1 U6201 ( .A(n5021), .B(n5087), .C(n10667), .D(
        \U_0/U_0/U_1/RCV_DATA [2]), .Y(n5086) );
  OAI22X1 U6202 ( .A(n9389), .B(n5023), .C(n10718), .D(n5088), .Y(n5087) );
  AOI22X1 U6203 ( .A(n10651), .B(\U_0/U_0/U_1/RCV_DATA [0]), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[38] ), .D(n5090), .Y(n5088) );
  NAND2X1 U6205 ( .A(n5076), .B(n10658), .Y(n5090) );
  NAND2X1 U6207 ( .A(n5061), .B(n10726), .Y(n5023) );
  NOR2X1 U6208 ( .A(n10736), .B(n10667), .Y(n5021) );
  AOI22X1 U6209 ( .A(n10712), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[38] ), .D(n9408), .Y(n5078) );
  NAND2X1 U6210 ( .A(n5092), .B(n5093), .Y(n9076) );
  AOI22X1 U6211 ( .A(n5094), .B(n5095), .C(n10712), .D(n9361), .Y(n5093) );
  OAI21X1 U6212 ( .A(n9356), .B(n5096), .C(n5097), .Y(n5095) );
  AOI22X1 U6213 ( .A(n5098), .B(n5065), .C(n10685), .D(n9404), .Y(n5097) );
  OAI21X1 U6215 ( .A(n9384), .B(n5067), .C(n5100), .Y(n5099) );
  AOI22X1 U6216 ( .A(n5035), .B(n5101), .C(n10736), .D(n9481), .Y(n5100) );
  OAI22X1 U6217 ( .A(n9389), .B(n5037), .C(n10667), .D(n5102), .Y(n5101) );
  AOI22X1 U6218 ( .A(n10719), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[37] ), .D(n5104), .Y(n5102) );
  NAND2X1 U6220 ( .A(n5076), .B(n10726), .Y(n5104) );
  NAND2X1 U6222 ( .A(n5061), .B(n10675), .Y(n5037) );
  NOR2X1 U6223 ( .A(n10614), .B(n10736), .Y(n5035) );
  AOI22X1 U6224 ( .A(n10661), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[37] ), .D(n9408), .Y(n5092) );
  NAND2X1 U6225 ( .A(n5106), .B(n5107), .Y(n9077) );
  AOI22X1 U6226 ( .A(n5108), .B(n5109), .C(n10661), .D(n9361), .Y(n5107) );
  OAI21X1 U6227 ( .A(n9356), .B(n5110), .C(n5111), .Y(n5109) );
  AOI22X1 U6228 ( .A(n5112), .B(n5080), .C(n10633), .D(n9404), .Y(n5111) );
  OAI21X1 U6230 ( .A(n9384), .B(n5082), .C(n5114), .Y(n5113) );
  AOI22X1 U6231 ( .A(n5049), .B(n5115), .C(n10614), .D(n9481), .Y(n5114) );
  OAI22X1 U6232 ( .A(n9389), .B(n5051), .C(n10736), .D(n5116), .Y(n5115) );
  AOI22X1 U6233 ( .A(n10668), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[36] ), .D(n5118), .Y(n5116) );
  NAND2X1 U6235 ( .A(n5076), .B(n10675), .Y(n5118) );
  NAND2X1 U6237 ( .A(n5061), .B(n10744), .Y(n5051) );
  NOR2X1 U6238 ( .A(n10685), .B(n10614), .Y(n5049) );
  AOI22X1 U6239 ( .A(n10729), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[36] ), .D(n9408), .Y(n5106) );
  NAND2X1 U6240 ( .A(n5120), .B(n5121), .Y(n9078) );
  AOI22X1 U6241 ( .A(n5122), .B(n5123), .C(n10729), .D(n9362), .Y(n5121) );
  OAI21X1 U6242 ( .A(n9356), .B(n5124), .C(n5125), .Y(n5123) );
  AOI22X1 U6243 ( .A(n5126), .B(n5094), .C(n10712), .D(n9404), .Y(n5125) );
  OAI21X1 U6245 ( .A(n9384), .B(n5096), .C(n5128), .Y(n5127) );
  AOI22X1 U6246 ( .A(n5065), .B(n5129), .C(n10685), .D(n9481), .Y(n5128) );
  OAI22X1 U6247 ( .A(n9389), .B(n5067), .C(n10614), .D(n5130), .Y(n5129) );
  AOI22X1 U6248 ( .A(n10737), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[35] ), .D(n5132), .Y(n5130) );
  NAND2X1 U6250 ( .A(n5076), .B(n10744), .Y(n5132) );
  NAND2X1 U6252 ( .A(n5061), .B(n10622), .Y(n5067) );
  NOR2X1 U6253 ( .A(n10633), .B(n10685), .Y(n5065) );
  AOI22X1 U6254 ( .A(n10678), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[35] ), .D(n9408), .Y(n5120) );
  NAND2X1 U6255 ( .A(n5134), .B(n5135), .Y(n9079) );
  AOI22X1 U6256 ( .A(n5136), .B(n5137), .C(n10678), .D(n9362), .Y(n5135) );
  OAI21X1 U6257 ( .A(n9356), .B(n5138), .C(n5139), .Y(n5137) );
  AOI22X1 U6258 ( .A(n5140), .B(n5108), .C(n10661), .D(n9404), .Y(n5139) );
  OAI21X1 U6260 ( .A(n9384), .B(n5110), .C(n5142), .Y(n5141) );
  AOI22X1 U6261 ( .A(n5080), .B(n5143), .C(n10633), .D(n9481), .Y(n5142) );
  OAI22X1 U6262 ( .A(n9389), .B(n5082), .C(n10685), .D(n5144), .Y(n5143) );
  AOI22X1 U6263 ( .A(n10615), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[34] ), .D(n5146), .Y(n5144) );
  NAND2X1 U6265 ( .A(n5076), .B(n10622), .Y(n5146) );
  NAND2X1 U6267 ( .A(n5061), .B(n10693), .Y(n5082) );
  NOR2X1 U6268 ( .A(n10712), .B(n10633), .Y(n5080) );
  AOI22X1 U6269 ( .A(n10747), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[34] ), .D(n4701), .Y(n5134) );
  NAND2X1 U6270 ( .A(n5148), .B(n5149), .Y(n9080) );
  AOI22X1 U6271 ( .A(n5150), .B(n5151), .C(n10747), .D(n9362), .Y(n5149) );
  OAI21X1 U6272 ( .A(n9357), .B(n5152), .C(n5153), .Y(n5151) );
  AOI22X1 U6273 ( .A(n5154), .B(n5122), .C(n10729), .D(n9404), .Y(n5153) );
  OAI21X1 U6275 ( .A(n9385), .B(n5124), .C(n5156), .Y(n5155) );
  AOI22X1 U6276 ( .A(n5094), .B(n5157), .C(n10712), .D(n9481), .Y(n5156) );
  OAI22X1 U6277 ( .A(n9389), .B(n5096), .C(n10633), .D(n5158), .Y(n5157) );
  AOI22X1 U6278 ( .A(n10686), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[33] ), .D(n5160), .Y(n5158) );
  NAND2X1 U6280 ( .A(n5076), .B(n10693), .Y(n5160) );
  NAND2X1 U6282 ( .A(n5061), .B(n10641), .Y(n5096) );
  NOR2X1 U6285 ( .A(n10661), .B(n10712), .Y(n5094) );
  AOI22X1 U6286 ( .A(n10625), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[33] ), .D(n4701), .Y(n5148) );
  NAND2X1 U6287 ( .A(n5162), .B(n5163), .Y(n9081) );
  AOI22X1 U6288 ( .A(n5164), .B(n5165), .C(n10625), .D(n9362), .Y(n5163) );
  OAI21X1 U6289 ( .A(n9357), .B(n5166), .C(n5167), .Y(n5165) );
  AOI22X1 U6290 ( .A(n5168), .B(n5136), .C(n10678), .D(n9404), .Y(n5167) );
  OAI21X1 U6292 ( .A(n9385), .B(n5138), .C(n5170), .Y(n5169) );
  AOI22X1 U6293 ( .A(n5108), .B(n5171), .C(n10661), .D(n9481), .Y(n5170) );
  OAI22X1 U6294 ( .A(n9390), .B(n5110), .C(n10712), .D(n5172), .Y(n5171) );
  AOI22X1 U6295 ( .A(n10634), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[32] ), .D(n5174), .Y(n5172) );
  NAND2X1 U6297 ( .A(n5076), .B(n10641), .Y(n5174) );
  NOR2X1 U6299 ( .A(n10758), .B(\U_0/U_0/U_1/U_8/address[4] ), .Y(n5060) );
  NAND2X1 U6301 ( .A(n5176), .B(n4946), .Y(n5110) );
  NOR2X1 U6302 ( .A(n10729), .B(n10661), .Y(n5108) );
  AOI22X1 U6303 ( .A(n10696), .B(n9414), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[32] ), .D(n4701), .Y(n5162) );
  NAND2X1 U6304 ( .A(n5178), .B(n5179), .Y(n9082) );
  AOI22X1 U6305 ( .A(n5180), .B(n5181), .C(n10696), .D(n9362), .Y(n5179) );
  OAI21X1 U6306 ( .A(n9357), .B(n5182), .C(n5183), .Y(n5181) );
  AOI22X1 U6307 ( .A(n5184), .B(n5150), .C(n10747), .D(n9404), .Y(n5183) );
  OAI21X1 U6309 ( .A(n9385), .B(n5152), .C(n5186), .Y(n5185) );
  AOI22X1 U6310 ( .A(n5122), .B(n5187), .C(n10729), .D(n9481), .Y(n5186) );
  OAI22X1 U6311 ( .A(n9390), .B(n5124), .C(n10661), .D(n5188), .Y(n5187) );
  AOI22X1 U6312 ( .A(n10703), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[31] ), .D(n5190), .Y(n5188) );
  NAND2X1 U6314 ( .A(n5191), .B(n10709), .Y(n5190) );
  NAND2X1 U6316 ( .A(n5176), .B(n4693), .Y(n5124) );
  NOR2X1 U6317 ( .A(n10678), .B(n10729), .Y(n5122) );
  AOI22X1 U6318 ( .A(n10643), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[31] ), .D(n4701), .Y(n5178) );
  NAND2X1 U6319 ( .A(n5193), .B(n5194), .Y(n9083) );
  AOI22X1 U6320 ( .A(n5195), .B(n5196), .C(n10643), .D(n9362), .Y(n5194) );
  OAI21X1 U6321 ( .A(n9357), .B(n5197), .C(n5198), .Y(n5196) );
  AOI22X1 U6322 ( .A(n5199), .B(n5164), .C(n10625), .D(n9404), .Y(n5198) );
  OAI21X1 U6324 ( .A(n9385), .B(n5166), .C(n5201), .Y(n5200) );
  AOI22X1 U6325 ( .A(n5136), .B(n5202), .C(n10678), .D(n9481), .Y(n5201) );
  OAI22X1 U6326 ( .A(n9390), .B(n5138), .C(n10729), .D(n5203), .Y(n5202) );
  AOI22X1 U6327 ( .A(n10652), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[30] ), .D(n5205), .Y(n5203) );
  NAND2X1 U6329 ( .A(n5191), .B(n10658), .Y(n5205) );
  NAND2X1 U6331 ( .A(n5176), .B(n4716), .Y(n5138) );
  NOR2X1 U6332 ( .A(n10747), .B(n10678), .Y(n5136) );
  AOI22X1 U6333 ( .A(n10704), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[30] ), .D(n9406), .Y(n5193) );
  NAND2X1 U6334 ( .A(n5207), .B(n5208), .Y(n9084) );
  AOI22X1 U6335 ( .A(n5209), .B(n5210), .C(n10704), .D(n9362), .Y(n5208) );
  OAI21X1 U6336 ( .A(n9357), .B(n5211), .C(n5212), .Y(n5210) );
  AOI22X1 U6337 ( .A(n5213), .B(n5180), .C(n10696), .D(n9403), .Y(n5212) );
  OAI21X1 U6339 ( .A(n9385), .B(n5182), .C(n5215), .Y(n5214) );
  AOI22X1 U6340 ( .A(n5150), .B(n5216), .C(n10747), .D(n9481), .Y(n5215) );
  OAI22X1 U6341 ( .A(n9390), .B(n5152), .C(n10678), .D(n5217), .Y(n5216) );
  AOI22X1 U6342 ( .A(n10720), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[29] ), .D(n5219), .Y(n5217) );
  NAND2X1 U6344 ( .A(n5191), .B(n10726), .Y(n5219) );
  NAND2X1 U6346 ( .A(n5176), .B(n4730), .Y(n5152) );
  NOR2X1 U6347 ( .A(n10625), .B(n10747), .Y(n5150) );
  AOI22X1 U6348 ( .A(n10653), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[29] ), .D(n4701), .Y(n5207) );
  NAND2X1 U6349 ( .A(n5221), .B(n5222), .Y(n9085) );
  AOI22X1 U6350 ( .A(n5223), .B(n5224), .C(n10653), .D(n9362), .Y(n5222) );
  OAI21X1 U6351 ( .A(n9357), .B(n5225), .C(n5226), .Y(n5224) );
  AOI22X1 U6352 ( .A(n5227), .B(n5195), .C(n10643), .D(n9403), .Y(n5226) );
  OAI21X1 U6354 ( .A(n9385), .B(n5197), .C(n5229), .Y(n5228) );
  AOI22X1 U6355 ( .A(n5164), .B(n5230), .C(n10625), .D(n9481), .Y(n5229) );
  OAI22X1 U6356 ( .A(n9390), .B(n5166), .C(n10747), .D(n5231), .Y(n5230) );
  AOI22X1 U6357 ( .A(n10669), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[28] ), .D(n5233), .Y(n5231) );
  NAND2X1 U6359 ( .A(n5191), .B(n10675), .Y(n5233) );
  NAND2X1 U6361 ( .A(n5176), .B(n4751), .Y(n5166) );
  NOR2X1 U6362 ( .A(n10696), .B(n10625), .Y(n5164) );
  AOI22X1 U6363 ( .A(n10721), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[28] ), .D(n9406), .Y(n5221) );
  NAND2X1 U6364 ( .A(n5235), .B(n5236), .Y(n9086) );
  AOI22X1 U6365 ( .A(n5237), .B(n5238), .C(n10721), .D(n9362), .Y(n5236) );
  OAI21X1 U6366 ( .A(n9357), .B(n5239), .C(n5240), .Y(n5238) );
  AOI22X1 U6367 ( .A(n5241), .B(n5209), .C(n10704), .D(n9405), .Y(n5240) );
  OAI21X1 U6369 ( .A(n9385), .B(n5211), .C(n5243), .Y(n5242) );
  AOI22X1 U6370 ( .A(n5180), .B(n5244), .C(n10696), .D(n9481), .Y(n5243) );
  OAI22X1 U6371 ( .A(n9390), .B(n5182), .C(n10625), .D(n5245), .Y(n5244) );
  AOI22X1 U6372 ( .A(n10738), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[27] ), .D(n5247), .Y(n5245) );
  NAND2X1 U6374 ( .A(n5191), .B(n10744), .Y(n5247) );
  NAND2X1 U6376 ( .A(n5176), .B(n4768), .Y(n5182) );
  NOR2X1 U6377 ( .A(n10643), .B(n10696), .Y(n5180) );
  AOI22X1 U6378 ( .A(n10670), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[27] ), .D(n4701), .Y(n5235) );
  NAND2X1 U6379 ( .A(n5249), .B(n5250), .Y(n9087) );
  AOI22X1 U6380 ( .A(n5251), .B(n5252), .C(n10670), .D(n9362), .Y(n5250) );
  OAI21X1 U6381 ( .A(n9357), .B(n5253), .C(n5254), .Y(n5252) );
  AOI22X1 U6382 ( .A(n5255), .B(n5223), .C(n10653), .D(n9404), .Y(n5254) );
  OAI21X1 U6384 ( .A(n9385), .B(n5225), .C(n5257), .Y(n5256) );
  AOI22X1 U6385 ( .A(n5195), .B(n5258), .C(n10643), .D(n9481), .Y(n5257) );
  OAI22X1 U6386 ( .A(n9390), .B(n5197), .C(n10696), .D(n5259), .Y(n5258) );
  AOI22X1 U6387 ( .A(n10616), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[26] ), .D(n5261), .Y(n5259) );
  NAND2X1 U6389 ( .A(n5191), .B(n10622), .Y(n5261) );
  NAND2X1 U6391 ( .A(n5176), .B(n4788), .Y(n5197) );
  NOR2X1 U6392 ( .A(n10704), .B(n10643), .Y(n5195) );
  AOI22X1 U6393 ( .A(n10739), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[26] ), .D(n9406), .Y(n5249) );
  NAND2X1 U6394 ( .A(n5263), .B(n5264), .Y(n9088) );
  AOI22X1 U6395 ( .A(n5265), .B(n5266), .C(n10739), .D(n9362), .Y(n5264) );
  OAI21X1 U6396 ( .A(n9357), .B(n5267), .C(n5268), .Y(n5266) );
  AOI22X1 U6397 ( .A(n5269), .B(n5237), .C(n10721), .D(n9405), .Y(n5268) );
  OAI21X1 U6399 ( .A(n9385), .B(n5239), .C(n5271), .Y(n5270) );
  AOI22X1 U6400 ( .A(n5209), .B(n5272), .C(n10704), .D(n9481), .Y(n5271) );
  OAI22X1 U6401 ( .A(n9390), .B(n5211), .C(n10643), .D(n5273), .Y(n5272) );
  AOI22X1 U6402 ( .A(n10687), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[25] ), .D(n5275), .Y(n5273) );
  NAND2X1 U6404 ( .A(n5191), .B(n10693), .Y(n5275) );
  NAND2X1 U6406 ( .A(n5176), .B(n4802), .Y(n5211) );
  NOR2X1 U6407 ( .A(n10653), .B(n10704), .Y(n5209) );
  AOI22X1 U6408 ( .A(n10617), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[25] ), .D(n9406), .Y(n5263) );
  NAND2X1 U6409 ( .A(n5277), .B(n5278), .Y(n9089) );
  AOI22X1 U6410 ( .A(n5279), .B(n5280), .C(n10617), .D(n9362), .Y(n5278) );
  OAI21X1 U6411 ( .A(n9357), .B(n5281), .C(n5282), .Y(n5280) );
  AOI22X1 U6412 ( .A(n5283), .B(n5251), .C(n10670), .D(n9403), .Y(n5282) );
  OAI21X1 U6414 ( .A(n9385), .B(n5253), .C(n5285), .Y(n5284) );
  AOI22X1 U6415 ( .A(n5223), .B(n5286), .C(n10653), .D(n9481), .Y(n5285) );
  OAI22X1 U6416 ( .A(n9390), .B(n5225), .C(n10704), .D(n5287), .Y(n5286) );
  AOI22X1 U6417 ( .A(n10635), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[24] ), .D(n5289), .Y(n5287) );
  NAND2X1 U6419 ( .A(n5191), .B(n10641), .Y(n5289) );
  NAND2X1 U6422 ( .A(n5291), .B(n10709), .Y(n5225) );
  NOR2X1 U6423 ( .A(n10721), .B(n10653), .Y(n5223) );
  AOI22X1 U6424 ( .A(n10688), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[24] ), .D(n9406), .Y(n5277) );
  NAND2X1 U6425 ( .A(n5293), .B(n5294), .Y(n9090) );
  AOI22X1 U6426 ( .A(n5295), .B(n5296), .C(n10688), .D(n9362), .Y(n5294) );
  OAI21X1 U6427 ( .A(n9357), .B(n5297), .C(n5298), .Y(n5296) );
  AOI22X1 U6428 ( .A(n5299), .B(n5265), .C(n10739), .D(n9404), .Y(n5298) );
  OAI21X1 U6430 ( .A(n9385), .B(n5267), .C(n5301), .Y(n5300) );
  AOI22X1 U6431 ( .A(n5237), .B(n5302), .C(n10721), .D(n9481), .Y(n5301) );
  OAI22X1 U6432 ( .A(n9390), .B(n5239), .C(n10653), .D(n5303), .Y(n5302) );
  AOI22X1 U6433 ( .A(n10705), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[23] ), .D(n5305), .Y(n5303) );
  NAND2X1 U6435 ( .A(n5306), .B(n10709), .Y(n5305) );
  NAND2X1 U6437 ( .A(n5291), .B(n10658), .Y(n5239) );
  NOR2X1 U6438 ( .A(n10670), .B(n10721), .Y(n5237) );
  AOI22X1 U6439 ( .A(n10636), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[23] ), .D(n9406), .Y(n5293) );
  NAND2X1 U6440 ( .A(n5308), .B(n5309), .Y(n9091) );
  AOI22X1 U6441 ( .A(n5310), .B(n5311), .C(n10636), .D(n9363), .Y(n5309) );
  OAI21X1 U6442 ( .A(n9357), .B(n5312), .C(n5313), .Y(n5311) );
  AOI22X1 U6443 ( .A(n5314), .B(n5279), .C(n10617), .D(n9405), .Y(n5313) );
  OAI21X1 U6445 ( .A(n9385), .B(n5281), .C(n5316), .Y(n5315) );
  AOI22X1 U6446 ( .A(n5251), .B(n5317), .C(n10670), .D(n9481), .Y(n5316) );
  OAI22X1 U6447 ( .A(n9390), .B(n5253), .C(n10721), .D(n5318), .Y(n5317) );
  AOI22X1 U6448 ( .A(n10654), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[22] ), .D(n5320), .Y(n5318) );
  NAND2X1 U6450 ( .A(n5306), .B(n10658), .Y(n5320) );
  NAND2X1 U6452 ( .A(n5291), .B(n10726), .Y(n5253) );
  NOR2X1 U6453 ( .A(n10739), .B(n10670), .Y(n5251) );
  AOI22X1 U6454 ( .A(n10711), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[22] ), .D(n9406), .Y(n5308) );
  NAND2X1 U6455 ( .A(n5322), .B(n5323), .Y(n9092) );
  AOI22X1 U6456 ( .A(n5324), .B(n5325), .C(n10711), .D(n9363), .Y(n5323) );
  OAI21X1 U6457 ( .A(n9357), .B(n5326), .C(n5327), .Y(n5325) );
  AOI22X1 U6458 ( .A(n5328), .B(n5295), .C(n10688), .D(n9403), .Y(n5327) );
  OAI21X1 U6460 ( .A(n9386), .B(n5297), .C(n5330), .Y(n5329) );
  AOI22X1 U6461 ( .A(n5265), .B(n5331), .C(n10739), .D(n9481), .Y(n5330) );
  OAI22X1 U6462 ( .A(n9390), .B(n5267), .C(n10670), .D(n5332), .Y(n5331) );
  AOI22X1 U6463 ( .A(n10722), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[21] ), .D(n5334), .Y(n5332) );
  NAND2X1 U6465 ( .A(n5306), .B(n10726), .Y(n5334) );
  NAND2X1 U6467 ( .A(n5291), .B(n10675), .Y(n5267) );
  NOR2X1 U6468 ( .A(n10617), .B(n10739), .Y(n5265) );
  AOI22X1 U6469 ( .A(n10660), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[21] ), .D(n9406), .Y(n5322) );
  NAND2X1 U6470 ( .A(n5336), .B(n5337), .Y(n9093) );
  AOI22X1 U6471 ( .A(n5338), .B(n5339), .C(n10660), .D(n9363), .Y(n5337) );
  OAI21X1 U6472 ( .A(n9358), .B(n5340), .C(n5341), .Y(n5339) );
  AOI22X1 U6473 ( .A(n5342), .B(n5310), .C(n10636), .D(n9404), .Y(n5341) );
  OAI21X1 U6475 ( .A(n9386), .B(n5312), .C(n5344), .Y(n5343) );
  AOI22X1 U6476 ( .A(n5279), .B(n5345), .C(n10617), .D(n9481), .Y(n5344) );
  OAI22X1 U6477 ( .A(n9391), .B(n5281), .C(n10739), .D(n5346), .Y(n5345) );
  AOI22X1 U6478 ( .A(n10671), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[20] ), .D(n5348), .Y(n5346) );
  NAND2X1 U6480 ( .A(n5306), .B(n10675), .Y(n5348) );
  NAND2X1 U6482 ( .A(n5291), .B(n10744), .Y(n5281) );
  NOR2X1 U6483 ( .A(n10688), .B(n10617), .Y(n5279) );
  AOI22X1 U6484 ( .A(n10728), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[20] ), .D(n9406), .Y(n5336) );
  NAND2X1 U6485 ( .A(n5350), .B(n5351), .Y(n9094) );
  AOI22X1 U6486 ( .A(n5352), .B(n5353), .C(n10728), .D(n9363), .Y(n5351) );
  OAI21X1 U6487 ( .A(n9358), .B(n5354), .C(n5355), .Y(n5353) );
  AOI22X1 U6488 ( .A(n5356), .B(n5324), .C(n10711), .D(n9405), .Y(n5355) );
  OAI21X1 U6490 ( .A(n9386), .B(n5326), .C(n5358), .Y(n5357) );
  AOI22X1 U6491 ( .A(n5295), .B(n5359), .C(n10688), .D(n9481), .Y(n5358) );
  OAI22X1 U6492 ( .A(n9391), .B(n5297), .C(n10617), .D(n5360), .Y(n5359) );
  AOI22X1 U6493 ( .A(n10740), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[19] ), .D(n5362), .Y(n5360) );
  NAND2X1 U6495 ( .A(n5306), .B(n10744), .Y(n5362) );
  NAND2X1 U6497 ( .A(n5291), .B(n10622), .Y(n5297) );
  NOR2X1 U6498 ( .A(n10636), .B(n10688), .Y(n5295) );
  AOI22X1 U6499 ( .A(n10677), .B(n9415), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[19] ), .D(n9406), .Y(n5350) );
  NAND2X1 U6500 ( .A(n5364), .B(n5365), .Y(n9095) );
  AOI22X1 U6501 ( .A(n5366), .B(n5367), .C(n10677), .D(n9363), .Y(n5365) );
  OAI21X1 U6502 ( .A(n9358), .B(n5368), .C(n5369), .Y(n5367) );
  AOI22X1 U6503 ( .A(n5370), .B(n5338), .C(n10660), .D(n9403), .Y(n5369) );
  OAI21X1 U6505 ( .A(n9386), .B(n5340), .C(n5372), .Y(n5371) );
  AOI22X1 U6506 ( .A(n5310), .B(n5373), .C(n10636), .D(n9481), .Y(n5372) );
  OAI22X1 U6507 ( .A(n9391), .B(n5312), .C(n10688), .D(n5374), .Y(n5373) );
  AOI22X1 U6508 ( .A(n10618), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[18] ), .D(n5376), .Y(n5374) );
  NAND2X1 U6510 ( .A(n5306), .B(n10622), .Y(n5376) );
  NAND2X1 U6512 ( .A(n5291), .B(n10693), .Y(n5312) );
  NOR2X1 U6513 ( .A(n10711), .B(n10636), .Y(n5310) );
  AOI22X1 U6514 ( .A(n10746), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[18] ), .D(n9406), .Y(n5364) );
  NAND2X1 U6515 ( .A(n5378), .B(n5379), .Y(n9096) );
  AOI22X1 U6516 ( .A(n5380), .B(n5381), .C(n10746), .D(n9363), .Y(n5379) );
  OAI21X1 U6517 ( .A(n9358), .B(n5382), .C(n5383), .Y(n5381) );
  AOI22X1 U6518 ( .A(n5384), .B(n5352), .C(n10728), .D(n9404), .Y(n5383) );
  OAI21X1 U6520 ( .A(n9386), .B(n5354), .C(n5386), .Y(n5385) );
  AOI22X1 U6521 ( .A(n5324), .B(n5387), .C(n10711), .D(n9481), .Y(n5386) );
  OAI22X1 U6522 ( .A(n9391), .B(n5326), .C(n10636), .D(n5388), .Y(n5387) );
  AOI22X1 U6523 ( .A(n10689), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[17] ), .D(n5390), .Y(n5388) );
  NAND2X1 U6525 ( .A(n5306), .B(n10693), .Y(n5390) );
  NAND2X1 U6527 ( .A(n5291), .B(n10641), .Y(n5326) );
  NOR2X1 U6530 ( .A(n10660), .B(n10711), .Y(n5324) );
  AOI22X1 U6531 ( .A(n10624), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[17] ), .D(n9406), .Y(n5378) );
  NAND2X1 U6532 ( .A(n5392), .B(n5393), .Y(n9097) );
  AOI22X1 U6533 ( .A(n5394), .B(n5395), .C(n10624), .D(n9363), .Y(n5393) );
  OAI21X1 U6534 ( .A(n9358), .B(n5396), .C(n5397), .Y(n5395) );
  AOI22X1 U6535 ( .A(n5398), .B(n5366), .C(n10677), .D(n9403), .Y(n5397) );
  OAI21X1 U6537 ( .A(n9386), .B(n5368), .C(n5400), .Y(n5399) );
  AOI22X1 U6538 ( .A(n5338), .B(n5401), .C(n10660), .D(n9481), .Y(n5400) );
  OAI22X1 U6539 ( .A(n9391), .B(n5340), .C(n10711), .D(n5402), .Y(n5401) );
  AOI22X1 U6540 ( .A(n10637), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[16] ), .D(n5404), .Y(n5402) );
  NAND2X1 U6542 ( .A(n5306), .B(n10641), .Y(n5404) );
  NOR2X1 U6544 ( .A(n10759), .B(\U_0/U_0/U_1/U_8/address[5] ), .Y(n5290) );
  NAND2X1 U6546 ( .A(n5406), .B(n4946), .Y(n5340) );
  NOR2X1 U6547 ( .A(n10728), .B(n10660), .Y(n5338) );
  AOI22X1 U6548 ( .A(n10695), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[16] ), .D(n9406), .Y(n5392) );
  NAND2X1 U6549 ( .A(n5408), .B(n5409), .Y(n9098) );
  AOI22X1 U6550 ( .A(n5410), .B(n5411), .C(n10695), .D(n9363), .Y(n5409) );
  OAI21X1 U6551 ( .A(n9358), .B(n5412), .C(n5413), .Y(n5411) );
  AOI22X1 U6552 ( .A(n5414), .B(n5380), .C(n10746), .D(n9403), .Y(n5413) );
  OAI21X1 U6554 ( .A(n9386), .B(n5382), .C(n5416), .Y(n5415) );
  AOI22X1 U6555 ( .A(n5352), .B(n5417), .C(n10728), .D(n9481), .Y(n5416) );
  OAI22X1 U6556 ( .A(n9391), .B(n5354), .C(n10660), .D(n5418), .Y(n5417) );
  AOI22X1 U6557 ( .A(n10706), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[15] ), .D(n5420), .Y(n5418) );
  NAND2X1 U6559 ( .A(n5421), .B(n10709), .Y(n5420) );
  NAND2X1 U6561 ( .A(n5406), .B(n4693), .Y(n5354) );
  NOR2X1 U6562 ( .A(n10677), .B(n10728), .Y(n5352) );
  AOI22X1 U6563 ( .A(n10642), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[15] ), .D(n9406), .Y(n5408) );
  NAND2X1 U6564 ( .A(n5423), .B(n5424), .Y(n9099) );
  AOI22X1 U6565 ( .A(n5425), .B(n5426), .C(n10642), .D(n9363), .Y(n5424) );
  OAI21X1 U6566 ( .A(n9358), .B(n5427), .C(n5428), .Y(n5426) );
  AOI22X1 U6567 ( .A(n5429), .B(n5394), .C(n10624), .D(n9403), .Y(n5428) );
  OAI21X1 U6569 ( .A(n9386), .B(n5396), .C(n5431), .Y(n5430) );
  AOI22X1 U6570 ( .A(n5366), .B(n5432), .C(n10677), .D(n9481), .Y(n5431) );
  OAI22X1 U6571 ( .A(n9391), .B(n5368), .C(n10728), .D(n5433), .Y(n5432) );
  AOI22X1 U6572 ( .A(n10655), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[14] ), .D(n5435), .Y(n5433) );
  NAND2X1 U6574 ( .A(n5421), .B(n10658), .Y(n5435) );
  NAND2X1 U6576 ( .A(n5406), .B(n4716), .Y(n5368) );
  NOR2X1 U6577 ( .A(n10746), .B(n10677), .Y(n5366) );
  AOI22X1 U6578 ( .A(n10707), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[14] ), .D(n4701), .Y(n5423) );
  NAND2X1 U6579 ( .A(n5437), .B(n5438), .Y(n9100) );
  AOI22X1 U6580 ( .A(n5439), .B(n5440), .C(n10707), .D(n9363), .Y(n5438) );
  OAI21X1 U6581 ( .A(n9358), .B(n5441), .C(n5442), .Y(n5440) );
  AOI22X1 U6582 ( .A(n5443), .B(n5410), .C(n10695), .D(n9403), .Y(n5442) );
  OAI21X1 U6584 ( .A(n9386), .B(n5412), .C(n5445), .Y(n5444) );
  AOI22X1 U6585 ( .A(n5380), .B(n5446), .C(n10746), .D(n9481), .Y(n5445) );
  OAI22X1 U6586 ( .A(n9391), .B(n5382), .C(n10677), .D(n5447), .Y(n5446) );
  AOI22X1 U6587 ( .A(n10723), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[13] ), .D(n5449), .Y(n5447) );
  NAND2X1 U6589 ( .A(n5421), .B(n10726), .Y(n5449) );
  NAND2X1 U6591 ( .A(n5406), .B(n4730), .Y(n5382) );
  NOR2X1 U6592 ( .A(n10624), .B(n10746), .Y(n5380) );
  AOI22X1 U6593 ( .A(n10656), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[13] ), .D(n9406), .Y(n5437) );
  NAND2X1 U6594 ( .A(n5451), .B(n5452), .Y(n9101) );
  AOI22X1 U6595 ( .A(n5453), .B(n5454), .C(n10656), .D(n9363), .Y(n5452) );
  OAI21X1 U6596 ( .A(n9358), .B(n5455), .C(n5456), .Y(n5454) );
  AOI22X1 U6597 ( .A(n5457), .B(n5425), .C(n10642), .D(n9403), .Y(n5456) );
  OAI21X1 U6599 ( .A(n9386), .B(n5427), .C(n5459), .Y(n5458) );
  AOI22X1 U6600 ( .A(n5394), .B(n5460), .C(n10624), .D(n9481), .Y(n5459) );
  OAI22X1 U6601 ( .A(n9391), .B(n5396), .C(n10746), .D(n5461), .Y(n5460) );
  AOI22X1 U6602 ( .A(n10672), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[12] ), .D(n5463), .Y(n5461) );
  NAND2X1 U6604 ( .A(n5421), .B(n10675), .Y(n5463) );
  NAND2X1 U6606 ( .A(n5406), .B(n4751), .Y(n5396) );
  NOR2X1 U6607 ( .A(n10695), .B(n10624), .Y(n5394) );
  AOI22X1 U6608 ( .A(n10724), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[12] ), .D(n4701), .Y(n5451) );
  NAND2X1 U6609 ( .A(n5465), .B(n5466), .Y(n9102) );
  AOI22X1 U6610 ( .A(n5467), .B(n5468), .C(n10724), .D(n9363), .Y(n5466) );
  OAI21X1 U6611 ( .A(n9358), .B(n5469), .C(n5470), .Y(n5468) );
  AOI22X1 U6612 ( .A(n5471), .B(n5439), .C(n10707), .D(n9403), .Y(n5470) );
  OAI21X1 U6614 ( .A(n9386), .B(n5441), .C(n5473), .Y(n5472) );
  AOI22X1 U6615 ( .A(n5410), .B(n5474), .C(n10695), .D(n9481), .Y(n5473) );
  OAI22X1 U6616 ( .A(n9391), .B(n5412), .C(n10624), .D(n5475), .Y(n5474) );
  AOI22X1 U6617 ( .A(n10741), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[11] ), .D(n5477), .Y(n5475) );
  NAND2X1 U6619 ( .A(n5421), .B(n10744), .Y(n5477) );
  NAND2X1 U6621 ( .A(n5406), .B(n4768), .Y(n5412) );
  NOR2X1 U6622 ( .A(n10642), .B(n10695), .Y(n5410) );
  AOI22X1 U6623 ( .A(n10673), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[11] ), .D(n4701), .Y(n5465) );
  NAND2X1 U6624 ( .A(n5479), .B(n5480), .Y(n9103) );
  AOI22X1 U6625 ( .A(n5481), .B(n5482), .C(n10673), .D(n9363), .Y(n5480) );
  OAI21X1 U6626 ( .A(n9358), .B(n5483), .C(n5484), .Y(n5482) );
  AOI22X1 U6627 ( .A(n5485), .B(n5453), .C(n10656), .D(n9403), .Y(n5484) );
  OAI21X1 U6629 ( .A(n9386), .B(n5455), .C(n5487), .Y(n5486) );
  AOI22X1 U6630 ( .A(n5425), .B(n5488), .C(n10642), .D(n9481), .Y(n5487) );
  OAI22X1 U6631 ( .A(n9391), .B(n5427), .C(n10695), .D(n5489), .Y(n5488) );
  AOI22X1 U6632 ( .A(n10619), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[10] ), .D(n5491), .Y(n5489) );
  NAND2X1 U6634 ( .A(n5421), .B(n10622), .Y(n5491) );
  NAND2X1 U6636 ( .A(n5406), .B(n4788), .Y(n5427) );
  NOR2X1 U6637 ( .A(n10707), .B(n10642), .Y(n5425) );
  AOI22X1 U6638 ( .A(n10742), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[10] ), .D(n9408), .Y(n5479) );
  NAND2X1 U6639 ( .A(n5493), .B(n5494), .Y(n9104) );
  AOI22X1 U6640 ( .A(n5495), .B(n5496), .C(n10742), .D(n9364), .Y(n5494) );
  OAI21X1 U6641 ( .A(n9358), .B(n5497), .C(n5498), .Y(n5496) );
  AOI22X1 U6642 ( .A(n5499), .B(n5467), .C(n10724), .D(n9403), .Y(n5498) );
  OAI21X1 U6644 ( .A(n9386), .B(n5469), .C(n5501), .Y(n5500) );
  AOI22X1 U6645 ( .A(n5439), .B(n5502), .C(n10707), .D(n9481), .Y(n5501) );
  OAI22X1 U6646 ( .A(n9391), .B(n5441), .C(n10642), .D(n5503), .Y(n5502) );
  AOI22X1 U6647 ( .A(n10690), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[9] ), .D(n5505), .Y(n5503) );
  NAND2X1 U6649 ( .A(n5421), .B(n10693), .Y(n5505) );
  NAND2X1 U6651 ( .A(n5406), .B(n4802), .Y(n5441) );
  NOR2X1 U6652 ( .A(n10756), .B(n4817), .Y(n4802) );
  NOR2X1 U6653 ( .A(n10656), .B(n10707), .Y(n5439) );
  AOI22X1 U6654 ( .A(n10620), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[9] ), .D(n4701), .Y(n5493) );
  NAND2X1 U6655 ( .A(n5507), .B(n5508), .Y(n9105) );
  AOI22X1 U6656 ( .A(n5509), .B(n5510), .C(n10620), .D(n9364), .Y(n5508) );
  OAI21X1 U6657 ( .A(n9358), .B(n5511), .C(n5512), .Y(n5510) );
  AOI22X1 U6658 ( .A(n5513), .B(n5481), .C(n10673), .D(n9403), .Y(n5512) );
  OAI21X1 U6660 ( .A(n9387), .B(n5483), .C(n5515), .Y(n5514) );
  AOI22X1 U6661 ( .A(n5453), .B(n5516), .C(n10656), .D(n9481), .Y(n5515) );
  OAI22X1 U6662 ( .A(n9391), .B(n5455), .C(n10707), .D(n5517), .Y(n5516) );
  AOI22X1 U6663 ( .A(n10638), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[8] ), .D(n5519), .Y(n5517) );
  NAND2X1 U6665 ( .A(n5421), .B(n10641), .Y(n5519) );
  NAND2X1 U6668 ( .A(n5521), .B(n10709), .Y(n5455) );
  NOR2X1 U6669 ( .A(n10724), .B(n10656), .Y(n5453) );
  AOI22X1 U6670 ( .A(n10691), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[8] ), .D(n9408), .Y(n5507) );
  NAND2X1 U6671 ( .A(n5523), .B(n5524), .Y(n9106) );
  AOI22X1 U6672 ( .A(n5525), .B(n5526), .C(n10691), .D(n9364), .Y(n5524) );
  OAI21X1 U6673 ( .A(n9359), .B(n5527), .C(n5528), .Y(n5526) );
  AOI22X1 U6674 ( .A(n5529), .B(n5495), .C(n10742), .D(n9403), .Y(n5528) );
  OAI21X1 U6676 ( .A(n9387), .B(n5497), .C(n5531), .Y(n5530) );
  AOI22X1 U6677 ( .A(n5467), .B(n5532), .C(n10724), .D(n9481), .Y(n5531) );
  OAI22X1 U6678 ( .A(n9392), .B(n5469), .C(n10656), .D(n5533), .Y(n5532) );
  AOI22X1 U6679 ( .A(n10708), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[7] ), .D(n5535), .Y(n5533) );
  NAND2X1 U6681 ( .A(n5536), .B(n10709), .Y(n5535) );
  NAND2X1 U6684 ( .A(n5521), .B(n10658), .Y(n5469) );
  NOR2X1 U6685 ( .A(n10673), .B(n10724), .Y(n5467) );
  AOI22X1 U6686 ( .A(n10639), .B(n9416), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[7] ), .D(n9408), .Y(n5523) );
  NAND2X1 U6687 ( .A(n5538), .B(n5539), .Y(n9107) );
  AOI22X1 U6688 ( .A(n5540), .B(n5541), .C(n10639), .D(n9364), .Y(n5539) );
  OAI21X1 U6689 ( .A(n9359), .B(n5542), .C(n5543), .Y(n5541) );
  AOI22X1 U6690 ( .A(n5544), .B(n5509), .C(n10620), .D(n9403), .Y(n5543) );
  OAI21X1 U6692 ( .A(n9387), .B(n5511), .C(n5546), .Y(n5545) );
  AOI22X1 U6693 ( .A(n5481), .B(n5547), .C(n10673), .D(n9481), .Y(n5546) );
  OAI22X1 U6694 ( .A(n9392), .B(n5483), .C(n10724), .D(n5548), .Y(n5547) );
  AOI22X1 U6695 ( .A(n10657), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[6] ), .D(n5550), .Y(n5548) );
  NAND2X1 U6697 ( .A(n5536), .B(n10658), .Y(n5550) );
  NAND2X1 U6700 ( .A(n5521), .B(n10726), .Y(n5483) );
  NOR2X1 U6701 ( .A(n10742), .B(n10673), .Y(n5481) );
  AOI22X1 U6702 ( .A(n10710), .B(n9412), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[6] ), .D(n9408), .Y(n5538) );
  NAND2X1 U6703 ( .A(n5552), .B(n5553), .Y(n9108) );
  AOI22X1 U6704 ( .A(n5554), .B(n5555), .C(n10659), .D(n9412), .Y(n5553) );
  OAI21X1 U6705 ( .A(n9359), .B(n5557), .C(n5558), .Y(n5555) );
  AOI22X1 U6706 ( .A(n5559), .B(n5525), .C(n10691), .D(n9403), .Y(n5558) );
  OAI21X1 U6708 ( .A(n9387), .B(n5527), .C(n5561), .Y(n5560) );
  AOI22X1 U6709 ( .A(n5495), .B(n5562), .C(n10742), .D(n9481), .Y(n5561) );
  OAI22X1 U6710 ( .A(n9392), .B(n5497), .C(n10673), .D(n5563), .Y(n5562) );
  AOI22X1 U6711 ( .A(n10725), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[5] ), .D(n5565), .Y(n5563) );
  NAND2X1 U6713 ( .A(n5536), .B(n10726), .Y(n5565) );
  NAND2X1 U6716 ( .A(n5521), .B(n10675), .Y(n5497) );
  NOR2X1 U6717 ( .A(n10620), .B(n10742), .Y(n5495) );
  AOI22X1 U6718 ( .A(n10710), .B(n9364), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[5] ), .D(n9408), .Y(n5552) );
  NAND2X1 U6719 ( .A(n5566), .B(n5567), .Y(n9109) );
  AOI22X1 U6720 ( .A(n5568), .B(n5569), .C(n10727), .D(n9412), .Y(n5567) );
  OAI21X1 U6721 ( .A(n9359), .B(n5571), .C(n5572), .Y(n5569) );
  AOI22X1 U6722 ( .A(n5573), .B(n5540), .C(n10639), .D(n9403), .Y(n5572) );
  OAI21X1 U6724 ( .A(n9387), .B(n5542), .C(n5575), .Y(n5574) );
  AOI22X1 U6725 ( .A(n5509), .B(n5576), .C(n10620), .D(n9481), .Y(n5575) );
  OAI22X1 U6726 ( .A(n9392), .B(n5511), .C(n10742), .D(n5577), .Y(n5576) );
  AOI22X1 U6727 ( .A(n10674), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[4] ), .D(n5579), .Y(n5577) );
  NAND2X1 U6729 ( .A(n5536), .B(n10675), .Y(n5579) );
  NAND2X1 U6732 ( .A(n5521), .B(n10744), .Y(n5511) );
  NOR2X1 U6733 ( .A(n10691), .B(n10620), .Y(n5509) );
  AOI22X1 U6734 ( .A(n10659), .B(n9364), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[4] ), .D(n9408), .Y(n5566) );
  OAI21X1 U6736 ( .A(n9407), .B(n10788), .C(n5580), .Y(n9110) );
  AOI22X1 U6737 ( .A(n5581), .B(n5582), .C(n10676), .D(n9412), .Y(n5580) );
  OAI21X1 U6738 ( .A(n4676), .B(n5584), .C(n5585), .Y(n5581) );
  OAI21X1 U6739 ( .A(n5586), .B(n5587), .C(n5584), .Y(n5585) );
  OAI21X1 U6740 ( .A(n9164), .B(n5571), .C(n5589), .Y(n5587) );
  NAND3X1 U6741 ( .A(n9410), .B(n5590), .C(n5554), .Y(n5589) );
  OAI21X1 U6742 ( .A(n9387), .B(n5557), .C(n5591), .Y(n5590) );
  AOI22X1 U6743 ( .A(n5525), .B(n5592), .C(n10691), .D(n9481), .Y(n5591) );
  OAI22X1 U6744 ( .A(n9392), .B(n5527), .C(n10620), .D(n5593), .Y(n5592) );
  AOI22X1 U6745 ( .A(n10743), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[3] ), .D(n5595), .Y(n5593) );
  NAND2X1 U6747 ( .A(n5536), .B(n10744), .Y(n5595) );
  NAND2X1 U6750 ( .A(n5521), .B(n10622), .Y(n5527) );
  NOR2X1 U6751 ( .A(n10639), .B(n10691), .Y(n5525) );
  NOR2X1 U6752 ( .A(n9359), .B(n5596), .Y(n5586) );
  OAI21X1 U6754 ( .A(n9407), .B(n10786), .C(n5597), .Y(n9111) );
  AOI22X1 U6755 ( .A(n5598), .B(n5599), .C(n10745), .D(n9412), .Y(n5597) );
  OAI21X1 U6756 ( .A(n4676), .B(n5582), .C(n5601), .Y(n5598) );
  OAI21X1 U6757 ( .A(n5602), .B(n5603), .C(n5582), .Y(n5601) );
  OAI21X1 U6758 ( .A(n9164), .B(n5596), .C(n5604), .Y(n5603) );
  NAND3X1 U6759 ( .A(n9410), .B(n5605), .C(n5568), .Y(n5604) );
  OAI21X1 U6760 ( .A(n9387), .B(n5571), .C(n5606), .Y(n5605) );
  AOI22X1 U6761 ( .A(n5540), .B(n5607), .C(n10639), .D(n9481), .Y(n5606) );
  OAI22X1 U6762 ( .A(n9392), .B(n5542), .C(n10691), .D(n5608), .Y(n5607) );
  AOI22X1 U6763 ( .A(n10621), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[2] ), .D(n5610), .Y(n5608) );
  NAND2X1 U6765 ( .A(n5536), .B(n10622), .Y(n5610) );
  NAND2X1 U6768 ( .A(n5521), .B(n10693), .Y(n5542) );
  NOR2X1 U6769 ( .A(n10710), .B(n10639), .Y(n5540) );
  NOR2X1 U6770 ( .A(n9359), .B(n5584), .Y(n5602) );
  OAI21X1 U6773 ( .A(n9407), .B(n10784), .C(n5611), .Y(n9112) );
  AOI22X1 U6774 ( .A(n5612), .B(n5613), .C(n10623), .D(n9412), .Y(n5611) );
  OAI22X1 U6776 ( .A(n4676), .B(n5599), .C(n10745), .D(n5615), .Y(n5612) );
  AOI22X1 U6777 ( .A(n5616), .B(n5582), .C(n10676), .D(n4743), .Y(n5615) );
  NOR2X1 U6778 ( .A(n9409), .B(n10764), .Y(n4743) );
  OAI21X1 U6780 ( .A(n9164), .B(n5584), .C(n5617), .Y(n5616) );
  NAND3X1 U6781 ( .A(n5618), .B(n5584), .C(n9410), .Y(n5617) );
  OAI21X1 U6782 ( .A(n9383), .B(n5596), .C(n5619), .Y(n5618) );
  AOI22X1 U6783 ( .A(n5554), .B(n5620), .C(n10710), .D(n9481), .Y(n5619) );
  OAI22X1 U6784 ( .A(n9392), .B(n5557), .C(n10639), .D(n5621), .Y(n5620) );
  AOI22X1 U6785 ( .A(n10692), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[1] ), .D(n5623), .Y(n5621) );
  NAND2X1 U6787 ( .A(n5536), .B(n10693), .Y(n5623) );
  NAND2X1 U6790 ( .A(n5521), .B(n10641), .Y(n5557) );
  NOR2X1 U6793 ( .A(\U_0/U_0/U_1/U_8/address[6] ), .B(
        \U_0/U_0/U_1/U_8/address[7] ), .Y(n4930) );
  NOR2X1 U6794 ( .A(n10659), .B(n10710), .Y(n5554) );
  OAI21X1 U6799 ( .A(n9407), .B(n10782), .C(n5624), .Y(n9113) );
  AOI22X1 U6800 ( .A(n5625), .B(n5626), .C(n10694), .D(n9412), .Y(n5624) );
  NOR2X1 U6801 ( .A(n9409), .B(n10761), .Y(n4671) );
  NAND2X1 U6805 ( .A(n10754), .B(n4788), .Y(n5626) );
  NOR2X1 U6806 ( .A(n4803), .B(n10756), .Y(n4788) );
  NAND3X1 U6807 ( .A(n10751), .B(n10752), .C(\U_0/U_0/U_1/U_8/address[0] ), 
        .Y(n4803) );
  OAI22X1 U6808 ( .A(n5631), .B(n5632), .C(n4676), .D(n5613), .Y(n5625) );
  NAND2X1 U6809 ( .A(n9411), .B(\U_0/U_0/U_1/RCV_DATA [6]), .Y(n4676) );
  OAI21X1 U6810 ( .A(\U_0/U_0/U_1/RCV_DATA [5]), .B(n5599), .C(n9411), .Y(
        n5632) );
  NOR2X1 U6811 ( .A(n5633), .B(n9408), .Y(n4678) );
  OAI21X1 U6812 ( .A(n10745), .B(n5634), .C(n5613), .Y(n5631) );
  NAND2X1 U6813 ( .A(n10754), .B(n4768), .Y(n5613) );
  NOR2X1 U6814 ( .A(n4787), .B(n10756), .Y(n4768) );
  NAND3X1 U6815 ( .A(n10681), .B(n10752), .C(\U_0/U_0/U_1/U_8/address[1] ), 
        .Y(n4787) );
  AOI22X1 U6816 ( .A(n10676), .B(n10766), .C(n5636), .D(n5637), .Y(n5634) );
  AOI21X1 U6817 ( .A(n5568), .B(n5638), .C(n10676), .Y(n5637) );
  OAI22X1 U6818 ( .A(n9388), .B(n5571), .C(n10710), .D(n5639), .Y(n5638) );
  AOI22X1 U6819 ( .A(n10640), .B(n9486), .C(
        \U_0/U_0/U_1/U_8/currentPlainKey[0] ), .D(n5641), .Y(n5639) );
  NAND2X1 U6821 ( .A(n5536), .B(n10641), .Y(n5641) );
  NAND3X1 U6823 ( .A(n10751), .B(n10752), .C(n10681), .Y(n4817) );
  NOR2X1 U6825 ( .A(\U_0/U_0/U_1/U_8/address[4] ), .B(
        \U_0/U_0/U_1/U_8/address[5] ), .Y(n5520) );
  NAND2X1 U6827 ( .A(n10754), .B(n4946), .Y(n5571) );
  NOR2X1 U6828 ( .A(n4698), .B(n10756), .Y(n4946) );
  NAND3X1 U6829 ( .A(\U_0/U_0/U_1/U_8/address[1] ), .B(
        \U_0/U_0/U_1/U_8/address[0] ), .C(\U_0/U_0/U_1/U_8/address[2] ), .Y(
        n4698) );
  NOR2X1 U6831 ( .A(n10727), .B(n10659), .Y(n5568) );
  AOI22X1 U6832 ( .A(n10659), .B(n9481), .C(n10727), .D(
        \U_0/U_0/U_1/RCV_DATA [3]), .Y(n5636) );
  NAND2X1 U6834 ( .A(n10754), .B(n4716), .Y(n5584) );
  NOR2X1 U6835 ( .A(n4733), .B(n10756), .Y(n4716) );
  NAND3X1 U6836 ( .A(\U_0/U_0/U_1/U_8/address[0] ), .B(n10751), .C(
        \U_0/U_0/U_1/U_8/address[2] ), .Y(n4733) );
  NAND2X1 U6838 ( .A(n10754), .B(n4693), .Y(n5596) );
  NOR2X1 U6839 ( .A(n4713), .B(n10756), .Y(n4693) );
  NAND3X1 U6840 ( .A(\U_0/U_0/U_1/U_8/address[1] ), .B(n10681), .C(
        \U_0/U_0/U_1/U_8/address[2] ), .Y(n4713) );
  NAND2X1 U6843 ( .A(n10754), .B(n4730), .Y(n5582) );
  NOR2X1 U6844 ( .A(n4748), .B(n10756), .Y(n4730) );
  NAND3X1 U6845 ( .A(n10681), .B(n10751), .C(\U_0/U_0/U_1/U_8/address[2] ), 
        .Y(n4748) );
  NAND2X1 U6847 ( .A(n10754), .B(n4751), .Y(n5599) );
  NOR2X1 U6848 ( .A(n4767), .B(n10756), .Y(n4751) );
  NAND3X1 U6850 ( .A(\U_0/U_0/U_1/U_8/address[0] ), .B(n10752), .C(
        \U_0/U_0/U_1/U_8/address[1] ), .Y(n4767) );
  NAND3X1 U6852 ( .A(\U_0/U_0/U_1/U_8/address[6] ), .B(n4820), .C(
        \U_0/U_0/U_1/U_8/address[7] ), .Y(n5642) );
  NOR2X1 U6853 ( .A(n10758), .B(n10759), .Y(n4820) );
  NAND2X1 U6858 ( .A(n5643), .B(n10602), .Y(n4701) );
  OAI21X1 U6859 ( .A(n9207), .B(n10780), .C(n5647), .Y(n9114) );
  NAND2X1 U6860 ( .A(\U_0/U_0/U_1/U_8/N1799 ), .B(n5648), .Y(n5647) );
  OAI21X1 U6861 ( .A(n9207), .B(n10779), .C(n5650), .Y(n9115) );
  NAND2X1 U6862 ( .A(\U_0/U_0/U_1/U_8/N1798 ), .B(n5648), .Y(n5650) );
  OAI21X1 U6863 ( .A(n9207), .B(n10778), .C(n5652), .Y(n9116) );
  NAND2X1 U6864 ( .A(\U_0/U_0/U_1/U_8/N1797 ), .B(n5648), .Y(n5652) );
  OAI21X1 U6866 ( .A(n9207), .B(n10777), .C(n5654), .Y(n9117) );
  NAND2X1 U6867 ( .A(\U_0/U_0/U_1/U_8/N1796 ), .B(n5648), .Y(n5654) );
  OAI21X1 U6869 ( .A(n9207), .B(n10776), .C(n5656), .Y(n9118) );
  NAND2X1 U6870 ( .A(\U_0/U_0/U_1/U_8/N1795 ), .B(n5648), .Y(n5656) );
  OAI21X1 U6871 ( .A(n9207), .B(n10775), .C(n5658), .Y(n9119) );
  NAND2X1 U6872 ( .A(\U_0/U_0/U_1/U_8/N1794 ), .B(n5648), .Y(n5658) );
  OAI21X1 U6873 ( .A(n9207), .B(n10774), .C(n5660), .Y(n9120) );
  NAND2X1 U6874 ( .A(\U_0/U_0/U_1/U_8/N1793 ), .B(n5648), .Y(n5660) );
  OAI21X1 U6876 ( .A(n9207), .B(n10773), .C(n5662), .Y(n9121) );
  NAND2X1 U6877 ( .A(\U_0/U_0/U_1/U_8/N1792 ), .B(n5648), .Y(n5662) );
  OAI22X1 U6880 ( .A(n9206), .B(n10772), .C(n10770), .D(n5665), .Y(n9122) );
  OAI22X1 U6882 ( .A(n9206), .B(n10770), .C(n10769), .D(n5665), .Y(n9123) );
  OAI22X1 U6884 ( .A(n9206), .B(n10769), .C(n10767), .D(n5665), .Y(n9124) );
  OAI22X1 U6886 ( .A(n9206), .B(n10767), .C(n10765), .D(n5665), .Y(n9125) );
  OAI22X1 U6888 ( .A(n9206), .B(n10765), .C(n10763), .D(n5665), .Y(n9126) );
  OAI22X1 U6890 ( .A(n9206), .B(n10763), .C(n10762), .D(n5665), .Y(n9127) );
  OAI22X1 U6892 ( .A(n9206), .B(n10762), .C(n10760), .D(n5665), .Y(n9128) );
  OAI22X1 U6894 ( .A(n9206), .B(n10760), .C(n5665), .D(n10567), .Y(n9129) );
  OAI21X1 U6896 ( .A(n5668), .B(n10681), .C(n5669), .Y(n9130) );
  OAI21X1 U6898 ( .A(n5668), .B(n10751), .C(n5669), .Y(n9131) );
  OAI21X1 U6900 ( .A(n5668), .B(n10752), .C(n5669), .Y(n9132) );
  OAI21X1 U6902 ( .A(n10541), .B(n10606), .C(n5672), .Y(n9133) );
  AOI21X1 U6903 ( .A(\U_0/U_0/U_1/U_8/address[3] ), .B(n10541), .C(n10542), 
        .Y(n5672) );
  OAI21X1 U6904 ( .A(n10541), .B(n10603), .C(n5675), .Y(n9134) );
  AOI21X1 U6905 ( .A(\U_0/U_0/U_1/U_8/address[4] ), .B(n10541), .C(n10542), 
        .Y(n5675) );
  OAI21X1 U6906 ( .A(n10541), .B(n10604), .C(n5677), .Y(n9135) );
  AOI21X1 U6907 ( .A(\U_0/U_0/U_1/U_8/address[5] ), .B(n10541), .C(n10542), 
        .Y(n5677) );
  OAI21X1 U6910 ( .A(n5668), .B(n10753), .C(n5669), .Y(n9136) );
  OAI21X1 U6912 ( .A(n5668), .B(n10755), .C(n5669), .Y(n9137) );
  NAND2X1 U6913 ( .A(\U_0/U_0/U_1/U_8/keyCount[3] ), .B(n5668), .Y(n5669) );
  NOR2X1 U6915 ( .A(n5680), .B(n5681), .Y(n5668) );
  NAND3X1 U6916 ( .A(n5682), .B(n10600), .C(n7748), .Y(n5681) );
  NOR2X1 U6917 ( .A(n5663), .B(RST), .Y(n7748) );
  NAND3X1 U6918 ( .A(n5684), .B(n10602), .C(n5685), .Y(n5680) );
  OAI21X1 U6919 ( .A(n5686), .B(n5687), .C(n5688), .Y(n9138) );
  NAND2X1 U6920 ( .A(\U_0/U_0/U_1/U_8/keyCount[3] ), .B(n5689), .Y(n5688) );
  OAI21X1 U6921 ( .A(\U_0/U_0/U_1/U_8/keyCount[2] ), .B(n5633), .C(n5690), .Y(
        n5689) );
  OAI21X1 U6922 ( .A(n5690), .B(n10604), .C(n5691), .Y(n9139) );
  NAND3X1 U6923 ( .A(\U_0/U_0/U_1/U_8/keyCount[0] ), .B(n10604), .C(n5692), 
        .Y(n5691) );
  NOR2X1 U6924 ( .A(n10603), .B(n5687), .Y(n5692) );
  AOI21X1 U6926 ( .A(n10603), .B(n10590), .C(n5694), .Y(n5690) );
  OAI21X1 U6927 ( .A(n9722), .B(n10603), .C(n5696), .Y(n9140) );
  NAND3X1 U6928 ( .A(\U_0/U_0/U_1/U_8/keyCount[0] ), .B(n10603), .C(n9721), 
        .Y(n5696) );
  OAI21X1 U6932 ( .A(\U_0/U_0/U_1/U_8/keyCount[0] ), .B(n5633), .C(n5643), .Y(
        n5694) );
  OAI22X1 U6933 ( .A(n5643), .B(n10606), .C(\U_0/U_0/U_1/U_8/keyCount[0] ), 
        .D(n5687), .Y(n9141) );
  NAND2X1 U6934 ( .A(n10590), .B(n5643), .Y(n5687) );
  NOR2X1 U6936 ( .A(n5699), .B(n5700), .Y(n5645) );
  NAND3X1 U6937 ( .A(n5701), .B(n5685), .C(n10600), .Y(n5700) );
  NAND3X1 U6938 ( .A(n5684), .B(n9520), .C(n5702), .Y(n5699) );
  NAND3X1 U6939 ( .A(n5702), .B(n5633), .C(n5703), .Y(n9142) );
  AOI21X1 U6940 ( .A(\U_0/U_0/U_1/U_8/state[1] ), .B(n5704), .C(n10596), .Y(
        n5703) );
  OAI21X1 U6941 ( .A(n10588), .B(n10607), .C(n5698), .Y(n9143) );
  OAI21X1 U6943 ( .A(n5708), .B(n5709), .C(n5710), .Y(n5704) );
  OAI21X1 U6944 ( .A(n10609), .B(\U_0/U_0/U_1/U_8/keyCount[3] ), .C(n10598), 
        .Y(n5709) );
  NAND2X1 U6946 ( .A(n10610), .B(n10589), .Y(n5708) );
  NAND3X1 U6947 ( .A(n5716), .B(n5717), .C(n5718), .Y(n9144) );
  AOI21X1 U6948 ( .A(n10590), .B(n5686), .C(n5719), .Y(n5718) );
  OAI21X1 U6949 ( .A(n10597), .B(n5710), .C(n5721), .Y(n5719) );
  OAI21X1 U6950 ( .A(n10599), .B(n10596), .C(\U_0/RBUF_FULL ), .Y(n5721) );
  NAND3X1 U6952 ( .A(n10610), .B(n10589), .C(n10598), .Y(n5717) );
  NOR2X1 U6955 ( .A(n5723), .B(n5724), .Y(n5716) );
  OAI21X1 U6957 ( .A(\U_0/RBUF_FULL ), .B(n10602), .C(n10595), .Y(n5726) );
  OAI22X1 U6959 ( .A(n5710), .B(n10605), .C(n5686), .D(n5633), .Y(n5728) );
  NAND3X1 U6960 ( .A(\U_0/U_0/U_1/U_8/keyCount[2] ), .B(
        \U_0/U_0/U_1/U_8/keyCount[1] ), .C(n5730), .Y(n5686) );
  NOR2X1 U6961 ( .A(\U_0/U_0/U_1/U_8/keyCount[3] ), .B(n10606), .Y(n5730) );
  OAI21X1 U6963 ( .A(\U_0/U_0/U_1/U_8/state[3] ), .B(n5731), .C(n5732), .Y(
        n5710) );
  NAND3X1 U6965 ( .A(n10600), .B(n5701), .C(n5733), .Y(n5725) );
  OAI21X1 U6966 ( .A(\U_0/U_0/U_1/OE ), .B(\U_0/U_0/U_1/SBE ), .C(n10598), .Y(
        n5733) );
  OAI21X1 U6968 ( .A(n10568), .B(n5735), .C(n5736), .Y(n9146) );
  NAND3X1 U6969 ( .A(n5737), .B(n5738), .C(\U_0/U_0/U_1/SET_RBUF_FULL ), .Y(
        n5736) );
  XNOR2X1 U6970 ( .A(n10570), .B(\U_0/U_0/U_1/U_2/nextState[0] ), .Y(n5735) );
  OAI21X1 U6971 ( .A(n5740), .B(n10577), .C(n5738), .Y(n9147) );
  OAI21X1 U6972 ( .A(n5740), .B(n10578), .C(n5738), .Y(n9148) );
  NAND2X1 U6973 ( .A(n5737), .B(n5743), .Y(n5740) );
  OAI21X1 U6974 ( .A(n10570), .B(n5744), .C(n5745), .Y(n9149) );
  NAND3X1 U6975 ( .A(n5737), .B(n5738), .C(\U_0/U_0/U_1/RBUF_LOAD ), .Y(n5745)
         );
  NAND2X1 U6976 ( .A(\U_0/U_0/U_1/U_2/nextState[2] ), .B(n10560), .Y(n5744) );
  OAI21X1 U6977 ( .A(n10576), .B(n5748), .C(n5749), .Y(n9150) );
  NAND2X1 U6978 ( .A(n5737), .B(n5738), .Y(n5748) );
  OAI21X1 U6979 ( .A(n10587), .B(n5751), .C(n5743), .Y(n9151) );
  NAND3X1 U6980 ( .A(n10560), .B(n10568), .C(\U_0/U_0/U_1/U_2/nextState[1] ), 
        .Y(n5743) );
  NAND2X1 U6981 ( .A(n5749), .B(n5737), .Y(n5751) );
  NAND2X1 U6982 ( .A(\U_0/U_0/U_1/U_2/nextState[2] ), .B(n10570), .Y(n5749) );
  OAI21X1 U6983 ( .A(n5752), .B(n10571), .C(n5738), .Y(n9152) );
  NAND3X1 U6984 ( .A(n10570), .B(n10568), .C(\U_0/U_0/U_1/U_2/nextState[0] ), 
        .Y(n5738) );
  NAND3X1 U6986 ( .A(n10570), .B(n10568), .C(n10560), .Y(n5737) );
  OAI22X1 U6990 ( .A(n9206), .B(n10567), .C(n5665), .D(n10566), .Y(n9153) );
  OAI22X1 U6991 ( .A(n9206), .B(n10566), .C(n10543), .D(n5665), .Y(n9154) );
  OAI21X1 U6995 ( .A(n5755), .B(n5756), .C(n5757), .Y(n5665) );
  NOR2X1 U6996 ( .A(\U_0/U_0/U_1/U_7/state[7] ), .B(\U_0/U_0/U_1/U_7/state[0] ), .Y(n5757) );
  OAI21X1 U6997 ( .A(n10583), .B(n5759), .C(n5760), .Y(n5756) );
  NAND3X1 U6998 ( .A(\U_0/U_0/U_1/U_7/state[6] ), .B(
        \U_0/U_0/U_1/U_7/state[1] ), .C(n5761), .Y(n5760) );
  AOI21X1 U6999 ( .A(n5762), .B(n5763), .C(\U_0/U_0/U_1/U_7/state[3] ), .Y(
        n5761) );
  NAND3X1 U7000 ( .A(n10583), .B(n10565), .C(\U_0/U_0/U_1/U_7/state[4] ), .Y(
        n5763) );
  NAND3X1 U7002 ( .A(\U_0/U_0/U_1/U_7/state[2] ), .B(n10586), .C(
        \U_0/U_0/U_1/U_7/state[5] ), .Y(n5762) );
  NAND2X1 U7003 ( .A(\U_0/U_0/U_1/U_7/state[4] ), .B(n5766), .Y(n5759) );
  AOI21X1 U7004 ( .A(n10563), .B(n10583), .C(n5768), .Y(n5755) );
  NAND2X1 U7005 ( .A(n5769), .B(n10586), .Y(n5768) );
  OAI21X1 U7007 ( .A(n5770), .B(n5771), .C(\U_0/U_0/U_1/U_7/state[2] ), .Y(
        n5769) );
  NAND2X1 U7008 ( .A(\U_0/U_0/U_1/U_7/state[3] ), .B(n10581), .Y(n5771) );
  OAI21X1 U7013 ( .A(\U_0/U_0/U_1/U_7/state[6] ), .B(n5773), .C(n5774), .Y(
        n5766) );
  NAND3X1 U7014 ( .A(\U_0/U_0/U_1/U_7/state[3] ), .B(
        \U_0/U_0/U_1/U_7/state[6] ), .C(n5775), .Y(n5774) );
  NOR2X1 U7015 ( .A(\U_0/U_0/U_1/U_7/state[5] ), .B(\U_0/U_0/U_1/U_7/state[1] ), .Y(n5775) );
  AOI22X1 U7016 ( .A(n5776), .B(\U_0/U_0/U_1/U_7/state[1] ), .C(n5777), .D(
        \U_0/U_0/U_1/U_7/state[5] ), .Y(n5773) );
  XNOR2X1 U7017 ( .A(\U_0/U_0/U_1/U_7/state[1] ), .B(
        \U_0/U_0/U_1/U_7/state[3] ), .Y(n5777) );
  NOR2X1 U7018 ( .A(\U_0/U_0/U_1/U_7/state[5] ), .B(\U_0/U_0/U_1/U_7/state[3] ), .Y(n5776) );
  OAI21X1 U7019 ( .A(n10579), .B(n5779), .C(n5780), .Y(n9155) );
  NAND2X1 U7020 ( .A(\U_0/U_0/U_1/U_7/N26 ), .B(n5781), .Y(n5780) );
  OAI21X1 U7022 ( .A(n5779), .B(n10580), .C(n5783), .Y(n9156) );
  NAND2X1 U7023 ( .A(\U_0/U_0/U_1/U_7/N27 ), .B(n5781), .Y(n5783) );
  OAI21X1 U7024 ( .A(n10582), .B(n5779), .C(n5785), .Y(n9157) );
  NAND2X1 U7025 ( .A(\U_0/U_0/U_1/U_7/N28 ), .B(n5781), .Y(n5785) );
  OAI21X1 U7026 ( .A(n10584), .B(n5779), .C(n5787), .Y(n9158) );
  NAND2X1 U7027 ( .A(\U_0/U_0/U_1/U_7/N29 ), .B(n5781), .Y(n5787) );
  OAI21X1 U7028 ( .A(n5779), .B(n10585), .C(n5789), .Y(n9159) );
  NAND2X1 U7029 ( .A(\U_0/U_0/U_1/U_7/N30 ), .B(n5781), .Y(n5789) );
  OAI21X1 U7031 ( .A(n10564), .B(n5779), .C(n5791), .Y(n9160) );
  NAND2X1 U7032 ( .A(\U_0/U_0/U_1/U_7/N31 ), .B(n5781), .Y(n5791) );
  OAI21X1 U7034 ( .A(n10562), .B(n5779), .C(n5793), .Y(n9161) );
  NAND2X1 U7035 ( .A(\U_0/U_0/U_1/U_7/N32 ), .B(n5781), .Y(n5793) );
  OAI21X1 U7037 ( .A(n5779), .B(n10561), .C(n5795), .Y(n9162) );
  NAND2X1 U7038 ( .A(\U_0/U_0/U_1/U_7/N33 ), .B(n5781), .Y(n5795) );
  NAND2X1 U7041 ( .A(n10578), .B(n5796), .Y(n5779) );
  NAND3X1 U7043 ( .A(\U_0/U_0/U_1/U_7/nextState[6] ), .B(
        \U_0/U_0/U_1/U_7/nextState[5] ), .C(n5799), .Y(n5798) );
  NOR2X1 U7044 ( .A(n10582), .B(n10584), .Y(n5799) );
  NAND3X1 U7047 ( .A(\U_0/U_0/U_1/U_7/nextState[0] ), .B(n10580), .C(n5800), 
        .Y(n5797) );
  NOR2X1 U7048 ( .A(\U_0/U_0/U_1/U_7/nextState[7] ), .B(
        \U_0/U_0/U_1/U_7/nextState[4] ), .Y(n5800) );
  NAND2X1 U7051 ( .A(n5685), .B(n3184), .Y(c_prog_error) );
  NAND2X1 U7053 ( .A(n10592), .B(n11344), .Y(c_key_error) );
  NOR2X1 U7054 ( .A(n5803), .B(n5804), .Y(\U_1/U_3/U_4/nextcount [3]) );
  XNOR2X1 U7055 ( .A(\U_1/U_3/U_4/count[3] ), .B(n5805), .Y(n5803) );
  NOR2X1 U7056 ( .A(n5806), .B(n12071), .Y(n5805) );
  AOI21X1 U7057 ( .A(n5808), .B(\U_1/U_3/U_4/state ), .C(n11640), .Y(
        \U_1/U_3/U_4/nextcount [2]) );
  XNOR2X1 U7058 ( .A(n5806), .B(n12071), .Y(n5808) );
  NOR2X1 U7059 ( .A(n5804), .B(n5810), .Y(\U_1/U_3/U_4/nextcount [1]) );
  OAI21X1 U7060 ( .A(\U_1/U_3/U_4/count[1] ), .B(\U_1/U_3/U_4/count[0] ), .C(
        n5806), .Y(n5810) );
  NAND2X1 U7061 ( .A(\U_1/U_3/U_4/count[1] ), .B(\U_1/U_3/U_4/count[0] ), .Y(
        n5806) );
  NAND3X1 U7062 ( .A(n814), .B(slave_is_sending), .C(\U_1/U_3/U_4/state ), .Y(
        n5804) );
  NAND3X1 U7063 ( .A(n12072), .B(n12071), .C(n12070), .Y(n814) );
  OAI21X1 U7067 ( .A(\U_1/U_3/U_4/count[0] ), .B(n11640), .C(
        \U_1/U_3/U_4/state ), .Y(\U_1/U_3/U_4/nextcount [0]) );
  NAND3X1 U7069 ( .A(n191), .B(n5813), .C(n5814), .Y(slave_is_sending) );
  AOI21X1 U7070 ( .A(n190), .B(n11644), .C(n5815), .Y(n5814) );
  NOR2X1 U7072 ( .A(n11654), .B(n11648), .Y(n191) );
  NAND3X1 U7073 ( .A(n5816), .B(n11652), .C(n5817), .Y(
        \U_1/U_3/U_3/nextstate [2]) );
  AOI22X1 U7074 ( .A(n5818), .B(n5819), .C(n5820), .D(\U_1/PDATA_READY ), .Y(
        n5817) );
  NOR2X1 U7075 ( .A(\U_1/U_3/U_3/state[1] ), .B(\U_1/U_3/U_3/state[0] ), .Y(
        n5820) );
  NOR2X1 U7076 ( .A(n5821), .B(n11646), .Y(n5818) );
  NAND3X1 U7077 ( .A(n5822), .B(n5823), .C(n11647), .Y(
        \U_1/U_3/U_3/nextstate [1]) );
  OAI22X1 U7079 ( .A(n11932), .B(n5827), .C(n237), .D(n2004), .Y(n5825) );
  NAND3X1 U7080 ( .A(n11648), .B(n862), .C(\U_1/U_3/U_3/count[0] ), .Y(n5822)
         );
  OAI21X1 U7082 ( .A(n11932), .B(n5823), .C(n5813), .Y(n5829) );
  NAND3X1 U7085 ( .A(\U_1/U_3/U_3/state[0] ), .B(n11655), .C(
        \U_1/U_3/U_3/state[1] ), .Y(n237) );
  NAND2X1 U7086 ( .A(n5831), .B(n11654), .Y(n5823) );
  AOI22X1 U7088 ( .A(n5832), .B(n11868), .C(n5819), .D(n2004), .Y(n5831) );
  OAI21X1 U7090 ( .A(n11652), .B(n11646), .C(n5834), .Y(n5828) );
  OAI21X1 U7092 ( .A(n11645), .B(n11866), .C(n11648), .Y(n5835) );
  NAND3X1 U7094 ( .A(n11651), .B(n11655), .C(\U_1/U_3/U_3/state[0] ), .Y(n865)
         );
  NOR2X1 U7097 ( .A(n5838), .B(\U_1/U_3/U_3/N188 ), .Y(n862) );
  NOR2X1 U7099 ( .A(n5839), .B(n5840), .Y(n2004) );
  NAND3X1 U7100 ( .A(\U_1/U_3/U_3/count[4] ), .B(\U_1/U_3/U_3/count[1] ), .C(
        \U_1/U_3/U_3/count[5] ), .Y(n5840) );
  NAND3X1 U7101 ( .A(\U_1/U_3/U_3/count[0] ), .B(\U_1/U_3/U_3/count[3] ), .C(
        n5841), .Y(n5839) );
  NOR2X1 U7102 ( .A(\U_1/U_3/U_3/N188 ), .B(n11870), .Y(n5841) );
  NOR2X1 U7105 ( .A(n11653), .B(\U_1/U_3/U_3/state[0] ), .Y(n5815) );
  AOI21X1 U7106 ( .A(\U_1/U_3/U_0/state[3] ), .B(n5842), .C(n11642), .Y(
        \U_1/U_3/U_0/nextstate [3]) );
  NAND2X1 U7107 ( .A(n5843), .B(n5844), .Y(\U_1/U_3/U_0/nextstate [2]) );
  AOI22X1 U7108 ( .A(n5845), .B(n5846), .C(n11629), .D(n11628), .Y(n5843) );
  OAI21X1 U7112 ( .A(n11635), .B(n5849), .C(n5844), .Y(n5852) );
  AOI22X1 U7113 ( .A(n11623), .B(n5854), .C(n11642), .D(n11622), .Y(n5844) );
  OAI21X1 U7114 ( .A(n5856), .B(n5857), .C(n5858), .Y(n5851) );
  NAND3X1 U7115 ( .A(\U_1/U_3/U_0/state[1] ), .B(n5850), .C(n5859), .Y(n5858)
         );
  NOR2X1 U7116 ( .A(\U_1/U_3/U_0/state[3] ), .B(\U_1/U_3/U_0/state[0] ), .Y(
        n5859) );
  OAI21X1 U7117 ( .A(n5860), .B(n5861), .C(n11635), .Y(n5850) );
  NAND2X1 U7118 ( .A(\U_1/U_3/d_encode ), .B(n11642), .Y(n5861) );
  NAND2X1 U7119 ( .A(n5862), .B(n5863), .Y(\U_1/U_3/U_0/nextstate [0]) );
  AOI22X1 U7120 ( .A(n5854), .B(n5864), .C(n11621), .D(n11629), .Y(n5863) );
  NAND3X1 U7122 ( .A(\U_1/U_3/d_encode ), .B(n11633), .C(n11630), .Y(n5856) );
  XNOR2X1 U7124 ( .A(\U_1/U_3/U_0/DE_holdout_last ), .B(n11631), .Y(n5860) );
  AOI22X1 U7125 ( .A(n11622), .B(n11633), .C(n5868), .D(n11623), .Y(n5862) );
  OAI21X1 U7126 ( .A(n5869), .B(n785), .C(n5870), .Y(\U_1/U_3/U_0/dm_tx_nxt )
         );
  AOI22X1 U7127 ( .A(n5854), .B(n5871), .C(\U_1/U_3/U_0/state[3] ), .D(n5842), 
        .Y(n5870) );
  OAI21X1 U7128 ( .A(\U_1/U_3/U_0/N59 ), .B(n12077), .C(n5872), .Y(n5871) );
  OAI21X1 U7129 ( .A(n11622), .B(n784), .C(n11631), .Y(n5872) );
  AOI21X1 U7130 ( .A(n11622), .B(\U_1/U_3/U_0/DE_holdout ), .C(n5873), .Y(
        n5869) );
  OAI22X1 U7131 ( .A(n5874), .B(n12076), .C(\U_1/U_3/d_encode ), .D(n5876), 
        .Y(n5873) );
  AOI22X1 U7132 ( .A(\U_1/U_3/U_0/DE_holdout ), .B(n784), .C(
        \U_1/U_3/U_0/DE_holdout_BS ), .D(n11623), .Y(n5876) );
  AOI22X1 U7133 ( .A(n784), .B(n11631), .C(n11623), .D(n12077), .Y(n5874) );
  NAND3X1 U7138 ( .A(n11638), .B(n11627), .C(n11636), .Y(n5877) );
  NAND2X1 U7139 ( .A(n5857), .B(n5849), .Y(n5864) );
  NAND3X1 U7140 ( .A(\U_1/U_3/U_0/state[0] ), .B(\U_1/U_3/U_0/state[1] ), .C(
        n5880), .Y(n5849) );
  NOR2X1 U7141 ( .A(\U_1/U_3/U_0/state[3] ), .B(\U_1/U_3/U_0/state[2] ), .Y(
        n5880) );
  NAND2X1 U7142 ( .A(n5846), .B(\U_1/U_3/U_0/state[0] ), .Y(n5857) );
  NAND3X1 U7144 ( .A(n11638), .B(n11627), .C(n5882), .Y(n5881) );
  NAND3X1 U7145 ( .A(n5882), .B(n11627), .C(\U_1/U_3/U_0/state[0] ), .Y(
        \U_1/U_3/U_0/N59 ) );
  OAI21X1 U7147 ( .A(n5883), .B(n11636), .C(n5884), .Y(
        \U_1/U_3/U_0/DE_holdout_nxt ) );
  OAI21X1 U7149 ( .A(n11637), .B(n5846), .C(n5888), .Y(n5886) );
  OAI21X1 U7150 ( .A(n5889), .B(n11631), .C(n5890), .Y(n5888) );
  NAND3X1 U7151 ( .A(n11631), .B(n12076), .C(n11633), .Y(n5890) );
  AOI21X1 U7154 ( .A(\U_1/U_3/d_encode ), .B(n11642), .C(n5854), .Y(n5889) );
  NOR2X1 U7155 ( .A(\U_1/U_3/U_0/state[1] ), .B(\U_1/U_3/U_0/state[3] ), .Y(
        n5846) );
  OAI21X1 U7156 ( .A(n11642), .B(n5842), .C(\U_1/U_3/U_0/state[3] ), .Y(n5885)
         );
  NAND3X1 U7157 ( .A(n11639), .B(n11637), .C(n11638), .Y(n5842) );
  NOR2X1 U7160 ( .A(n11639), .B(n11637), .Y(n5882) );
  AOI22X1 U7163 ( .A(n5892), .B(n11642), .C(\U_1/U_3/U_0/state[0] ), .D(n5893), 
        .Y(n5883) );
  OAI21X1 U7164 ( .A(\U_1/U_3/U_0/DE_holdout_BS ), .B(n11634), .C(n5895), .Y(
        n5893) );
  NAND3X1 U7165 ( .A(\U_1/U_3/U_0/DE_holdout_BS ), .B(n11633), .C(
        \U_1/U_3/d_encode ), .Y(n5895) );
  NAND2X1 U7167 ( .A(\U_1/U_3/SHIFT_ENABLE_E ), .B(n11642), .Y(n785) );
  OAI21X1 U7169 ( .A(\U_1/U_3/d_encode ), .B(n5896), .C(n11635), .Y(n5868) );
  NOR2X1 U7171 ( .A(n5896), .B(\U_1/U_3/SHIFT_ENABLE_E ), .Y(n5854) );
  OAI21X1 U7173 ( .A(n5821), .B(n5897), .C(n5898), .Y(n5896) );
  NAND2X1 U7174 ( .A(\U_1/U_3/U_3/N187 ), .B(n11643), .Y(n5898) );
  OAI21X1 U7176 ( .A(n5899), .B(n5900), .C(n190), .Y(n5816) );
  NOR2X1 U7177 ( .A(n11656), .B(n11653), .Y(n190) );
  NOR2X1 U7179 ( .A(n11655), .B(\U_1/U_3/U_3/state[1] ), .Y(n877) );
  NAND3X1 U7180 ( .A(\U_1/U_3/U_3/count[2] ), .B(n5832), .C(
        \U_1/U_3/U_3/count[3] ), .Y(n5900) );
  NAND3X1 U7181 ( .A(n11872), .B(n11867), .C(n11869), .Y(n5899) );
  NAND2X1 U7185 ( .A(n5832), .B(n11868), .Y(n5897) );
  NAND3X1 U7187 ( .A(n5901), .B(n11871), .C(n5902), .Y(n5838) );
  NOR2X1 U7188 ( .A(\U_1/U_3/U_3/count[2] ), .B(\U_1/U_3/U_3/count[1] ), .Y(
        n5902) );
  NOR2X1 U7190 ( .A(\U_1/U_3/U_3/count[5] ), .B(\U_1/U_3/U_3/count[4] ), .Y(
        n5901) );
  NOR2X1 U7191 ( .A(n11644), .B(\U_1/U_3/U_3/count[0] ), .Y(n5832) );
  NOR2X1 U7193 ( .A(\U_1/U_3/U_0/state[0] ), .B(n5903), .Y(n5892) );
  XNOR2X1 U7194 ( .A(\U_1/U_3/SHIFT_ENABLE_E ), .B(\U_1/U_3/U_0/DE_holdout ), 
        .Y(n5903) );
  NOR2X1 U7195 ( .A(n5904), .B(n5905), .Y(\U_1/U_2/U_7/nextcount [3]) );
  NAND2X1 U7196 ( .A(n5906), .B(n5907), .Y(n5905) );
  XOR2X1 U7197 ( .A(\U_1/U_2/U_7/count[3] ), .B(n5908), .Y(n5906) );
  NOR2X1 U7198 ( .A(n5909), .B(n11560), .Y(n5908) );
  AOI21X1 U7199 ( .A(n5911), .B(n5912), .C(n5913), .Y(
        \U_1/U_2/U_7/nextcount [2]) );
  XNOR2X1 U7200 ( .A(n5909), .B(n11560), .Y(n5912) );
  NOR2X1 U7202 ( .A(n5904), .B(n5915), .Y(\U_1/U_2/U_7/nextcount [1]) );
  OAI21X1 U7203 ( .A(\U_1/U_2/U_7/count[1] ), .B(\U_1/U_2/U_7/count[0] ), .C(
        n5909), .Y(n5915) );
  NAND2X1 U7204 ( .A(\U_1/U_2/U_7/count[1] ), .B(\U_1/U_2/U_7/count[0] ), .Y(
        n5909) );
  OAI21X1 U7205 ( .A(n5913), .B(n5916), .C(\U_1/U_2/U_7/state ), .Y(
        \U_1/U_2/U_7/nextcount [0]) );
  NOR2X1 U7206 ( .A(n9715), .B(n11616), .Y(n5916) );
  NAND2X1 U7207 ( .A(n5919), .B(n5920), .Y(\U_1/U_2/U_5/nextstate [3]) );
  NOR2X1 U7208 ( .A(n5921), .B(n5922), .Y(n5920) );
  OAI21X1 U7209 ( .A(\U_1/U_2/U_5/state[1] ), .B(n5923), .C(n5924), .Y(n5922)
         );
  NAND3X1 U7210 ( .A(n5925), .B(n11555), .C(BSE_S), .Y(n5924) );
  AOI21X1 U7211 ( .A(\U_1/U_2/U_5/state[3] ), .B(n5927), .C(n5928), .Y(n5923)
         );
  OAI21X1 U7212 ( .A(n5929), .B(n5930), .C(n5931), .Y(n5928) );
  NAND3X1 U7213 ( .A(\U_1/U_2/U_5/state[0] ), .B(\U_1/U_2/U_5/state[2] ), .C(
        n9715), .Y(n5931) );
  NAND2X1 U7214 ( .A(n5932), .B(n9301), .Y(n5930) );
  OAI21X1 U7215 ( .A(n9301), .B(n5929), .C(n2112), .Y(n5927) );
  OAI21X1 U7216 ( .A(n11570), .B(n5934), .C(n5935), .Y(n5921) );
  NAND2X1 U7217 ( .A(n2016), .B(n11557), .Y(n5934) );
  AOI21X1 U7220 ( .A(n11553), .B(n9698), .C(n5937), .Y(n5919) );
  OAI22X1 U7221 ( .A(n9698), .B(n2110), .C(n5938), .D(n11569), .Y(n5937) );
  NAND3X1 U7222 ( .A(n11554), .B(n5941), .C(n5942), .Y(
        \U_1/U_2/U_5/nextstate [2]) );
  NOR2X1 U7223 ( .A(n5943), .B(n5944), .Y(n5942) );
  OAI22X1 U7224 ( .A(\U_1/U_2/U_5/N170 ), .B(n9204), .C(n9715), .D(n2114), .Y(
        n5944) );
  NAND3X1 U7225 ( .A(\U_1/U_2/U_5/state[2] ), .B(n11577), .C(n5932), .Y(n2114)
         );
  NAND3X1 U7226 ( .A(n5935), .B(n2130), .C(n5945), .Y(n5943) );
  OAI21X1 U7227 ( .A(n11551), .B(n11553), .C(n2142), .Y(n5945) );
  NAND2X1 U7229 ( .A(n9202), .B(n5948), .Y(n2130) );
  AOI22X1 U7230 ( .A(BSE_S), .B(n5949), .C(n11556), .D(n9698), .Y(n5941) );
  OAI21X1 U7233 ( .A(n11555), .B(n11577), .C(n2109), .Y(n5951) );
  AOI21X1 U7234 ( .A(n5925), .B(n2115), .C(n5952), .Y(n2109) );
  OAI22X1 U7235 ( .A(n9203), .B(n2016), .C(n5938), .D(n5953), .Y(n5952) );
  NOR2X1 U7236 ( .A(n5954), .B(\U_1/U_2/U_5/count[3] ), .Y(n2016) );
  NAND3X1 U7237 ( .A(\U_1/U_2/U_5/state[2] ), .B(n5955), .C(
        \U_1/U_2/U_5/state[1] ), .Y(n1888) );
  OAI21X1 U7239 ( .A(BSE_S), .B(n5956), .C(n5957), .Y(
        \U_1/U_2/U_5/nextstate [1]) );
  AOI21X1 U7240 ( .A(n9202), .B(n5958), .C(n11547), .Y(n5957) );
  NOR2X1 U7241 ( .A(n2034), .B(n5959), .Y(n5956) );
  OAI21X1 U7242 ( .A(n9202), .B(n5960), .C(n5947), .Y(n5959) );
  AOI22X1 U7243 ( .A(n11550), .B(n2142), .C(n11553), .D(n11572), .Y(n5960) );
  OAI21X1 U7245 ( .A(n5938), .B(n11569), .C(n5963), .Y(n2034) );
  OAI22X1 U7247 ( .A(n5964), .B(n5965), .C(n11577), .D(n5966), .Y(
        \U_1/U_2/U_5/nextstate [0]) );
  OAI21X1 U7248 ( .A(n11552), .B(n5968), .C(n5969), .Y(n5966) );
  NAND3X1 U7249 ( .A(n5929), .B(n9301), .C(n5970), .Y(n5969) );
  OAI21X1 U7250 ( .A(n11544), .B(n9698), .C(n5972), .Y(n5970) );
  AOI22X1 U7251 ( .A(n9697), .B(\U_1/U_2/U_5/state[3] ), .C(n5955), .D(n11569), 
        .Y(n5972) );
  NOR2X1 U7253 ( .A(n5974), .B(n5975), .Y(n5953) );
  NAND3X1 U7254 ( .A(n9317), .B(n9302), .C(n5976), .Y(n5975) );
  NOR2X1 U7255 ( .A(n9307), .B(n9305), .Y(n5976) );
  NAND3X1 U7257 ( .A(n9308), .B(n9310), .C(n5977), .Y(n5974) );
  NOR2X1 U7258 ( .A(n9315), .B(n9313), .Y(n5977) );
  NAND2X1 U7263 ( .A(\U_1/U_2/U_5/state[3] ), .B(\U_1/U_2/U_5/state[2] ), .Y(
        n5968) );
  OAI21X1 U7264 ( .A(\U_1/U_2/U_5/state[0] ), .B(n2112), .C(n5979), .Y(n5965)
         );
  NAND2X1 U7265 ( .A(n5980), .B(n11558), .Y(n5979) );
  OAI21X1 U7266 ( .A(n5978), .B(n5982), .C(n5983), .Y(n5980) );
  OAI21X1 U7267 ( .A(n9715), .B(n11552), .C(\U_1/U_2/U_5/state[2] ), .Y(n5983)
         );
  NAND2X1 U7269 ( .A(n5929), .B(n9301), .Y(n5982) );
  NAND3X1 U7270 ( .A(\U_1/U_2/U_5/state[0] ), .B(n9698), .C(n2142), .Y(n5978)
         );
  NOR2X1 U7271 ( .A(n11576), .B(n5954), .Y(n2142) );
  NAND3X1 U7272 ( .A(n11574), .B(n11575), .C(n11573), .Y(n5954) );
  NAND2X1 U7277 ( .A(n5914), .B(n9301), .Y(n2112) );
  OAI21X1 U7278 ( .A(n11552), .B(n5984), .C(n11577), .Y(n5964) );
  NAND2X1 U7279 ( .A(\U_1/U_2/U_5/state[3] ), .B(n5985), .Y(n5984) );
  OAI22X1 U7280 ( .A(n9301), .B(n9698), .C(\U_1/U_2/U_5/state[2] ), .D(n5914), 
        .Y(n5985) );
  OAI21X1 U7283 ( .A(n11565), .B(n9708), .C(n5929), .Y(n5986) );
  NAND3X1 U7284 ( .A(\U_1/U_2/U_1/state[3] ), .B(n11564), .C(n5989), .Y(n5929)
         );
  NOR2X1 U7285 ( .A(\U_1/U_2/U_1/state[2] ), .B(\U_1/U_2/U_1/state[1] ), .Y(
        n5989) );
  AOI21X1 U7287 ( .A(n9706), .B(n768), .C(n9202), .Y(\U_1/U_2/U_1/N31 ) );
  AOI22X1 U7288 ( .A(n2161), .B(n2164), .C(n9708), .D(n2155), .Y(n768) );
  OAI22X1 U7290 ( .A(n5992), .B(n9707), .C(n767), .D(n9708), .Y(n5991) );
  AOI21X1 U7291 ( .A(n5994), .B(n5995), .C(n9202), .Y(\U_1/U_2/U_1/N29 ) );
  AOI22X1 U7292 ( .A(n2163), .B(n2161), .C(n5996), .D(n2165), .Y(n5995) );
  OAI21X1 U7293 ( .A(\U_1/U_2/U_1/state[0] ), .B(n5992), .C(n774), .Y(n2165)
         );
  NAND2X1 U7294 ( .A(n5997), .B(n11564), .Y(n774) );
  NAND3X1 U7295 ( .A(n11568), .B(n11567), .C(\U_1/U_2/U_1/state[2] ), .Y(n5992) );
  NAND2X1 U7296 ( .A(n767), .B(n770), .Y(n2163) );
  NAND3X1 U7297 ( .A(n11568), .B(n11567), .C(\U_1/U_2/U_1/state[0] ), .Y(n770)
         );
  NAND3X1 U7299 ( .A(\U_1/U_2/U_1/state[0] ), .B(\U_1/U_2/U_1/state[1] ), .C(
        n5997), .Y(n767) );
  NOR2X1 U7300 ( .A(\U_1/U_2/U_1/state[2] ), .B(\U_1/U_2/U_1/state[3] ), .Y(
        n5997) );
  AOI22X1 U7301 ( .A(n9707), .B(n2155), .C(n2164), .D(n9708), .Y(n5994) );
  NOR2X1 U7303 ( .A(n2161), .B(n6000), .Y(n5996) );
  NOR2X1 U7304 ( .A(n11564), .B(n6001), .Y(n2164) );
  NOR2X1 U7306 ( .A(n6001), .B(\U_1/U_2/U_1/state[0] ), .Y(n2155) );
  NAND3X1 U7307 ( .A(\U_1/U_2/U_1/state[1] ), .B(n11567), .C(
        \U_1/U_2/U_1/state[2] ), .Y(n6001) );
  NAND2X1 U7310 ( .A(n9716), .B(n6000), .Y(n772) );
  XNOR2X1 U7311 ( .A(DPRS), .B(n11566), .Y(n6000) );
  NAND3X1 U7314 ( .A(n9718), .B(n11559), .C(\U_1/U_2/U_7/count[3] ), .Y(n2161)
         );
  NAND3X1 U7316 ( .A(n11617), .B(n11560), .C(n11616), .Y(n5907) );
  NAND3X1 U7321 ( .A(n11546), .B(n5914), .C(\U_1/U_2/U_7/state ), .Y(n5904) );
  NAND2X1 U7322 ( .A(n6005), .B(n9513), .Y(n5914) );
  XOR2X1 U7323 ( .A(\U_1/U_2/U_0/DP_hold2 ), .B(\U_1/U_2/U_0/DP_hold1 ), .Y(
        n6005) );
  NOR3X1 U7325 ( .A(n5958), .B(n11547), .C(n5949), .Y(n5913) );
  NAND3X1 U7326 ( .A(n5938), .B(n5963), .C(n11549), .Y(n5949) );
  NAND2X1 U7328 ( .A(n2108), .B(n5947), .Y(n5948) );
  NAND2X1 U7329 ( .A(n5932), .B(n5925), .Y(n5947) );
  NOR2X1 U7330 ( .A(n11550), .B(n11553), .Y(n2108) );
  NAND3X1 U7332 ( .A(\U_1/U_2/U_5/state[3] ), .B(n5925), .C(
        \U_1/U_2/U_5/state[0] ), .Y(n6006) );
  NAND3X1 U7334 ( .A(n11577), .B(n9301), .C(n5932), .Y(n6007) );
  NAND3X1 U7336 ( .A(\U_1/U_2/U_5/state[2] ), .B(n11577), .C(n2115), .Y(n5963)
         );
  NOR2X1 U7337 ( .A(n11558), .B(\U_1/U_2/U_5/state[0] ), .Y(n2115) );
  NAND2X1 U7338 ( .A(n5925), .B(n5955), .Y(n5938) );
  NOR2X1 U7339 ( .A(n11577), .B(\U_1/U_2/U_5/state[2] ), .Y(n5925) );
  NAND3X1 U7341 ( .A(\U_1/U_2/U_5/state[1] ), .B(\U_1/U_2/U_5/state[2] ), .C(
        n5932), .Y(n6008) );
  NOR2X1 U7342 ( .A(n11552), .B(\U_1/U_2/U_5/state[3] ), .Y(n5932) );
  NAND2X1 U7343 ( .A(n2110), .B(n5935), .Y(n5958) );
  NAND3X1 U7344 ( .A(\U_1/U_2/U_5/state[2] ), .B(n11577), .C(n6009), .Y(n5935)
         );
  NOR2X1 U7345 ( .A(n11558), .B(n11552), .Y(n6009) );
  NAND3X1 U7348 ( .A(n5955), .B(n11577), .C(\U_1/U_2/U_5/state[2] ), .Y(n2110)
         );
  NOR2X1 U7350 ( .A(\U_1/U_2/U_5/state[3] ), .B(\U_1/U_2/U_5/state[0] ), .Y(
        n5955) );
  NAND3X1 U7362 ( .A(n6010), .B(n6011), .C(n6012), .Y(
        \U_1/U_1/U_0/nextState [2]) );
  OAI21X1 U7363 ( .A(n11649), .B(n6014), .C(n11659), .Y(n6012) );
  NAND3X1 U7364 ( .A(n6016), .B(n11842), .C(\U_1/U_1/U_0/state[2] ), .Y(n6011)
         );
  OAI21X1 U7365 ( .A(n11830), .B(n6018), .C(\U_1/U_1/U_0/state[1] ), .Y(n6016)
         );
  NAND3X1 U7366 ( .A(\U_1/U_1/U_0/state[0] ), .B(n11657), .C(
        \U_1/U_1/U_0/state[1] ), .Y(n6010) );
  OAI21X1 U7367 ( .A(\U_1/U_1/U_0/state[2] ), .B(n11841), .C(n6019), .Y(
        \U_1/U_1/U_0/nextState [1]) );
  OAI21X1 U7368 ( .A(n6020), .B(n11659), .C(n11649), .Y(n6019) );
  OAI21X1 U7370 ( .A(\U_1/U_1/U_0/state[1] ), .B(n11842), .C(n6022), .Y(n6021)
         );
  OAI21X1 U7371 ( .A(\U_1/U_1/U_0/state[2] ), .B(n6022), .C(n6023), .Y(
        \U_1/U_1/U_0/nextState [0]) );
  AOI22X1 U7372 ( .A(n6024), .B(n6025), .C(n11658), .D(n6018), .Y(n6023) );
  AOI21X1 U7374 ( .A(n6014), .B(n11659), .C(n6020), .Y(n6027) );
  NOR2X1 U7375 ( .A(n6022), .B(n11830), .Y(n6020) );
  NAND3X1 U7377 ( .A(n6029), .B(n9643), .C(n6031), .Y(n6028) );
  NOR2X1 U7378 ( .A(\U_1/U_1/BYTE_COUNT [1]), .B(\U_1/U_1/BYTE_COUNT [0]), .Y(
        n6031) );
  NOR2X1 U7380 ( .A(\U_1/U_1/U_0/N39 ), .B(\U_1/U_1/BYTE_COUNT [3]), .Y(n6029)
         );
  NAND3X1 U7382 ( .A(\U_1/U_1/U_0/state[0] ), .B(n11843), .C(
        \U_1/U_1/U_0/state[2] ), .Y(n6032) );
  NAND2X1 U7384 ( .A(\U_1/U_1/OUT_OPCODE [0]), .B(\U_1/U_1/OUT_OPCODE [1]), 
        .Y(n6014) );
  OAI21X1 U7385 ( .A(n11649), .B(n6033), .C(n11657), .Y(n6025) );
  AOI21X1 U7387 ( .A(\U_1/U_1/U_0/N40 ), .B(n9202), .C(\U_1/U_1/U_0/N39 ), .Y(
        n6033) );
  NOR2X1 U7388 ( .A(DPRS), .B(DMRS), .Y(n2159) );
  OAI21X1 U7390 ( .A(n5819), .B(n5821), .C(n11650), .Y(n6018) );
  OAI22X1 U7392 ( .A(n11656), .B(n236), .C(\U_1/PDATA_READY ), .D(n5827), .Y(
        n6034) );
  NAND3X1 U7393 ( .A(n11651), .B(n11655), .C(n11656), .Y(n5827) );
  NAND2X1 U7395 ( .A(\U_1/U_3/U_3/state[1] ), .B(\U_1/U_3/U_3/state[2] ), .Y(
        n236) );
  NAND3X1 U7396 ( .A(n11656), .B(n11655), .C(\U_1/U_3/U_3/state[1] ), .Y(n5821) );
  NOR2X1 U7399 ( .A(\U_1/U_1/U_0/state[1] ), .B(\U_1/U_1/U_0/state[0] ), .Y(
        n6024) );
  NAND2X1 U7400 ( .A(\U_1/U_1/U_0/state[1] ), .B(n11842), .Y(n6022) );
  OAI21X1 U7402 ( .A(n11345), .B(n11533), .C(n6037), .Y(
        \U_1/U_0/U_1/U_8/nextParityError ) );
  OAI21X1 U7404 ( .A(n6040), .B(n6041), .C(n3223), .Y(n6038) );
  NAND3X1 U7405 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[0] ), .B(
        \U_1/U_0/U_1/U_8/parityAccumulator[1] ), .C(n6042), .Y(n6041) );
  NOR2X1 U7406 ( .A(n11528), .B(n11527), .Y(n6042) );
  NAND3X1 U7409 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[4] ), .B(
        \U_1/U_0/U_1/U_8/parityAccumulator[5] ), .C(n6043), .Y(n6040) );
  NOR2X1 U7410 ( .A(n11532), .B(n11531), .Y(n6043) );
  NOR2X1 U7414 ( .A(n6044), .B(n6045), .Y(\U_1/U_0/U_1/U_5/sb_detect_flag ) );
  NAND2X1 U7415 ( .A(\U_1/U_0/U_1/SBC_EN ), .B(n11329), .Y(n6045) );
  NOR2X1 U7416 ( .A(n11339), .B(n6046), .Y(\U_1/U_0/U_1/U_5/SBE_prime ) );
  NAND2X1 U7417 ( .A(n6044), .B(n11329), .Y(n6046) );
  NAND2X1 U7419 ( .A(\U_1/U_0/U_1/STOP_DATA [1]), .B(n11319), .Y(n6044) );
  OAI21X1 U7422 ( .A(n11326), .B(n11321), .C(n6049), .Y(
        \U_1/U_0/U_1/U_2/nextState[2] ) );
  AOI21X1 U7423 ( .A(n6050), .B(\U_1/U_0/U_1/U_2/state[1] ), .C(n6051), .Y(
        n6049) );
  OAI21X1 U7425 ( .A(n6052), .B(n11324), .C(n6054), .Y(
        \U_1/U_0/U_1/U_2/nextState[1] ) );
  NOR2X1 U7426 ( .A(n6055), .B(n6051), .Y(n6054) );
  NOR2X1 U7427 ( .A(n11326), .B(n6052), .Y(n6051) );
  OAI21X1 U7430 ( .A(\U_1/U_0/U_1/U_2/state[2] ), .B(n6056), .C(n11321), .Y(
        \U_1/U_0/U_1/U_2/nextState[0] ) );
  NOR2X1 U7432 ( .A(n11325), .B(\U_1/U_0/U_1/U_2/state[0] ), .Y(n6055) );
  AOI21X1 U7433 ( .A(\U_1/U_0/U_1/SB_DETECT ), .B(\U_1/U_0/U_1/U_2/state[1] ), 
        .C(n6058), .Y(n6056) );
  OAI21X1 U7434 ( .A(\U_1/U_0/U_1/U_2/N99 ), .B(n6052), .C(n6059), .Y(n6058)
         );
  NAND2X1 U7435 ( .A(n6060), .B(\U_1/U_0/U_1/U_0/Q_int2 ), .Y(n6059) );
  NOR2X1 U7436 ( .A(\U_1/U_0/U_1/U_2/state[0] ), .B(\U_1/U_0/U_1/U_0/Q_int ), 
        .Y(n6060) );
  NAND2X1 U7437 ( .A(\U_1/U_0/U_1/U_2/state[0] ), .B(n11325), .Y(n6052) );
  NOR2X1 U7448 ( .A(n11361), .B(n11328), .Y(\U_1/U_0/U_1/U_1/OE_prime ) );
  NOR2X1 U7451 ( .A(n6061), .B(n11909), .Y(n6958) );
  AOI22X1 U7453 ( .A(n9197), .B(\U_1/U_0/U_0/prefillCounter[7] ), .C(
        \U_1/U_0/U_0/extratemp[7] ), .D(n11918), .Y(n6063) );
  OAI21X1 U7454 ( .A(n11892), .B(n12033), .C(n6065), .Y(n6061) );
  AOI22X1 U7455 ( .A(n307), .B(DATA_IN_S[7]), .C(\U_1/U_0/U_0/fdata [7]), .D(
        n6066), .Y(n6065) );
  NOR2X1 U7456 ( .A(n6067), .B(n11908), .Y(n6957) );
  AOI22X1 U7458 ( .A(n9197), .B(\U_1/U_0/U_0/prefillCounter[6] ), .C(
        \U_1/U_0/U_0/extratemp[6] ), .D(n11918), .Y(n6069) );
  OAI21X1 U7459 ( .A(n11892), .B(n12030), .C(n6070), .Y(n6067) );
  AOI22X1 U7460 ( .A(n307), .B(DATA_IN_S[6]), .C(\U_1/U_0/U_0/fdata [6]), .D(
        n6066), .Y(n6070) );
  NOR2X1 U7461 ( .A(n6071), .B(n11907), .Y(n6956) );
  AOI22X1 U7463 ( .A(n9197), .B(\U_1/U_0/U_0/prefillCounter[5] ), .C(
        \U_1/U_0/U_0/extratemp[5] ), .D(n11918), .Y(n6073) );
  OAI21X1 U7464 ( .A(n11892), .B(n12027), .C(n6074), .Y(n6071) );
  AOI22X1 U7465 ( .A(n307), .B(DATA_IN_S[5]), .C(\U_1/U_0/U_0/fdata [5]), .D(
        n6066), .Y(n6074) );
  NOR2X1 U7466 ( .A(n6075), .B(n11906), .Y(n6955) );
  AOI22X1 U7468 ( .A(n9197), .B(\U_1/U_0/U_0/prefillCounter[4] ), .C(
        \U_1/U_0/U_0/extratemp[4] ), .D(n11918), .Y(n6077) );
  OAI21X1 U7469 ( .A(n11892), .B(n12024), .C(n6078), .Y(n6075) );
  AOI22X1 U7470 ( .A(n307), .B(DATA_IN_S[4]), .C(\U_1/U_0/U_0/fdata [4]), .D(
        n6066), .Y(n6078) );
  NOR2X1 U7471 ( .A(n6079), .B(n11905), .Y(n6954) );
  AOI22X1 U7473 ( .A(n9197), .B(\U_1/U_0/U_0/prefillCounter[3] ), .C(
        \U_1/U_0/U_0/extratemp[3] ), .D(n11918), .Y(n6081) );
  OAI21X1 U7474 ( .A(n11892), .B(n12022), .C(n6082), .Y(n6079) );
  AOI22X1 U7475 ( .A(n307), .B(DATA_IN_S[3]), .C(\U_1/U_0/U_0/fdata [3]), .D(
        n6066), .Y(n6082) );
  NOR2X1 U7476 ( .A(n6083), .B(n11904), .Y(n6953) );
  AOI22X1 U7478 ( .A(n9197), .B(\U_1/U_0/U_0/prefillCounter[2] ), .C(
        \U_1/U_0/U_0/extratemp[2] ), .D(n11918), .Y(n6085) );
  OAI21X1 U7479 ( .A(n11892), .B(n12020), .C(n6086), .Y(n6083) );
  AOI22X1 U7480 ( .A(n307), .B(DATA_IN_S[2]), .C(\U_1/U_0/U_0/fdata [2]), .D(
        n6066), .Y(n6086) );
  NOR2X1 U7481 ( .A(n6087), .B(n11903), .Y(n6952) );
  AOI22X1 U7483 ( .A(n9197), .B(\U_1/U_0/U_0/prefillCounter[1] ), .C(
        \U_1/U_0/U_0/extratemp[1] ), .D(n11918), .Y(n6089) );
  OAI21X1 U7484 ( .A(n11892), .B(n12018), .C(n6090), .Y(n6087) );
  AOI22X1 U7485 ( .A(n307), .B(DATA_IN_S[1]), .C(\U_1/U_0/U_0/fdata [1]), .D(
        n6066), .Y(n6090) );
  NOR2X1 U7486 ( .A(n6091), .B(n11902), .Y(n6951) );
  AOI22X1 U7488 ( .A(n9197), .B(\U_1/U_0/U_0/prefillCounter[0] ), .C(
        \U_1/U_0/U_0/extratemp[0] ), .D(n11918), .Y(n6093) );
  OAI21X1 U7489 ( .A(n11892), .B(n12016), .C(n6094), .Y(n6091) );
  AOI22X1 U7490 ( .A(n307), .B(DATA_IN_S[0]), .C(\U_1/U_0/U_0/fdata [0]), .D(
        n6066), .Y(n6094) );
  NAND3X1 U7491 ( .A(n11881), .B(n6095), .C(n11898), .Y(n6066) );
  NAND3X1 U7493 ( .A(n316), .B(n11912), .C(n6096), .Y(n300) );
  NOR2X1 U7494 ( .A(n6097), .B(n6098), .Y(n6096) );
  NAND3X1 U7497 ( .A(n1033), .B(n1016), .C(n6101), .Y(n6100) );
  AOI22X1 U7498 ( .A(n6102), .B(n6103), .C(n11920), .D(n9196), .Y(n6101) );
  NOR2X1 U7499 ( .A(n6106), .B(n6107), .Y(n6949) );
  NAND2X1 U7500 ( .A(n6108), .B(n6109), .Y(n6107) );
  AOI22X1 U7501 ( .A(\U_1/U_0/U_0/inti[7] ), .B(n956), .C(
        \U_1/U_0/U_0/intj[7] ), .D(n11914), .Y(n6109) );
  AOI22X1 U7502 ( .A(\U_1/U_0/U_0/N448 ), .B(n6110), .C(
        \U_1/U_0/U_0/prefillCounter[7] ), .D(n9197), .Y(n6108) );
  NAND2X1 U7503 ( .A(n6111), .B(n6112), .Y(n6106) );
  AOI22X1 U7504 ( .A(\U_1/U_0/U_0/N503 ), .B(n11899), .C(n6099), .D(
        \U_1/U_0/U_0/temp[7] ), .Y(n6112) );
  AOI22X1 U7505 ( .A(\U_1/U_0/U_0/sj[7] ), .B(n9199), .C(
        \U_1/U_0/U_0/faddr [7]), .D(n6113), .Y(n6111) );
  NOR2X1 U7506 ( .A(n6114), .B(n6115), .Y(n6948) );
  NAND2X1 U7507 ( .A(n6116), .B(n6117), .Y(n6115) );
  AOI22X1 U7508 ( .A(\U_1/U_0/U_0/inti[6] ), .B(n956), .C(
        \U_1/U_0/U_0/intj[6] ), .D(n11914), .Y(n6117) );
  AOI22X1 U7509 ( .A(\U_1/U_0/U_0/N447 ), .B(n6110), .C(
        \U_1/U_0/U_0/prefillCounter[6] ), .D(n9197), .Y(n6116) );
  NAND2X1 U7510 ( .A(n6118), .B(n6119), .Y(n6114) );
  AOI22X1 U7511 ( .A(\U_1/U_0/U_0/N502 ), .B(n11899), .C(\U_1/U_0/U_0/temp[6] ), .D(n6099), .Y(n6119) );
  AOI22X1 U7512 ( .A(\U_1/U_0/U_0/sj[6] ), .B(n9199), .C(
        \U_1/U_0/U_0/faddr [6]), .D(n6113), .Y(n6118) );
  NOR2X1 U7513 ( .A(n6120), .B(n6121), .Y(n6947) );
  NAND2X1 U7514 ( .A(n6122), .B(n6123), .Y(n6121) );
  AOI22X1 U7515 ( .A(\U_1/U_0/U_0/inti[5] ), .B(n956), .C(
        \U_1/U_0/U_0/intj[5] ), .D(n11914), .Y(n6123) );
  AOI22X1 U7516 ( .A(\U_1/U_0/U_0/N446 ), .B(n6110), .C(
        \U_1/U_0/U_0/prefillCounter[5] ), .D(n9197), .Y(n6122) );
  NAND2X1 U7517 ( .A(n6124), .B(n6125), .Y(n6120) );
  AOI22X1 U7518 ( .A(\U_1/U_0/U_0/N501 ), .B(n11899), .C(\U_1/U_0/U_0/temp[5] ), .D(n6099), .Y(n6125) );
  AOI22X1 U7519 ( .A(\U_1/U_0/U_0/sj[5] ), .B(n9199), .C(
        \U_1/U_0/U_0/faddr [5]), .D(n6113), .Y(n6124) );
  NOR2X1 U7520 ( .A(n6126), .B(n6127), .Y(n6946) );
  NAND2X1 U7521 ( .A(n6128), .B(n6129), .Y(n6127) );
  AOI22X1 U7522 ( .A(\U_1/U_0/U_0/inti[4] ), .B(n956), .C(
        \U_1/U_0/U_0/intj[4] ), .D(n11914), .Y(n6129) );
  AOI22X1 U7523 ( .A(\U_1/U_0/U_0/N445 ), .B(n6110), .C(
        \U_1/U_0/U_0/prefillCounter[4] ), .D(n9197), .Y(n6128) );
  NAND2X1 U7524 ( .A(n6130), .B(n6131), .Y(n6126) );
  AOI22X1 U7525 ( .A(\U_1/U_0/U_0/N500 ), .B(n11899), .C(\U_1/U_0/U_0/temp[4] ), .D(n6099), .Y(n6131) );
  AOI22X1 U7526 ( .A(\U_1/U_0/U_0/sj[4] ), .B(n9199), .C(
        \U_1/U_0/U_0/faddr [4]), .D(n6113), .Y(n6130) );
  NOR2X1 U7527 ( .A(n6132), .B(n6133), .Y(n6945) );
  NAND2X1 U7528 ( .A(n6134), .B(n6135), .Y(n6133) );
  AOI22X1 U7529 ( .A(\U_1/U_0/U_0/inti[3] ), .B(n956), .C(
        \U_1/U_0/U_0/intj[3] ), .D(n11914), .Y(n6135) );
  AOI22X1 U7530 ( .A(\U_1/U_0/U_0/N444 ), .B(n6110), .C(
        \U_1/U_0/U_0/prefillCounter[3] ), .D(n9197), .Y(n6134) );
  NAND2X1 U7531 ( .A(n6136), .B(n6137), .Y(n6132) );
  AOI22X1 U7532 ( .A(\U_1/U_0/U_0/N499 ), .B(n11899), .C(\U_1/U_0/U_0/temp[3] ), .D(n6099), .Y(n6137) );
  AOI22X1 U7533 ( .A(\U_1/U_0/U_0/sj[3] ), .B(n9199), .C(
        \U_1/U_0/U_0/faddr [3]), .D(n6113), .Y(n6136) );
  NOR2X1 U7534 ( .A(n6138), .B(n6139), .Y(n6944) );
  NAND2X1 U7535 ( .A(n6140), .B(n6141), .Y(n6139) );
  AOI22X1 U7536 ( .A(\U_1/U_0/U_0/inti[2] ), .B(n956), .C(
        \U_1/U_0/U_0/intj[2] ), .D(n11914), .Y(n6141) );
  AOI22X1 U7537 ( .A(\U_1/U_0/U_0/N443 ), .B(n6110), .C(
        \U_1/U_0/U_0/prefillCounter[2] ), .D(n9197), .Y(n6140) );
  NAND2X1 U7538 ( .A(n6142), .B(n6143), .Y(n6138) );
  AOI22X1 U7539 ( .A(\U_1/U_0/U_0/N498 ), .B(n11899), .C(\U_1/U_0/U_0/temp[2] ), .D(n6099), .Y(n6143) );
  AOI22X1 U7540 ( .A(\U_1/U_0/U_0/sj[2] ), .B(n9199), .C(
        \U_1/U_0/U_0/faddr [2]), .D(n6113), .Y(n6142) );
  NOR2X1 U7541 ( .A(n6144), .B(n6145), .Y(n6943) );
  NAND2X1 U7542 ( .A(n6146), .B(n6147), .Y(n6145) );
  AOI22X1 U7543 ( .A(\U_1/U_0/U_0/inti[1] ), .B(n956), .C(
        \U_1/U_0/U_0/intj[1] ), .D(n11914), .Y(n6147) );
  AOI22X1 U7544 ( .A(\U_1/U_0/U_0/N442 ), .B(n6110), .C(
        \U_1/U_0/U_0/prefillCounter[1] ), .D(n9197), .Y(n6146) );
  NAND2X1 U7545 ( .A(n6148), .B(n6149), .Y(n6144) );
  AOI22X1 U7546 ( .A(\U_1/U_0/U_0/N497 ), .B(n11899), .C(\U_1/U_0/U_0/temp[1] ), .D(n6099), .Y(n6149) );
  AOI22X1 U7547 ( .A(\U_1/U_0/U_0/sj[1] ), .B(n9199), .C(
        \U_1/U_0/U_0/faddr [1]), .D(n6113), .Y(n6148) );
  OAI21X1 U7549 ( .A(\U_1/U_0/U_0/state[3] ), .B(n11888), .C(n11898), .Y(n6150) );
  NAND3X1 U7551 ( .A(n1007), .B(n1008), .C(n6153), .Y(n6152) );
  NAND2X1 U7553 ( .A(n11901), .B(n6155), .Y(n1007) );
  NAND3X1 U7555 ( .A(n1098), .B(n980), .C(n1099), .Y(n1004) );
  NOR2X1 U7556 ( .A(n6157), .B(n6158), .Y(n6942) );
  NAND2X1 U7557 ( .A(n6159), .B(n6160), .Y(n6158) );
  AOI22X1 U7558 ( .A(\U_1/U_0/U_0/inti[0] ), .B(n956), .C(
        \U_1/U_0/U_0/intj[0] ), .D(n11914), .Y(n6160) );
  AOI22X1 U7559 ( .A(n11923), .B(n6110), .C(\U_1/U_0/U_0/prefillCounter[0] ), 
        .D(n9197), .Y(n6159) );
  NAND2X1 U7560 ( .A(n6161), .B(n6162), .Y(n6157) );
  AOI22X1 U7561 ( .A(\U_1/U_0/U_0/N496 ), .B(n11899), .C(\U_1/U_0/U_0/temp[0] ), .D(n6099), .Y(n6162) );
  AOI22X1 U7562 ( .A(\U_1/U_0/U_0/sj[0] ), .B(n9199), .C(
        \U_1/U_0/U_0/faddr [0]), .D(n6113), .Y(n6161) );
  NAND2X1 U7563 ( .A(n316), .B(n6095), .Y(n6113) );
  NOR2X1 U7564 ( .A(n918), .B(n11910), .Y(n316) );
  OAI21X1 U7565 ( .A(n11929), .B(n6165), .C(n6166), .Y(n918) );
  NOR2X1 U7566 ( .A(n11882), .B(n11915), .Y(n6166) );
  OAI21X1 U7569 ( .A(\U_1/U_0/U_0/state[3] ), .B(n11930), .C(n6170), .Y(n6168)
         );
  OAI21X1 U7570 ( .A(n931), .B(n6171), .C(n6172), .Y(n6167) );
  AOI21X1 U7571 ( .A(n11344), .B(n6173), .C(n11882), .Y(n6172) );
  OAI21X1 U7573 ( .A(n931), .B(n6174), .C(n6175), .Y(n6173) );
  OAI22X1 U7574 ( .A(n11844), .B(n11846), .C(n11911), .D(n11922), .Y(n6175) );
  NAND2X1 U7576 ( .A(n5819), .B(\U_1/B_READY ), .Y(n6174) );
  NAND3X1 U7577 ( .A(n6178), .B(n11894), .C(n6180), .Y(
        \U_1/U_0/U_0/nextState [3]) );
  AOI21X1 U7578 ( .A(n6181), .B(n6155), .C(n6182), .Y(n6180) );
  NAND2X1 U7579 ( .A(n320), .B(n1097), .Y(n6182) );
  NOR2X1 U7580 ( .A(n9286), .B(\U_1/U_0/U_0/state[1] ), .Y(n6181) );
  AOI22X1 U7581 ( .A(n11344), .B(n11910), .C(n6183), .D(n9196), .Y(n6178) );
  NAND3X1 U7582 ( .A(n6184), .B(n11894), .C(n6185), .Y(
        \U_1/U_0/U_0/nextState [2]) );
  AOI21X1 U7583 ( .A(n9196), .B(n11931), .C(n6187), .Y(n6185) );
  NAND2X1 U7584 ( .A(n322), .B(n6188), .Y(n6187) );
  OAI21X1 U7586 ( .A(n11924), .B(n1008), .C(n6191), .Y(n6189) );
  NOR2X1 U7587 ( .A(n11895), .B(n11899), .Y(n6191) );
  AOI22X1 U7590 ( .A(n11344), .B(n6192), .C(n6183), .D(n6193), .Y(n6184) );
  OAI22X1 U7591 ( .A(n6194), .B(n1096), .C(n11919), .D(n6196), .Y(n6192) );
  NAND3X1 U7592 ( .A(n11343), .B(n6198), .C(n6199), .Y(
        \U_1/U_0/U_0/nextState [1]) );
  NOR2X1 U7593 ( .A(n6200), .B(n6201), .Y(n6199) );
  OAI21X1 U7594 ( .A(n6202), .B(n6203), .C(n6204), .Y(n6201) );
  NAND3X1 U7595 ( .A(n6205), .B(n11934), .C(n6206), .Y(n6203) );
  NOR2X1 U7596 ( .A(\U_1/U_0/U_0/prefillCounter[2] ), .B(
        \U_1/U_0/U_0/prefillCounter[1] ), .Y(n6206) );
  NAND3X1 U7598 ( .A(n6207), .B(n11939), .C(n6208), .Y(n6202) );
  NOR2X1 U7599 ( .A(\U_1/U_0/U_0/prefillCounter[4] ), .B(
        \U_1/U_0/U_0/prefillCounter[3] ), .Y(n6208) );
  NOR2X1 U7601 ( .A(\U_1/U_0/U_0/prefillCounter[7] ), .B(
        \U_1/U_0/U_0/prefillCounter[6] ), .Y(n6207) );
  NAND2X1 U7602 ( .A(n1001), .B(n6165), .Y(n6200) );
  AOI22X1 U7603 ( .A(n6209), .B(n6210), .C(n6211), .D(n6212), .Y(n6198) );
  OAI21X1 U7604 ( .A(n11925), .B(n6171), .C(n11928), .Y(n6212) );
  OAI21X1 U7606 ( .A(n6216), .B(n5819), .C(\U_1/B_READY ), .Y(n6194) );
  NOR2X1 U7607 ( .A(n11916), .B(n6218), .Y(n6209) );
  OAI21X1 U7609 ( .A(n6171), .B(n11919), .C(n6220), .Y(n6219) );
  NAND2X1 U7611 ( .A(n6196), .B(n11344), .Y(n6171) );
  NOR2X1 U7612 ( .A(n6222), .B(n11844), .Y(n6196) );
  NAND3X1 U7615 ( .A(n318), .B(n9198), .C(n6220), .Y(n6224) );
  NOR2X1 U7616 ( .A(n6225), .B(n6226), .Y(n6220) );
  OAI21X1 U7617 ( .A(\U_1/U_0/U_0/permuteComplete ), .B(n1008), .C(n11892), 
        .Y(n6226) );
  OAI21X1 U7619 ( .A(n6227), .B(n11927), .C(n320), .Y(n308) );
  NAND3X1 U7620 ( .A(n980), .B(n6188), .C(n322), .Y(n6225) );
  NOR2X1 U7621 ( .A(n6205), .B(n11918), .Y(n318) );
  NAND3X1 U7622 ( .A(n1099), .B(n1097), .C(n6229), .Y(n6223) );
  OAI21X1 U7623 ( .A(n6230), .B(n6231), .C(n11344), .Y(n6229) );
  NAND3X1 U7625 ( .A(n6039), .B(n11352), .C(n11345), .Y(n6218) );
  NAND3X1 U7627 ( .A(n3181), .B(n11346), .C(n6234), .Y(n6232) );
  NOR2X1 U7628 ( .A(n11353), .B(n6236), .Y(n6234) );
  NAND2X1 U7629 ( .A(n3201), .B(n3183), .Y(n6236) );
  NAND3X1 U7630 ( .A(n6237), .B(n11357), .C(\U_1/U_0/U_1/U_8/state[0] ), .Y(
        n3183) );
  NAND3X1 U7633 ( .A(\U_1/U_0/U_1/U_8/state[2] ), .B(n11359), .C(n3230), .Y(
        n3184) );
  NAND2X1 U7635 ( .A(n3132), .B(n3197), .Y(n3162) );
  NAND3X1 U7636 ( .A(\U_1/U_0/U_1/U_8/state[0] ), .B(n6237), .C(
        \U_1/U_0/U_1/U_8/state[2] ), .Y(n3197) );
  NAND3X1 U7637 ( .A(n11349), .B(n11357), .C(n6237), .Y(n3132) );
  AOI21X1 U7638 ( .A(n11359), .B(n11351), .C(n11348), .Y(n3181) );
  NAND3X1 U7640 ( .A(n6237), .B(n11349), .C(\U_1/U_0/U_1/U_8/state[2] ), .Y(
        n3200) );
  NOR2X1 U7642 ( .A(n11360), .B(\U_1/U_0/U_1/U_8/state[3] ), .Y(n6237) );
  NOR2X1 U7645 ( .A(n11359), .B(n3231), .Y(n3223) );
  NAND2X1 U7646 ( .A(n3230), .B(n11357), .Y(n3231) );
  NOR2X1 U7647 ( .A(\U_1/U_0/U_1/U_8/state[1] ), .B(\U_1/U_0/U_1/U_8/state[0] ), .Y(n3230) );
  NAND2X1 U7648 ( .A(\U_1/U_0/U_1/U_8/parityError ), .B(n3222), .Y(n6039) );
  NOR2X1 U7649 ( .A(n6238), .B(n11357), .Y(n3222) );
  NAND3X1 U7651 ( .A(n11360), .B(n11359), .C(\U_1/U_0/U_1/U_8/state[0] ), .Y(
        n6238) );
  OAI22X1 U7654 ( .A(\U_1/U_0/U_0/state[3] ), .B(n6240), .C(\U_1/B_READY ), 
        .D(n1096), .Y(n6231) );
  OAI21X1 U7655 ( .A(n11846), .B(n6241), .C(n6242), .Y(n6230) );
  NAND3X1 U7656 ( .A(n6222), .B(n11845), .C(n11911), .Y(n6242) );
  NOR2X1 U7658 ( .A(n11847), .B(n11865), .Y(n5819) );
  NAND2X1 U7659 ( .A(n11865), .B(n11847), .Y(n6222) );
  NAND2X1 U7661 ( .A(\U_1/B_READY ), .B(n6221), .Y(n6241) );
  NOR2X1 U7663 ( .A(n11847), .B(\U_1/PRGA_OPCODE[1] ), .Y(n6216) );
  NOR2X1 U7665 ( .A(n6243), .B(n11886), .Y(n1097) );
  OAI21X1 U7666 ( .A(n11890), .B(n12034), .C(n6247), .Y(
        \U_1/U_0/U_0/nextProcessedData[7] ) );
  AOI22X1 U7667 ( .A(n6243), .B(n6248), .C(\U_1/PRGA_IN [7]), .D(n11886), .Y(
        n6247) );
  XNOR2X1 U7668 ( .A(n12033), .B(\U_1/U_0/U_0/delaydata [7]), .Y(n6248) );
  OAI21X1 U7671 ( .A(n11890), .B(n12031), .C(n6250), .Y(
        \U_1/U_0/U_0/nextProcessedData[6] ) );
  AOI22X1 U7672 ( .A(n6243), .B(n6251), .C(\U_1/PRGA_IN [6]), .D(n11886), .Y(
        n6250) );
  XNOR2X1 U7673 ( .A(n12030), .B(\U_1/U_0/U_0/delaydata [6]), .Y(n6251) );
  OAI21X1 U7676 ( .A(n11890), .B(n12028), .C(n6253), .Y(
        \U_1/U_0/U_0/nextProcessedData[5] ) );
  AOI22X1 U7677 ( .A(n6243), .B(n6254), .C(\U_1/PRGA_IN [5]), .D(n11886), .Y(
        n6253) );
  XNOR2X1 U7678 ( .A(n12027), .B(\U_1/U_0/U_0/delaydata [5]), .Y(n6254) );
  OAI21X1 U7681 ( .A(n11890), .B(n12025), .C(n6256), .Y(
        \U_1/U_0/U_0/nextProcessedData[4] ) );
  AOI22X1 U7682 ( .A(n6243), .B(n6257), .C(\U_1/PRGA_IN [4]), .D(n11886), .Y(
        n6256) );
  XNOR2X1 U7683 ( .A(n12024), .B(\U_1/U_0/U_0/delaydata [4]), .Y(n6257) );
  OAI21X1 U7686 ( .A(n11890), .B(n12023), .C(n6259), .Y(
        \U_1/U_0/U_0/nextProcessedData[3] ) );
  AOI22X1 U7687 ( .A(n6243), .B(n6260), .C(\U_1/PRGA_IN [3]), .D(n11886), .Y(
        n6259) );
  XNOR2X1 U7688 ( .A(n12022), .B(\U_1/U_0/U_0/delaydata [3]), .Y(n6260) );
  OAI21X1 U7691 ( .A(n11890), .B(n12021), .C(n6262), .Y(
        \U_1/U_0/U_0/nextProcessedData[2] ) );
  AOI22X1 U7692 ( .A(n6243), .B(n6263), .C(\U_1/PRGA_IN [2]), .D(n11886), .Y(
        n6262) );
  XNOR2X1 U7693 ( .A(n12020), .B(\U_1/U_0/U_0/delaydata [2]), .Y(n6263) );
  OAI21X1 U7696 ( .A(n11890), .B(n12019), .C(n6265), .Y(
        \U_1/U_0/U_0/nextProcessedData[1] ) );
  AOI22X1 U7697 ( .A(n6243), .B(n6266), .C(\U_1/PRGA_IN [1]), .D(n11886), .Y(
        n6265) );
  XNOR2X1 U7698 ( .A(n12018), .B(\U_1/U_0/U_0/delaydata [1]), .Y(n6266) );
  OAI21X1 U7701 ( .A(n11890), .B(n12017), .C(n6268), .Y(
        \U_1/U_0/U_0/nextProcessedData[0] ) );
  AOI22X1 U7702 ( .A(n6243), .B(n6269), .C(\U_1/PRGA_IN [0]), .D(n11886), .Y(
        n6268) );
  NAND2X1 U7704 ( .A(n11887), .B(n6215), .Y(n6204) );
  XNOR2X1 U7706 ( .A(n12016), .B(\U_1/U_0/U_0/delaydata [0]), .Y(n6269) );
  NAND3X1 U7711 ( .A(n6273), .B(n6274), .C(n6275), .Y(n6272) );
  NOR2X1 U7712 ( .A(n6276), .B(n6277), .Y(n6275) );
  NAND2X1 U7713 ( .A(n9200), .B(n912), .Y(n6277) );
  NAND2X1 U7714 ( .A(n6103), .B(n6193), .Y(n912) );
  OAI21X1 U7716 ( .A(n6227), .B(n11927), .C(n1033), .Y(n956) );
  NAND2X1 U7717 ( .A(n6278), .B(n6211), .Y(n1033) );
  NAND3X1 U7719 ( .A(n1001), .B(n322), .C(n1018), .Y(n6276) );
  NAND2X1 U7720 ( .A(n6278), .B(n6183), .Y(n1018) );
  NAND2X1 U7721 ( .A(n6099), .B(n9286), .Y(n322) );
  NAND3X1 U7722 ( .A(n9196), .B(n9286), .C(n6211), .Y(n1001) );
  NOR2X1 U7723 ( .A(n11910), .B(n6097), .Y(n6274) );
  NAND3X1 U7724 ( .A(n1098), .B(n321), .C(n1099), .Y(n6097) );
  NAND2X1 U7725 ( .A(n6278), .B(n6271), .Y(n1099) );
  NOR2X1 U7726 ( .A(n11928), .B(n11930), .Y(n6278) );
  NAND2X1 U7727 ( .A(n6102), .B(n11901), .Y(n321) );
  NAND3X1 U7728 ( .A(n9196), .B(n9286), .C(n6183), .Y(n1098) );
  NOR2X1 U7730 ( .A(n6221), .B(n11911), .Y(n921) );
  OAI21X1 U7732 ( .A(n6183), .B(n6211), .C(n6215), .Y(n1096) );
  NOR2X1 U7733 ( .A(n11930), .B(n11925), .Y(n6215) );
  NAND2X1 U7734 ( .A(n931), .B(n6177), .Y(n6221) );
  NAND3X1 U7735 ( .A(n6271), .B(n9286), .C(n6102), .Y(n6177) );
  NAND2X1 U7736 ( .A(n6102), .B(n11920), .Y(n931) );
  NOR2X1 U7737 ( .A(n11914), .B(n1054), .Y(n6273) );
  NAND3X1 U7738 ( .A(n1089), .B(n9168), .C(n6280), .Y(n1054) );
  NOR2X1 U7739 ( .A(n11896), .B(n11895), .Y(n6280) );
  NAND2X1 U7741 ( .A(n6102), .B(n6156), .Y(n980) );
  NAND2X1 U7743 ( .A(n6099), .B(n11930), .Y(n6188) );
  NOR2X1 U7744 ( .A(n11929), .B(n6227), .Y(n6099) );
  NAND2X1 U7747 ( .A(n6103), .B(n9196), .Y(n1016) );
  NAND2X1 U7748 ( .A(n6156), .B(n6155), .Y(n320) );
  NOR2X1 U7749 ( .A(n6227), .B(n9286), .Y(n6156) );
  NAND2X1 U7750 ( .A(\U_1/U_0/U_0/state[1] ), .B(n11917), .Y(n6227) );
  NOR2X1 U7751 ( .A(n6282), .B(n6283), .Y(n1089) );
  NAND3X1 U7752 ( .A(n6284), .B(n1008), .C(n9198), .Y(n6283) );
  OAI21X1 U7754 ( .A(n11929), .B(n6240), .C(n11921), .Y(n6110) );
  NOR2X1 U7756 ( .A(n6240), .B(n11925), .Y(n307) );
  NAND2X1 U7759 ( .A(n6103), .B(n6155), .Y(n1008) );
  OAI21X1 U7760 ( .A(n6155), .B(n9196), .C(n11901), .Y(n6284) );
  NOR2X1 U7762 ( .A(n11926), .B(\U_1/U_0/U_0/state[2] ), .Y(n6155) );
  NAND3X1 U7763 ( .A(n1020), .B(n11913), .C(n9179), .Y(n6282) );
  NAND2X1 U7767 ( .A(n6211), .B(n11930), .Y(n6165) );
  NOR2X1 U7768 ( .A(n11917), .B(\U_1/U_0/U_0/state[1] ), .Y(n6211) );
  NOR2X1 U7770 ( .A(n6095), .B(n11931), .Y(n6205) );
  NAND3X1 U7771 ( .A(n11917), .B(n11930), .C(n6193), .Y(n6095) );
  NAND2X1 U7772 ( .A(n11920), .B(n6193), .Y(n1020) );
  NOR2X1 U7773 ( .A(\U_1/U_0/U_0/state[2] ), .B(\U_1/U_0/U_0/state[3] ), .Y(
        n6193) );
  NAND2X1 U7775 ( .A(n6271), .B(n11930), .Y(n6240) );
  AOI21X1 U7778 ( .A(n6103), .B(n6102), .C(n11918), .Y(n6170) );
  NAND3X1 U7780 ( .A(n6271), .B(n9286), .C(n9196), .Y(n304) );
  NOR2X1 U7781 ( .A(n11933), .B(\U_1/U_0/U_0/state[3] ), .Y(n6105) );
  NOR2X1 U7782 ( .A(\U_1/U_0/U_0/state[0] ), .B(\U_1/U_0/U_0/state[1] ), .Y(
        n6271) );
  NOR2X1 U7783 ( .A(n11933), .B(n11926), .Y(n6102) );
  NOR2X1 U7786 ( .A(n11916), .B(n9286), .Y(n6103) );
  NOR2X1 U7788 ( .A(n11917), .B(n11931), .Y(n6183) );
  NAND3X1 U7791 ( .A(n6287), .B(n6288), .C(n6289), .Y(\U_1/U_0/U_0/N479 ) );
  NOR2X1 U7792 ( .A(n6290), .B(n6291), .Y(n6289) );
  OAI22X1 U7793 ( .A(n11967), .B(n6293), .C(n11948), .D(n6294), .Y(n6291) );
  OAI22X1 U7796 ( .A(n11951), .B(n6296), .C(n11959), .D(n6298), .Y(n6290) );
  AOI22X1 U7799 ( .A(n11981), .B(\U_1/U_0/U_0/keyTable[5][0] ), .C(n11980), 
        .D(\U_1/U_0/U_0/keyTable[4][0] ), .Y(n6288) );
  AOI22X1 U7800 ( .A(n11983), .B(\U_1/U_0/U_0/keyTable[7][0] ), .C(n11982), 
        .D(\U_1/U_0/U_0/keyTable[6][0] ), .Y(n6287) );
  NAND3X1 U7801 ( .A(n6303), .B(n6304), .C(n6305), .Y(\U_1/U_0/U_0/N478 ) );
  NOR2X1 U7802 ( .A(n6306), .B(n6307), .Y(n6305) );
  OAI22X1 U7803 ( .A(n11968), .B(n6293), .C(n11947), .D(n6294), .Y(n6307) );
  OAI22X1 U7806 ( .A(n11952), .B(n6296), .C(n11960), .D(n6298), .Y(n6306) );
  AOI22X1 U7809 ( .A(n11981), .B(\U_1/U_0/U_0/keyTable[5][1] ), .C(n11980), 
        .D(\U_1/U_0/U_0/keyTable[4][1] ), .Y(n6304) );
  AOI22X1 U7810 ( .A(n11983), .B(\U_1/U_0/U_0/keyTable[7][1] ), .C(n11982), 
        .D(\U_1/U_0/U_0/keyTable[6][1] ), .Y(n6303) );
  NAND3X1 U7811 ( .A(n6311), .B(n6312), .C(n6313), .Y(\U_1/U_0/U_0/N477 ) );
  NOR2X1 U7812 ( .A(n6314), .B(n6315), .Y(n6313) );
  OAI22X1 U7813 ( .A(n11969), .B(n6293), .C(n11946), .D(n6294), .Y(n6315) );
  OAI22X1 U7816 ( .A(n11953), .B(n6296), .C(n11961), .D(n6298), .Y(n6314) );
  AOI22X1 U7819 ( .A(n11981), .B(\U_1/U_0/U_0/keyTable[5][2] ), .C(n11980), 
        .D(\U_1/U_0/U_0/keyTable[4][2] ), .Y(n6312) );
  AOI22X1 U7820 ( .A(n11983), .B(\U_1/U_0/U_0/keyTable[7][2] ), .C(n11982), 
        .D(\U_1/U_0/U_0/keyTable[6][2] ), .Y(n6311) );
  NAND3X1 U7821 ( .A(n6319), .B(n6320), .C(n6321), .Y(\U_1/U_0/U_0/N476 ) );
  NOR2X1 U7822 ( .A(n6322), .B(n6323), .Y(n6321) );
  OAI22X1 U7823 ( .A(n11970), .B(n6293), .C(n11945), .D(n6294), .Y(n6323) );
  OAI22X1 U7826 ( .A(n11954), .B(n6296), .C(n11962), .D(n6298), .Y(n6322) );
  AOI22X1 U7829 ( .A(n11981), .B(\U_1/U_0/U_0/keyTable[5][3] ), .C(n11980), 
        .D(\U_1/U_0/U_0/keyTable[4][3] ), .Y(n6320) );
  AOI22X1 U7830 ( .A(n11983), .B(\U_1/U_0/U_0/keyTable[7][3] ), .C(n11982), 
        .D(\U_1/U_0/U_0/keyTable[6][3] ), .Y(n6319) );
  NAND3X1 U7831 ( .A(n6327), .B(n6328), .C(n6329), .Y(\U_1/U_0/U_0/N475 ) );
  NOR2X1 U7832 ( .A(n6330), .B(n6331), .Y(n6329) );
  OAI22X1 U7833 ( .A(n11971), .B(n6293), .C(n11944), .D(n6294), .Y(n6331) );
  OAI22X1 U7836 ( .A(n11955), .B(n6296), .C(n11963), .D(n6298), .Y(n6330) );
  AOI22X1 U7839 ( .A(n11981), .B(\U_1/U_0/U_0/keyTable[5][4] ), .C(n11980), 
        .D(\U_1/U_0/U_0/keyTable[4][4] ), .Y(n6328) );
  AOI22X1 U7840 ( .A(n11983), .B(\U_1/U_0/U_0/keyTable[7][4] ), .C(n11982), 
        .D(\U_1/U_0/U_0/keyTable[6][4] ), .Y(n6327) );
  NAND3X1 U7841 ( .A(n6336), .B(n6337), .C(n6338), .Y(\U_1/U_0/U_0/N474 ) );
  NOR2X1 U7842 ( .A(n6339), .B(n6340), .Y(n6338) );
  OAI22X1 U7843 ( .A(n11972), .B(n6293), .C(n11943), .D(n6294), .Y(n6340) );
  OAI22X1 U7846 ( .A(n11956), .B(n6296), .C(n11964), .D(n6298), .Y(n6339) );
  AOI22X1 U7849 ( .A(n11981), .B(\U_1/U_0/U_0/keyTable[5][5] ), .C(n11980), 
        .D(\U_1/U_0/U_0/keyTable[4][5] ), .Y(n6337) );
  AOI22X1 U7850 ( .A(n11983), .B(\U_1/U_0/U_0/keyTable[7][5] ), .C(n11982), 
        .D(\U_1/U_0/U_0/keyTable[6][5] ), .Y(n6336) );
  NAND3X1 U7851 ( .A(n6345), .B(n6346), .C(n6347), .Y(\U_1/U_0/U_0/N473 ) );
  NOR2X1 U7852 ( .A(n6348), .B(n6349), .Y(n6347) );
  OAI22X1 U7853 ( .A(n11973), .B(n6293), .C(n11942), .D(n6294), .Y(n6349) );
  OAI22X1 U7856 ( .A(n11957), .B(n6296), .C(n11965), .D(n6298), .Y(n6348) );
  AOI22X1 U7859 ( .A(n11981), .B(\U_1/U_0/U_0/keyTable[5][6] ), .C(n11980), 
        .D(\U_1/U_0/U_0/keyTable[4][6] ), .Y(n6346) );
  AOI22X1 U7860 ( .A(n11983), .B(\U_1/U_0/U_0/keyTable[7][6] ), .C(n11982), 
        .D(\U_1/U_0/U_0/keyTable[6][6] ), .Y(n6345) );
  NAND3X1 U7861 ( .A(n6354), .B(n6355), .C(n6356), .Y(\U_1/U_0/U_0/N472 ) );
  NOR2X1 U7862 ( .A(n6357), .B(n6358), .Y(n6356) );
  OAI22X1 U7863 ( .A(n11949), .B(n6293), .C(n11950), .D(n6294), .Y(n6358) );
  NAND3X1 U7864 ( .A(n11984), .B(n11979), .C(n12052), .Y(n6294) );
  NAND3X1 U7866 ( .A(n11984), .B(n11979), .C(\U_1/U_0/U_0/keyi[0] ), .Y(n6293)
         );
  OAI22X1 U7868 ( .A(n11958), .B(n6296), .C(n11966), .D(n6298), .Y(n6357) );
  NAND3X1 U7869 ( .A(n12052), .B(n11979), .C(\U_1/U_0/U_0/keyi[1] ), .Y(n6298)
         );
  NAND3X1 U7871 ( .A(\U_1/U_0/U_0/keyi[0] ), .B(n11979), .C(
        \U_1/U_0/U_0/keyi[1] ), .Y(n6296) );
  AOI22X1 U7874 ( .A(n11981), .B(\U_1/U_0/U_0/keyTable[5][7] ), .C(n11980), 
        .D(\U_1/U_0/U_0/keyTable[4][7] ), .Y(n6355) );
  NAND3X1 U7876 ( .A(n12052), .B(n11984), .C(\U_1/U_0/U_0/keyi[2] ), .Y(n6363)
         );
  NAND3X1 U7878 ( .A(\U_1/U_0/U_0/keyi[0] ), .B(n11984), .C(
        \U_1/U_0/U_0/keyi[2] ), .Y(n6364) );
  AOI22X1 U7880 ( .A(n11983), .B(\U_1/U_0/U_0/keyTable[7][7] ), .C(n11982), 
        .D(\U_1/U_0/U_0/keyTable[6][7] ), .Y(n6354) );
  NAND3X1 U7882 ( .A(\U_1/U_0/U_0/keyi[1] ), .B(n12052), .C(
        \U_1/U_0/U_0/keyi[2] ), .Y(n6365) );
  NAND3X1 U7885 ( .A(\U_1/U_0/U_0/keyi[1] ), .B(\U_1/U_0/U_0/keyi[0] ), .C(
        \U_1/U_0/U_0/keyi[2] ), .Y(n6366) );
  NOR2X1 U7886 ( .A(n6367), .B(n6368), .Y(\U_0/U_3/U_4/nextcount [3]) );
  XNOR2X1 U7887 ( .A(\U_0/U_3/U_4/count[3] ), .B(n6369), .Y(n6367) );
  NOR2X1 U7888 ( .A(n6370), .B(n11305), .Y(n6369) );
  AOI21X1 U7889 ( .A(n6372), .B(\U_0/U_3/U_4/state ), .C(n10888), .Y(
        \U_0/U_3/U_4/nextcount [2]) );
  XNOR2X1 U7890 ( .A(n6370), .B(n11305), .Y(n6372) );
  NOR2X1 U7891 ( .A(n6368), .B(n6374), .Y(\U_0/U_3/U_4/nextcount [1]) );
  OAI21X1 U7892 ( .A(\U_0/U_3/U_4/count[1] ), .B(\U_0/U_3/U_4/count[0] ), .C(
        n6370), .Y(n6374) );
  NAND2X1 U7893 ( .A(\U_0/U_3/U_4/count[1] ), .B(\U_0/U_3/U_4/count[0] ), .Y(
        n6370) );
  NAND3X1 U7894 ( .A(n3336), .B(host_is_sending), .C(\U_0/U_3/U_4/state ), .Y(
        n6368) );
  NAND3X1 U7895 ( .A(n11306), .B(n11305), .C(n11304), .Y(n3336) );
  OAI21X1 U7899 ( .A(\U_0/U_3/U_4/count[0] ), .B(n10888), .C(
        \U_0/U_3/U_4/state ), .Y(\U_0/U_3/U_4/nextcount [0]) );
  NAND3X1 U7901 ( .A(n6377), .B(n477), .C(n10890), .Y(host_is_sending) );
  OAI21X1 U7903 ( .A(n518), .B(\U_0/U_3/U_3/N188 ), .C(n519), .Y(n6379) );
  NOR2X1 U7904 ( .A(n10902), .B(n10896), .Y(n477) );
  NAND3X1 U7905 ( .A(n6380), .B(n519), .C(n6381), .Y(
        \U_0/U_3/U_3/nextstate [2]) );
  AOI22X1 U7906 ( .A(n6382), .B(n6383), .C(n6384), .D(\U_0/PDATA_READY ), .Y(
        n6381) );
  NOR2X1 U7907 ( .A(\U_0/U_3/U_3/state[1] ), .B(\U_0/U_3/U_3/state[0] ), .Y(
        n6384) );
  NOR2X1 U7908 ( .A(n6385), .B(n10894), .Y(n6382) );
  NAND3X1 U7909 ( .A(n6386), .B(n6387), .C(n10895), .Y(
        \U_0/U_3/U_3/nextstate [1]) );
  OAI22X1 U7911 ( .A(n11181), .B(n6391), .C(n522), .D(n4501), .Y(n6389) );
  NAND3X1 U7912 ( .A(n10896), .B(n3384), .C(\U_0/U_3/U_3/count[0] ), .Y(n6386)
         );
  OAI21X1 U7914 ( .A(n11181), .B(n6387), .C(n6377), .Y(n6393) );
  NAND2X1 U7916 ( .A(n3398), .B(n10904), .Y(n473) );
  NAND3X1 U7917 ( .A(\U_0/U_3/U_3/state[0] ), .B(n10903), .C(
        \U_0/U_3/U_3/state[1] ), .Y(n522) );
  NAND2X1 U7918 ( .A(n6395), .B(n10902), .Y(n6387) );
  AOI22X1 U7920 ( .A(n6396), .B(n11116), .C(n6383), .D(n4501), .Y(n6395) );
  OAI21X1 U7922 ( .A(n519), .B(n10894), .C(n6398), .Y(n6392) );
  OAI21X1 U7924 ( .A(n10893), .B(n11114), .C(n10896), .Y(n6399) );
  NAND3X1 U7926 ( .A(n10901), .B(n10903), .C(\U_0/U_3/U_3/state[0] ), .Y(n3387) );
  NOR2X1 U7929 ( .A(n6402), .B(\U_0/U_3/U_3/N188 ), .Y(n3384) );
  NOR2X1 U7931 ( .A(n6403), .B(n6404), .Y(n4501) );
  NAND3X1 U7932 ( .A(\U_0/U_3/U_3/count[4] ), .B(\U_0/U_3/U_3/count[1] ), .C(
        \U_0/U_3/U_3/count[5] ), .Y(n6404) );
  NAND3X1 U7933 ( .A(\U_0/U_3/U_3/count[0] ), .B(\U_0/U_3/U_3/count[3] ), .C(
        n6405), .Y(n6403) );
  NOR2X1 U7934 ( .A(\U_0/U_3/U_3/N188 ), .B(n11118), .Y(n6405) );
  NAND3X1 U7936 ( .A(n10904), .B(n10901), .C(\U_0/U_3/U_3/state[2] ), .Y(n519)
         );
  AOI21X1 U7937 ( .A(\U_0/U_3/U_0/state[3] ), .B(n6406), .C(n10891), .Y(
        \U_0/U_3/U_0/nextstate [3]) );
  NAND2X1 U7938 ( .A(n6407), .B(n6408), .Y(\U_0/U_3/U_0/nextstate [2]) );
  AOI22X1 U7939 ( .A(n6409), .B(n6410), .C(n10877), .D(n10876), .Y(n6407) );
  OAI21X1 U7943 ( .A(n10883), .B(n6413), .C(n6408), .Y(n6416) );
  AOI22X1 U7944 ( .A(n10871), .B(n6418), .C(n10891), .D(n10870), .Y(n6408) );
  OAI21X1 U7945 ( .A(n6420), .B(n6421), .C(n6422), .Y(n6415) );
  NAND3X1 U7946 ( .A(\U_0/U_3/U_0/state[1] ), .B(n6414), .C(n6423), .Y(n6422)
         );
  NOR2X1 U7947 ( .A(\U_0/U_3/U_0/state[3] ), .B(\U_0/U_3/U_0/state[0] ), .Y(
        n6423) );
  OAI21X1 U7948 ( .A(n6424), .B(n6425), .C(n10883), .Y(n6414) );
  NAND2X1 U7949 ( .A(\U_0/U_3/d_encode ), .B(n10891), .Y(n6425) );
  NAND2X1 U7950 ( .A(n6426), .B(n6427), .Y(\U_0/U_3/U_0/nextstate [0]) );
  AOI22X1 U7951 ( .A(n6418), .B(n6428), .C(n10869), .D(n10877), .Y(n6427) );
  NAND3X1 U7953 ( .A(\U_0/U_3/d_encode ), .B(n10881), .C(n10878), .Y(n6420) );
  XNOR2X1 U7955 ( .A(\U_0/U_3/U_0/DE_holdout_last ), .B(n10879), .Y(n6424) );
  AOI22X1 U7956 ( .A(n10870), .B(n10881), .C(n6432), .D(n10871), .Y(n6426) );
  OAI21X1 U7957 ( .A(n6433), .B(n3307), .C(n6434), .Y(\U_0/U_3/U_0/dm_tx_nxt )
         );
  AOI22X1 U7958 ( .A(n6418), .B(n6435), .C(\U_0/U_3/U_0/state[3] ), .D(n6406), 
        .Y(n6434) );
  OAI21X1 U7959 ( .A(\U_0/U_3/U_0/N59 ), .B(n11311), .C(n6436), .Y(n6435) );
  OAI21X1 U7960 ( .A(n10870), .B(n3306), .C(n10879), .Y(n6436) );
  AOI21X1 U7961 ( .A(n10870), .B(\U_0/U_3/U_0/DE_holdout ), .C(n6437), .Y(
        n6433) );
  OAI22X1 U7962 ( .A(n6438), .B(n11310), .C(\U_0/U_3/d_encode ), .D(n6440), 
        .Y(n6437) );
  AOI22X1 U7963 ( .A(\U_0/U_3/U_0/DE_holdout ), .B(n3306), .C(
        \U_0/U_3/U_0/DE_holdout_BS ), .D(n10871), .Y(n6440) );
  AOI22X1 U7964 ( .A(n3306), .B(n10879), .C(n10871), .D(n11311), .Y(n6438) );
  NAND3X1 U7969 ( .A(n10886), .B(n10875), .C(n10884), .Y(n6441) );
  NAND2X1 U7970 ( .A(n6421), .B(n6413), .Y(n6428) );
  NAND3X1 U7971 ( .A(\U_0/U_3/U_0/state[0] ), .B(\U_0/U_3/U_0/state[1] ), .C(
        n6444), .Y(n6413) );
  NOR2X1 U7972 ( .A(\U_0/U_3/U_0/state[3] ), .B(\U_0/U_3/U_0/state[2] ), .Y(
        n6444) );
  NAND2X1 U7973 ( .A(n6410), .B(\U_0/U_3/U_0/state[0] ), .Y(n6421) );
  NAND3X1 U7975 ( .A(n10886), .B(n10875), .C(n6446), .Y(n6445) );
  NAND3X1 U7976 ( .A(n6446), .B(n10875), .C(\U_0/U_3/U_0/state[0] ), .Y(
        \U_0/U_3/U_0/N59 ) );
  OAI21X1 U7978 ( .A(n6447), .B(n10884), .C(n6448), .Y(
        \U_0/U_3/U_0/DE_holdout_nxt ) );
  OAI21X1 U7980 ( .A(n10885), .B(n6410), .C(n6452), .Y(n6450) );
  OAI21X1 U7981 ( .A(n6453), .B(n10879), .C(n6454), .Y(n6452) );
  NAND3X1 U7982 ( .A(n10879), .B(n11310), .C(n10881), .Y(n6454) );
  AOI21X1 U7985 ( .A(\U_0/U_3/d_encode ), .B(n10891), .C(n6418), .Y(n6453) );
  NOR2X1 U7986 ( .A(\U_0/U_3/U_0/state[1] ), .B(\U_0/U_3/U_0/state[3] ), .Y(
        n6410) );
  OAI21X1 U7987 ( .A(n10891), .B(n6406), .C(\U_0/U_3/U_0/state[3] ), .Y(n6449)
         );
  NAND3X1 U7988 ( .A(n10887), .B(n10885), .C(n10886), .Y(n6406) );
  NOR2X1 U7991 ( .A(n10887), .B(n10885), .Y(n6446) );
  AOI22X1 U7994 ( .A(n6456), .B(n10891), .C(\U_0/U_3/U_0/state[0] ), .D(n6457), 
        .Y(n6447) );
  OAI21X1 U7995 ( .A(\U_0/U_3/U_0/DE_holdout_BS ), .B(n10882), .C(n6459), .Y(
        n6457) );
  NAND3X1 U7996 ( .A(\U_0/U_3/U_0/DE_holdout_BS ), .B(n10881), .C(
        \U_0/U_3/d_encode ), .Y(n6459) );
  NAND2X1 U7998 ( .A(\U_0/U_3/SHIFT_ENABLE_E ), .B(n10891), .Y(n3307) );
  OAI21X1 U8000 ( .A(\U_0/U_3/d_encode ), .B(n6460), .C(n10883), .Y(n6432) );
  NOR2X1 U8002 ( .A(n6460), .B(\U_0/U_3/SHIFT_ENABLE_E ), .Y(n6418) );
  OAI21X1 U8004 ( .A(n6385), .B(n6461), .C(n6462), .Y(n6460) );
  NAND2X1 U8005 ( .A(\U_0/U_3/U_3/N187 ), .B(n10892), .Y(n6462) );
  OAI21X1 U8007 ( .A(n6463), .B(n6464), .C(n10897), .Y(n6380) );
  NAND3X1 U8009 ( .A(\U_0/U_3/U_3/state[0] ), .B(n10901), .C(
        \U_0/U_3/U_3/state[2] ), .Y(n518) );
  NAND3X1 U8010 ( .A(\U_0/U_3/U_3/count[2] ), .B(n6396), .C(
        \U_0/U_3/U_3/count[3] ), .Y(n6464) );
  NAND3X1 U8011 ( .A(n11120), .B(n11115), .C(n11117), .Y(n6463) );
  NAND2X1 U8015 ( .A(n6396), .B(n11116), .Y(n6461) );
  NAND3X1 U8017 ( .A(n6465), .B(n11119), .C(n6466), .Y(n6402) );
  NOR2X1 U8018 ( .A(\U_0/U_3/U_3/count[2] ), .B(\U_0/U_3/U_3/count[1] ), .Y(
        n6466) );
  NOR2X1 U8020 ( .A(\U_0/U_3/U_3/count[5] ), .B(\U_0/U_3/U_3/count[4] ), .Y(
        n6465) );
  NOR2X1 U8021 ( .A(n9335), .B(\U_0/U_3/U_3/count[0] ), .Y(n6396) );
  NOR2X1 U8023 ( .A(\U_0/U_3/U_0/state[0] ), .B(n6467), .Y(n6456) );
  XNOR2X1 U8024 ( .A(\U_0/U_3/SHIFT_ENABLE_E ), .B(\U_0/U_3/U_0/DE_holdout ), 
        .Y(n6467) );
  NOR2X1 U8025 ( .A(n6468), .B(n6469), .Y(\U_0/U_2/U_7/nextcount [3]) );
  NAND2X1 U8026 ( .A(n6470), .B(n6471), .Y(n6469) );
  XOR2X1 U8027 ( .A(\U_0/U_2/U_7/count[3] ), .B(n6472), .Y(n6470) );
  NOR2X1 U8028 ( .A(n6473), .B(n10808), .Y(n6472) );
  AOI21X1 U8029 ( .A(n6475), .B(n6476), .C(n6477), .Y(
        \U_0/U_2/U_7/nextcount [2]) );
  XNOR2X1 U8030 ( .A(n6473), .B(n10808), .Y(n6476) );
  NOR2X1 U8032 ( .A(n6468), .B(n6479), .Y(\U_0/U_2/U_7/nextcount [1]) );
  OAI21X1 U8033 ( .A(\U_0/U_2/U_7/count[1] ), .B(\U_0/U_2/U_7/count[0] ), .C(
        n6473), .Y(n6479) );
  NAND2X1 U8034 ( .A(\U_0/U_2/U_7/count[1] ), .B(\U_0/U_2/U_7/count[0] ), .Y(
        n6473) );
  OAI21X1 U8035 ( .A(n6477), .B(n6480), .C(\U_0/U_2/U_7/state ), .Y(
        \U_0/U_2/U_7/nextcount [0]) );
  NOR2X1 U8036 ( .A(n9709), .B(n10864), .Y(n6480) );
  NAND2X1 U8037 ( .A(n6483), .B(n6484), .Y(\U_0/U_2/U_5/nextstate [3]) );
  NOR2X1 U8038 ( .A(n6485), .B(n6486), .Y(n6484) );
  OAI21X1 U8039 ( .A(\U_0/U_2/U_5/state[1] ), .B(n6487), .C(n6488), .Y(n6486)
         );
  NAND3X1 U8040 ( .A(n6489), .B(n10803), .C(BSE_H), .Y(n6488) );
  AOI21X1 U8041 ( .A(\U_0/U_2/U_5/state[3] ), .B(n6491), .C(n6492), .Y(n6487)
         );
  OAI21X1 U8042 ( .A(n6493), .B(n6494), .C(n6495), .Y(n6492) );
  NAND3X1 U8043 ( .A(\U_0/U_2/U_5/state[0] ), .B(\U_0/U_2/U_5/state[2] ), .C(
        n9709), .Y(n6495) );
  NAND2X1 U8044 ( .A(n6496), .B(n9336), .Y(n6494) );
  OAI21X1 U8045 ( .A(n9336), .B(n6493), .C(n4613), .Y(n6491) );
  OAI21X1 U8046 ( .A(n10818), .B(n6498), .C(n6499), .Y(n6485) );
  NAND2X1 U8047 ( .A(n4517), .B(n10805), .Y(n6498) );
  AOI21X1 U8050 ( .A(n10801), .B(n9690), .C(n6501), .Y(n6483) );
  OAI22X1 U8051 ( .A(n9690), .B(n4611), .C(n6502), .D(n10817), .Y(n6501) );
  NAND3X1 U8052 ( .A(n10802), .B(n6505), .C(n6506), .Y(
        \U_0/U_2/U_5/nextstate [2]) );
  NOR2X1 U8053 ( .A(n6507), .B(n6508), .Y(n6506) );
  OAI22X1 U8054 ( .A(\U_0/U_2/U_5/N170 ), .B(n9194), .C(n9709), .D(n4615), .Y(
        n6508) );
  NAND3X1 U8055 ( .A(\U_0/U_2/U_5/state[2] ), .B(n10825), .C(n6496), .Y(n4615)
         );
  NAND3X1 U8056 ( .A(n6499), .B(n4631), .C(n6509), .Y(n6507) );
  OAI21X1 U8057 ( .A(n10799), .B(n10801), .C(n4643), .Y(n6509) );
  NAND2X1 U8059 ( .A(n9192), .B(n6512), .Y(n4631) );
  AOI22X1 U8060 ( .A(BSE_H), .B(n6513), .C(n10804), .D(n9690), .Y(n6505) );
  OAI21X1 U8063 ( .A(n10803), .B(n10825), .C(n4610), .Y(n6515) );
  AOI21X1 U8064 ( .A(n6489), .B(n4616), .C(n6516), .Y(n4610) );
  OAI22X1 U8065 ( .A(n9193), .B(n4517), .C(n6502), .D(n6517), .Y(n6516) );
  NOR2X1 U8066 ( .A(n6518), .B(\U_0/U_2/U_5/count[3] ), .Y(n4517) );
  NAND3X1 U8067 ( .A(\U_0/U_2/U_5/state[2] ), .B(n6519), .C(
        \U_0/U_2/U_5/state[1] ), .Y(n4391) );
  OAI21X1 U8069 ( .A(BSE_H), .B(n6520), .C(n6521), .Y(
        \U_0/U_2/U_5/nextstate [1]) );
  AOI21X1 U8070 ( .A(n9192), .B(n6522), .C(n10795), .Y(n6521) );
  NOR2X1 U8071 ( .A(n4535), .B(n6523), .Y(n6520) );
  OAI21X1 U8072 ( .A(n9192), .B(n6524), .C(n6511), .Y(n6523) );
  AOI22X1 U8073 ( .A(n10798), .B(n4643), .C(n10801), .D(n10820), .Y(n6524) );
  OAI21X1 U8075 ( .A(n6502), .B(n10817), .C(n6527), .Y(n4535) );
  OAI22X1 U8077 ( .A(n6528), .B(n6529), .C(n10825), .D(n6530), .Y(
        \U_0/U_2/U_5/nextstate [0]) );
  OAI21X1 U8078 ( .A(n10800), .B(n6532), .C(n6533), .Y(n6530) );
  NAND3X1 U8079 ( .A(n6493), .B(n9336), .C(n6534), .Y(n6533) );
  OAI21X1 U8080 ( .A(n10792), .B(n9690), .C(n6536), .Y(n6534) );
  AOI22X1 U8081 ( .A(n9689), .B(\U_0/U_2/U_5/state[3] ), .C(n6519), .D(n10817), 
        .Y(n6536) );
  NOR2X1 U8083 ( .A(n6538), .B(n6539), .Y(n6517) );
  NAND3X1 U8084 ( .A(n9352), .B(n9337), .C(n6540), .Y(n6539) );
  NOR2X1 U8085 ( .A(n9342), .B(n9340), .Y(n6540) );
  NAND3X1 U8087 ( .A(n9343), .B(n9345), .C(n6541), .Y(n6538) );
  NOR2X1 U8088 ( .A(n9350), .B(n9348), .Y(n6541) );
  NAND2X1 U8093 ( .A(\U_0/U_2/U_5/state[3] ), .B(\U_0/U_2/U_5/state[2] ), .Y(
        n6532) );
  OAI21X1 U8094 ( .A(\U_0/U_2/U_5/state[0] ), .B(n4613), .C(n6543), .Y(n6529)
         );
  NAND2X1 U8095 ( .A(n6544), .B(n10806), .Y(n6543) );
  OAI21X1 U8096 ( .A(n6542), .B(n6546), .C(n6547), .Y(n6544) );
  OAI21X1 U8097 ( .A(n9709), .B(n10800), .C(\U_0/U_2/U_5/state[2] ), .Y(n6547)
         );
  NAND2X1 U8099 ( .A(n6493), .B(n9336), .Y(n6546) );
  NAND3X1 U8100 ( .A(\U_0/U_2/U_5/state[0] ), .B(n9690), .C(n4643), .Y(n6542)
         );
  NOR2X1 U8101 ( .A(n10824), .B(n6518), .Y(n4643) );
  NAND3X1 U8102 ( .A(n10822), .B(n10823), .C(n10821), .Y(n6518) );
  NAND2X1 U8107 ( .A(n6478), .B(n9336), .Y(n4613) );
  OAI21X1 U8108 ( .A(n10800), .B(n6548), .C(n10825), .Y(n6528) );
  NAND2X1 U8109 ( .A(\U_0/U_2/U_5/state[3] ), .B(n6549), .Y(n6548) );
  OAI22X1 U8110 ( .A(n9336), .B(n9690), .C(\U_0/U_2/U_5/state[2] ), .D(n6478), 
        .Y(n6549) );
  OAI21X1 U8113 ( .A(n10813), .B(n9705), .C(n6493), .Y(n6550) );
  NAND3X1 U8114 ( .A(\U_0/U_2/U_1/state[3] ), .B(n10812), .C(n6553), .Y(n6493)
         );
  NOR2X1 U8115 ( .A(\U_0/U_2/U_1/state[2] ), .B(\U_0/U_2/U_1/state[1] ), .Y(
        n6553) );
  AOI21X1 U8117 ( .A(n9703), .B(n754), .C(n9192), .Y(\U_0/U_2/U_1/N31 ) );
  AOI22X1 U8118 ( .A(n4662), .B(n4665), .C(n9705), .D(n4656), .Y(n754) );
  OAI22X1 U8120 ( .A(n6556), .B(n9704), .C(n753), .D(n9705), .Y(n6555) );
  AOI21X1 U8121 ( .A(n6558), .B(n6559), .C(n9192), .Y(\U_0/U_2/U_1/N29 ) );
  AOI22X1 U8122 ( .A(n4664), .B(n4662), .C(n6560), .D(n4666), .Y(n6559) );
  OAI21X1 U8123 ( .A(\U_0/U_2/U_1/state[0] ), .B(n6556), .C(n760), .Y(n4666)
         );
  NAND2X1 U8124 ( .A(n6561), .B(n10812), .Y(n760) );
  NAND3X1 U8125 ( .A(n10816), .B(n10815), .C(\U_0/U_2/U_1/state[2] ), .Y(n6556) );
  NAND2X1 U8126 ( .A(n753), .B(n756), .Y(n4664) );
  NAND3X1 U8127 ( .A(n10816), .B(n10815), .C(\U_0/U_2/U_1/state[0] ), .Y(n756)
         );
  NAND3X1 U8129 ( .A(\U_0/U_2/U_1/state[0] ), .B(\U_0/U_2/U_1/state[1] ), .C(
        n6561), .Y(n753) );
  NOR2X1 U8130 ( .A(\U_0/U_2/U_1/state[2] ), .B(\U_0/U_2/U_1/state[3] ), .Y(
        n6561) );
  AOI22X1 U8131 ( .A(n9704), .B(n4656), .C(n4665), .D(n9705), .Y(n6558) );
  NOR2X1 U8133 ( .A(n4662), .B(n6564), .Y(n6560) );
  NOR2X1 U8134 ( .A(n10812), .B(n6565), .Y(n4665) );
  NOR2X1 U8136 ( .A(n6565), .B(\U_0/U_2/U_1/state[0] ), .Y(n4656) );
  NAND3X1 U8137 ( .A(\U_0/U_2/U_1/state[1] ), .B(n10815), .C(
        \U_0/U_2/U_1/state[2] ), .Y(n6565) );
  NAND2X1 U8140 ( .A(n9710), .B(n6564), .Y(n758) );
  XNOR2X1 U8141 ( .A(DPRH), .B(n10814), .Y(n6564) );
  NAND3X1 U8144 ( .A(n9712), .B(n10807), .C(\U_0/U_2/U_7/count[3] ), .Y(n4662)
         );
  NAND3X1 U8146 ( .A(n10865), .B(n10808), .C(n10864), .Y(n6471) );
  NAND3X1 U8151 ( .A(n10794), .B(n6478), .C(\U_0/U_2/U_7/state ), .Y(n6468) );
  NAND2X1 U8152 ( .A(n6569), .B(n9514), .Y(n6478) );
  XOR2X1 U8154 ( .A(\U_0/U_2/U_0/DP_hold2 ), .B(\U_0/U_2/U_0/DP_hold1 ), .Y(
        n6569) );
  NOR3X1 U8156 ( .A(n6522), .B(n10795), .C(n6513), .Y(n6477) );
  NAND3X1 U8157 ( .A(n6502), .B(n6527), .C(n10797), .Y(n6513) );
  NAND2X1 U8159 ( .A(n4609), .B(n6511), .Y(n6512) );
  NAND2X1 U8160 ( .A(n6496), .B(n6489), .Y(n6511) );
  NOR2X1 U8161 ( .A(n10798), .B(n10801), .Y(n4609) );
  NAND3X1 U8163 ( .A(\U_0/U_2/U_5/state[3] ), .B(n6489), .C(
        \U_0/U_2/U_5/state[0] ), .Y(n6570) );
  NAND3X1 U8165 ( .A(n10825), .B(n9336), .C(n6496), .Y(n6571) );
  NAND3X1 U8167 ( .A(\U_0/U_2/U_5/state[2] ), .B(n10825), .C(n4616), .Y(n6527)
         );
  NOR2X1 U8168 ( .A(n10806), .B(\U_0/U_2/U_5/state[0] ), .Y(n4616) );
  NAND2X1 U8169 ( .A(n6489), .B(n6519), .Y(n6502) );
  NOR2X1 U8170 ( .A(n10825), .B(\U_0/U_2/U_5/state[2] ), .Y(n6489) );
  NAND3X1 U8172 ( .A(\U_0/U_2/U_5/state[1] ), .B(\U_0/U_2/U_5/state[2] ), .C(
        n6496), .Y(n6572) );
  NOR2X1 U8173 ( .A(n10800), .B(\U_0/U_2/U_5/state[3] ), .Y(n6496) );
  NAND2X1 U8174 ( .A(n4611), .B(n6499), .Y(n6522) );
  NAND3X1 U8175 ( .A(\U_0/U_2/U_5/state[2] ), .B(n10825), .C(n6573), .Y(n6499)
         );
  NOR2X1 U8176 ( .A(n10806), .B(n10800), .Y(n6573) );
  NAND3X1 U8179 ( .A(n6519), .B(n10825), .C(\U_0/U_2/U_5/state[2] ), .Y(n4611)
         );
  NOR2X1 U8181 ( .A(\U_0/U_2/U_5/state[3] ), .B(\U_0/U_2/U_5/state[0] ), .Y(
        n6519) );
  NAND3X1 U8193 ( .A(n6574), .B(n6575), .C(n6576), .Y(
        \U_0/U_1/U_0/nextState [2]) );
  OAI21X1 U8194 ( .A(n10899), .B(n6578), .C(n10907), .Y(n6576) );
  NAND3X1 U8195 ( .A(n6580), .B(n11090), .C(\U_0/U_1/U_0/state[2] ), .Y(n6575)
         );
  OAI21X1 U8196 ( .A(n11078), .B(n6582), .C(\U_0/U_1/U_0/state[1] ), .Y(n6580)
         );
  NAND3X1 U8197 ( .A(\U_0/U_1/U_0/state[0] ), .B(n10905), .C(
        \U_0/U_1/U_0/state[1] ), .Y(n6574) );
  OAI21X1 U8198 ( .A(\U_0/U_1/U_0/state[2] ), .B(n11089), .C(n6583), .Y(
        \U_0/U_1/U_0/nextState [1]) );
  OAI21X1 U8199 ( .A(n6584), .B(n10907), .C(n10899), .Y(n6583) );
  OAI21X1 U8201 ( .A(\U_0/U_1/U_0/state[1] ), .B(n11090), .C(n6586), .Y(n6585)
         );
  OAI21X1 U8202 ( .A(\U_0/U_1/U_0/state[2] ), .B(n6586), .C(n6587), .Y(
        \U_0/U_1/U_0/nextState [0]) );
  AOI22X1 U8203 ( .A(n6588), .B(n6589), .C(n10906), .D(n6582), .Y(n6587) );
  AOI21X1 U8205 ( .A(n6578), .B(n10907), .C(n6584), .Y(n6591) );
  NOR2X1 U8206 ( .A(n6586), .B(n11078), .Y(n6584) );
  NAND3X1 U8208 ( .A(n6593), .B(n9648), .C(n6595), .Y(n6592) );
  NOR2X1 U8209 ( .A(\U_0/U_1/BYTE_COUNT [1]), .B(\U_0/U_1/BYTE_COUNT [0]), .Y(
        n6595) );
  NOR2X1 U8211 ( .A(\U_0/U_1/U_0/N39 ), .B(\U_0/U_1/BYTE_COUNT [3]), .Y(n6593)
         );
  NAND3X1 U8213 ( .A(\U_0/U_1/U_0/state[0] ), .B(n11091), .C(
        \U_0/U_1/U_0/state[2] ), .Y(n6596) );
  NAND2X1 U8215 ( .A(\U_0/U_1/OUT_OPCODE [0]), .B(\U_0/U_1/OUT_OPCODE [1]), 
        .Y(n6578) );
  OAI21X1 U8216 ( .A(n10899), .B(n6597), .C(n10905), .Y(n6589) );
  AOI21X1 U8218 ( .A(\U_0/U_1/U_0/N40 ), .B(n9192), .C(\U_0/U_1/U_0/N39 ), .Y(
        n6597) );
  NOR2X1 U8219 ( .A(DPRH), .B(DMRH), .Y(n4660) );
  OAI21X1 U8221 ( .A(n6383), .B(n6385), .C(n6598), .Y(n6582) );
  AOI21X1 U8222 ( .A(n3398), .B(\U_0/U_3/U_3/state[0] ), .C(n3400), .Y(n6598)
         );
  NOR2X1 U8223 ( .A(n6391), .B(\U_0/PDATA_READY ), .Y(n3400) );
  NAND3X1 U8224 ( .A(n10901), .B(n10903), .C(n10904), .Y(n6391) );
  NOR2X1 U8225 ( .A(n10901), .B(n10903), .Y(n3398) );
  NAND3X1 U8227 ( .A(n10904), .B(n10903), .C(\U_0/U_3/U_3/state[1] ), .Y(n6385) );
  NOR2X1 U8230 ( .A(\U_0/U_1/U_0/state[1] ), .B(\U_0/U_1/U_0/state[0] ), .Y(
        n6588) );
  NAND2X1 U8231 ( .A(\U_0/U_1/U_0/state[1] ), .B(n11090), .Y(n6586) );
  OAI21X1 U8233 ( .A(n10593), .B(n10781), .C(n6601), .Y(
        \U_0/U_0/U_1/U_8/nextParityError ) );
  OAI21X1 U8235 ( .A(n6604), .B(n6605), .C(n5724), .Y(n6602) );
  NAND3X1 U8236 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[0] ), .B(
        \U_0/U_0/U_1/U_8/parityAccumulator[1] ), .C(n6606), .Y(n6605) );
  NOR2X1 U8237 ( .A(n10776), .B(n10775), .Y(n6606) );
  NAND3X1 U8240 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[4] ), .B(
        \U_0/U_0/U_1/U_8/parityAccumulator[5] ), .C(n6607), .Y(n6604) );
  NOR2X1 U8241 ( .A(n10780), .B(n10779), .Y(n6607) );
  NOR2X1 U8245 ( .A(n6608), .B(n6609), .Y(\U_0/U_0/U_1/U_5/sb_detect_flag ) );
  NAND2X1 U8246 ( .A(\U_0/U_0/U_1/SBC_EN ), .B(n10577), .Y(n6609) );
  NOR2X1 U8247 ( .A(n10587), .B(n6610), .Y(\U_0/U_0/U_1/U_5/SBE_prime ) );
  NAND2X1 U8248 ( .A(n6608), .B(n10577), .Y(n6610) );
  NAND2X1 U8250 ( .A(\U_0/U_0/U_1/STOP_DATA [1]), .B(n10567), .Y(n6608) );
  OAI21X1 U8253 ( .A(n10574), .B(n10569), .C(n6613), .Y(
        \U_0/U_0/U_1/U_2/nextState[2] ) );
  AOI21X1 U8254 ( .A(n6614), .B(\U_0/U_0/U_1/U_2/state[1] ), .C(n6615), .Y(
        n6613) );
  OAI21X1 U8256 ( .A(n6616), .B(n10572), .C(n6618), .Y(
        \U_0/U_0/U_1/U_2/nextState[1] ) );
  NOR2X1 U8257 ( .A(n6619), .B(n6615), .Y(n6618) );
  NOR2X1 U8258 ( .A(n10574), .B(n6616), .Y(n6615) );
  OAI21X1 U8261 ( .A(\U_0/U_0/U_1/U_2/state[2] ), .B(n6620), .C(n10569), .Y(
        \U_0/U_0/U_1/U_2/nextState[0] ) );
  NOR2X1 U8263 ( .A(n10573), .B(\U_0/U_0/U_1/U_2/state[0] ), .Y(n6619) );
  AOI21X1 U8264 ( .A(\U_0/U_0/U_1/SB_DETECT ), .B(\U_0/U_0/U_1/U_2/state[1] ), 
        .C(n6622), .Y(n6620) );
  OAI21X1 U8265 ( .A(\U_0/U_0/U_1/U_2/N99 ), .B(n6616), .C(n6623), .Y(n6622)
         );
  NAND2X1 U8266 ( .A(n6624), .B(\U_0/U_0/U_1/U_0/Q_int2 ), .Y(n6623) );
  NOR2X1 U8267 ( .A(\U_0/U_0/U_1/U_2/state[0] ), .B(\U_0/U_0/U_1/U_0/Q_int ), 
        .Y(n6624) );
  NAND2X1 U8268 ( .A(\U_0/U_0/U_1/U_2/state[0] ), .B(n10573), .Y(n6616) );
  NOR2X1 U8279 ( .A(n10609), .B(n10576), .Y(\U_0/U_0/U_1/U_1/OE_prime ) );
  NOR2X1 U8283 ( .A(n6626), .B(n6627), .Y(n6940) );
  OAI22X1 U8284 ( .A(n11155), .B(n11172), .C(n11137), .D(n11205), .Y(n6627) );
  OAI21X1 U8286 ( .A(n11129), .B(n11254), .C(n6630), .Y(n6626) );
  AOI22X1 U8287 ( .A(n9188), .B(DATA_IN_H[7]), .C(n11163), .D(
        \U_0/U_0/U_0/extratemp[7] ), .Y(n6630) );
  NOR2X1 U8289 ( .A(n6633), .B(n6634), .Y(n6939) );
  OAI22X1 U8290 ( .A(n11155), .B(n11180), .C(n11137), .D(n11198), .Y(n6634) );
  OAI21X1 U8292 ( .A(n11129), .B(n11234), .C(n6635), .Y(n6633) );
  AOI22X1 U8293 ( .A(n9188), .B(DATA_IN_H[6]), .C(n11163), .D(
        \U_0/U_0/U_0/extratemp[6] ), .Y(n6635) );
  NOR2X1 U8295 ( .A(n6636), .B(n6637), .Y(n6938) );
  OAI22X1 U8296 ( .A(n11155), .B(n11179), .C(n11137), .D(n11204), .Y(n6637) );
  OAI21X1 U8297 ( .A(n11129), .B(n11235), .C(n6638), .Y(n6636) );
  AOI22X1 U8298 ( .A(n9188), .B(DATA_IN_H[5]), .C(n11163), .D(
        \U_0/U_0/U_0/extratemp[5] ), .Y(n6638) );
  NOR2X1 U8300 ( .A(n6639), .B(n6640), .Y(n6937) );
  OAI22X1 U8301 ( .A(n11155), .B(n11178), .C(n11137), .D(n11203), .Y(n6640) );
  OAI21X1 U8303 ( .A(n11129), .B(n11236), .C(n6641), .Y(n6639) );
  AOI22X1 U8304 ( .A(n9188), .B(DATA_IN_H[4]), .C(n11163), .D(
        \U_0/U_0/U_0/extratemp[4] ), .Y(n6641) );
  NOR2X1 U8306 ( .A(n6642), .B(n6643), .Y(n6936) );
  OAI22X1 U8307 ( .A(n11155), .B(n11177), .C(n11137), .D(n11202), .Y(n6643) );
  OAI21X1 U8309 ( .A(n11129), .B(n11237), .C(n6644), .Y(n6642) );
  AOI22X1 U8310 ( .A(n9188), .B(DATA_IN_H[3]), .C(n11163), .D(
        \U_0/U_0/U_0/extratemp[3] ), .Y(n6644) );
  NOR2X1 U8312 ( .A(n6645), .B(n6646), .Y(n6935) );
  OAI22X1 U8313 ( .A(n11155), .B(n11176), .C(n11137), .D(n11201), .Y(n6646) );
  OAI21X1 U8314 ( .A(n11129), .B(n11238), .C(n6647), .Y(n6645) );
  AOI22X1 U8315 ( .A(n9188), .B(DATA_IN_H[2]), .C(n11163), .D(
        \U_0/U_0/U_0/extratemp[2] ), .Y(n6647) );
  NOR2X1 U8317 ( .A(n6648), .B(n6649), .Y(n6934) );
  OAI22X1 U8318 ( .A(n11155), .B(n11175), .C(n11137), .D(n11200), .Y(n6649) );
  OAI21X1 U8319 ( .A(n11129), .B(n11239), .C(n6650), .Y(n6648) );
  AOI22X1 U8320 ( .A(n9188), .B(DATA_IN_H[1]), .C(n11163), .D(
        \U_0/U_0/U_0/extratemp[1] ), .Y(n6650) );
  NOR2X1 U8322 ( .A(n6651), .B(n6652), .Y(n6933) );
  OAI22X1 U8323 ( .A(n11155), .B(n11174), .C(n11137), .D(n11199), .Y(n6652) );
  OAI21X1 U8326 ( .A(n11129), .B(n11240), .C(n6653), .Y(n6651) );
  AOI22X1 U8327 ( .A(n9188), .B(DATA_IN_H[0]), .C(n11163), .D(
        \U_0/U_0/U_0/extratemp[0] ), .Y(n6653) );
  NAND3X1 U8331 ( .A(n11130), .B(n562), .C(n6655), .Y(n6654) );
  NOR2X1 U8332 ( .A(n3673), .B(n6656), .Y(n6655) );
  NAND2X1 U8333 ( .A(n11149), .B(n3504), .Y(n6656) );
  NAND3X1 U8335 ( .A(n568), .B(n9166), .C(n3501), .Y(n6658) );
  NOR2X1 U8336 ( .A(n6660), .B(n3571), .Y(n568) );
  OAI21X1 U8337 ( .A(n6661), .B(n6662), .C(n6663), .Y(n3571) );
  OAI22X1 U8339 ( .A(n6662), .B(n6664), .C(n11161), .D(n6661), .Y(n6660) );
  NOR2X1 U8340 ( .A(n6666), .B(n6667), .Y(n6931) );
  NAND2X1 U8341 ( .A(n6668), .B(n6669), .Y(n6667) );
  AOI22X1 U8342 ( .A(\U_0/U_0/U_0/intj[7] ), .B(n6670), .C(\U_0/U_0/U_0/N448 ), 
        .D(n6671), .Y(n6669) );
  AOI22X1 U8343 ( .A(\U_0/U_0/U_0/inti[7] ), .B(n3674), .C(\U_0/U_0/U_0/N503 ), 
        .D(n6672), .Y(n6668) );
  NAND2X1 U8344 ( .A(n6673), .B(n6674), .Y(n6666) );
  AOI22X1 U8345 ( .A(\U_0/U_0/U_0/temp[7] ), .B(n9187), .C(\U_0/U_0/U_0/sj[7] ), .D(n6676), .Y(n6674) );
  AOI22X1 U8346 ( .A(\U_0/U_0/U_0/faddr [7]), .B(n6677), .C(
        \U_0/U_0/U_0/prefillCounter[7] ), .D(n3570), .Y(n6673) );
  NOR2X1 U8347 ( .A(n6678), .B(n6679), .Y(n6930) );
  NAND2X1 U8348 ( .A(n6680), .B(n6681), .Y(n6679) );
  AOI22X1 U8349 ( .A(\U_0/U_0/U_0/intj[6] ), .B(n6670), .C(\U_0/U_0/U_0/N447 ), 
        .D(n6671), .Y(n6681) );
  AOI22X1 U8350 ( .A(\U_0/U_0/U_0/inti[6] ), .B(n3674), .C(\U_0/U_0/U_0/N502 ), 
        .D(n6672), .Y(n6680) );
  NAND2X1 U8351 ( .A(n6682), .B(n6683), .Y(n6678) );
  AOI22X1 U8352 ( .A(\U_0/U_0/U_0/temp[6] ), .B(n9187), .C(\U_0/U_0/U_0/sj[6] ), .D(n6676), .Y(n6683) );
  AOI22X1 U8353 ( .A(\U_0/U_0/U_0/faddr [6]), .B(n6677), .C(
        \U_0/U_0/U_0/prefillCounter[6] ), .D(n3570), .Y(n6682) );
  NOR2X1 U8354 ( .A(n6684), .B(n6685), .Y(n6929) );
  NAND2X1 U8355 ( .A(n6686), .B(n6687), .Y(n6685) );
  AOI22X1 U8356 ( .A(\U_0/U_0/U_0/intj[5] ), .B(n6670), .C(\U_0/U_0/U_0/N446 ), 
        .D(n6671), .Y(n6687) );
  AOI22X1 U8357 ( .A(\U_0/U_0/U_0/inti[5] ), .B(n3674), .C(\U_0/U_0/U_0/N501 ), 
        .D(n6672), .Y(n6686) );
  NAND2X1 U8358 ( .A(n6688), .B(n6689), .Y(n6684) );
  AOI22X1 U8359 ( .A(\U_0/U_0/U_0/temp[5] ), .B(n9187), .C(\U_0/U_0/U_0/sj[5] ), .D(n6676), .Y(n6689) );
  AOI22X1 U8360 ( .A(\U_0/U_0/U_0/faddr [5]), .B(n6677), .C(
        \U_0/U_0/U_0/prefillCounter[5] ), .D(n3570), .Y(n6688) );
  NOR2X1 U8361 ( .A(n6690), .B(n6691), .Y(n6928) );
  NAND2X1 U8362 ( .A(n6692), .B(n6693), .Y(n6691) );
  AOI22X1 U8363 ( .A(\U_0/U_0/U_0/intj[4] ), .B(n6670), .C(\U_0/U_0/U_0/N445 ), 
        .D(n6671), .Y(n6693) );
  AOI22X1 U8364 ( .A(\U_0/U_0/U_0/inti[4] ), .B(n3674), .C(\U_0/U_0/U_0/N500 ), 
        .D(n6672), .Y(n6692) );
  NAND2X1 U8365 ( .A(n6694), .B(n6695), .Y(n6690) );
  AOI22X1 U8366 ( .A(\U_0/U_0/U_0/temp[4] ), .B(n9187), .C(\U_0/U_0/U_0/sj[4] ), .D(n6676), .Y(n6695) );
  AOI22X1 U8367 ( .A(\U_0/U_0/U_0/faddr [4]), .B(n6677), .C(
        \U_0/U_0/U_0/prefillCounter[4] ), .D(n3570), .Y(n6694) );
  NOR2X1 U8368 ( .A(n6696), .B(n6697), .Y(n6927) );
  NAND2X1 U8369 ( .A(n6698), .B(n6699), .Y(n6697) );
  AOI22X1 U8370 ( .A(\U_0/U_0/U_0/intj[3] ), .B(n6670), .C(\U_0/U_0/U_0/N444 ), 
        .D(n6671), .Y(n6699) );
  AOI22X1 U8371 ( .A(\U_0/U_0/U_0/inti[3] ), .B(n3674), .C(\U_0/U_0/U_0/N499 ), 
        .D(n6672), .Y(n6698) );
  NAND2X1 U8372 ( .A(n6700), .B(n6701), .Y(n6696) );
  AOI22X1 U8373 ( .A(\U_0/U_0/U_0/temp[3] ), .B(n9187), .C(\U_0/U_0/U_0/sj[3] ), .D(n6676), .Y(n6701) );
  AOI22X1 U8374 ( .A(\U_0/U_0/U_0/faddr [3]), .B(n6677), .C(
        \U_0/U_0/U_0/prefillCounter[3] ), .D(n3570), .Y(n6700) );
  NOR2X1 U8375 ( .A(n6702), .B(n6703), .Y(n6926) );
  NAND2X1 U8376 ( .A(n6704), .B(n6705), .Y(n6703) );
  AOI22X1 U8377 ( .A(\U_0/U_0/U_0/intj[2] ), .B(n6670), .C(\U_0/U_0/U_0/N443 ), 
        .D(n6671), .Y(n6705) );
  AOI22X1 U8378 ( .A(\U_0/U_0/U_0/inti[2] ), .B(n3674), .C(\U_0/U_0/U_0/N498 ), 
        .D(n6672), .Y(n6704) );
  NAND2X1 U8379 ( .A(n6706), .B(n6707), .Y(n6702) );
  AOI22X1 U8380 ( .A(\U_0/U_0/U_0/temp[2] ), .B(n9187), .C(\U_0/U_0/U_0/sj[2] ), .D(n6676), .Y(n6707) );
  AOI22X1 U8381 ( .A(\U_0/U_0/U_0/faddr [2]), .B(n6677), .C(
        \U_0/U_0/U_0/prefillCounter[2] ), .D(n3570), .Y(n6706) );
  NOR2X1 U8382 ( .A(n6708), .B(n6709), .Y(n6925) );
  NAND2X1 U8383 ( .A(n6710), .B(n6711), .Y(n6709) );
  AOI22X1 U8384 ( .A(\U_0/U_0/U_0/intj[1] ), .B(n6670), .C(\U_0/U_0/U_0/N442 ), 
        .D(n6671), .Y(n6711) );
  AOI22X1 U8385 ( .A(\U_0/U_0/U_0/inti[1] ), .B(n3674), .C(\U_0/U_0/U_0/N497 ), 
        .D(n6672), .Y(n6710) );
  NAND2X1 U8386 ( .A(n6712), .B(n6713), .Y(n6708) );
  AOI22X1 U8387 ( .A(\U_0/U_0/U_0/temp[1] ), .B(n9187), .C(\U_0/U_0/U_0/sj[1] ), .D(n6676), .Y(n6713) );
  AOI22X1 U8388 ( .A(\U_0/U_0/U_0/faddr [1]), .B(n6677), .C(
        \U_0/U_0/U_0/prefillCounter[1] ), .D(n3570), .Y(n6712) );
  NAND3X1 U8390 ( .A(n3501), .B(n11153), .C(n6714), .Y(n3444) );
  AOI21X1 U8391 ( .A(n6715), .B(n11167), .C(n6717), .Y(n6714) );
  NAND2X1 U8393 ( .A(n3558), .B(n3572), .Y(n3673) );
  NAND2X1 U8394 ( .A(n6718), .B(n3670), .Y(n3572) );
  NOR2X1 U8395 ( .A(n6719), .B(n11147), .Y(n3501) );
  NOR2X1 U8396 ( .A(n6721), .B(n6722), .Y(n6924) );
  NAND2X1 U8397 ( .A(n6723), .B(n6724), .Y(n6722) );
  AOI22X1 U8398 ( .A(\U_0/U_0/U_0/intj[0] ), .B(n6670), .C(n11242), .D(n6671), 
        .Y(n6724) );
  AOI22X1 U8399 ( .A(\U_0/U_0/U_0/inti[0] ), .B(n3674), .C(\U_0/U_0/U_0/N496 ), 
        .D(n6672), .Y(n6723) );
  OAI21X1 U8400 ( .A(n6725), .B(n11169), .C(n3583), .Y(n3674) );
  NAND2X1 U8401 ( .A(n3670), .B(n6727), .Y(n3583) );
  NAND2X1 U8402 ( .A(n6728), .B(n6729), .Y(n6721) );
  AOI22X1 U8403 ( .A(\U_0/U_0/U_0/temp[0] ), .B(n9187), .C(\U_0/U_0/U_0/sj[0] ), .D(n6676), .Y(n6729) );
  AOI22X1 U8404 ( .A(\U_0/U_0/U_0/faddr [0]), .B(n6677), .C(
        \U_0/U_0/U_0/prefillCounter[0] ), .D(n3570), .Y(n6728) );
  OAI21X1 U8405 ( .A(n11170), .B(n6731), .C(n562), .Y(n6677) );
  NOR2X1 U8406 ( .A(n3443), .B(n3438), .Y(n562) );
  NAND3X1 U8407 ( .A(n3503), .B(n6625), .C(n6732), .Y(n3443) );
  NAND2X1 U8408 ( .A(n11156), .B(n11171), .Y(n6731) );
  NAND2X1 U8409 ( .A(n6735), .B(n6736), .Y(\U_0/U_0/U_0/nextState [4]) );
  AOI22X1 U8410 ( .A(n10592), .B(n6737), .C(n10591), .D(n3655), .Y(n6736) );
  OAI21X1 U8411 ( .A(n11158), .B(n6739), .C(n6740), .Y(n6737) );
  OAI21X1 U8412 ( .A(n11092), .B(n11094), .C(n3476), .Y(n6740) );
  NAND2X1 U8413 ( .A(n6741), .B(n6742), .Y(n3476) );
  NAND2X1 U8414 ( .A(n6383), .B(\U_0/B_READY ), .Y(n6739) );
  AOI21X1 U8415 ( .A(n9320), .B(n11167), .C(n3477), .Y(n6735) );
  NAND3X1 U8416 ( .A(n569), .B(n6625), .C(n9189), .Y(n3477) );
  NAND3X1 U8418 ( .A(n6743), .B(n11142), .C(n6745), .Y(
        \U_0/U_0/U_0/nextState [3]) );
  NOR2X1 U8419 ( .A(n6746), .B(n6747), .Y(n6745) );
  OAI21X1 U8420 ( .A(n6732), .B(n6748), .C(n6749), .Y(n6747) );
  NAND3X1 U8421 ( .A(n11173), .B(n11171), .C(n6751), .Y(n6749) );
  NAND2X1 U8422 ( .A(n566), .B(n6625), .Y(n6746) );
  AOI22X1 U8423 ( .A(n6718), .B(n11166), .C(n6753), .D(
        \U_0/U_0/U_0/permuteComplete ), .Y(n6743) );
  NAND3X1 U8424 ( .A(n6754), .B(n11132), .C(n6756), .Y(
        \U_0/U_0/U_0/nextState [2]) );
  AOI21X1 U8425 ( .A(n10592), .B(n6757), .C(n6758), .Y(n6756) );
  OAI21X1 U8426 ( .A(\U_0/U_0/U_0/state[1] ), .B(n6661), .C(n11131), .Y(n6758)
         );
  OAI22X1 U8427 ( .A(n6759), .B(n6742), .C(n11157), .D(n6761), .Y(n6757) );
  AOI22X1 U8430 ( .A(n6718), .B(n6764), .C(n6753), .D(
        \U_0/U_0/U_0/permuteComplete ), .Y(n6754) );
  NAND3X1 U8431 ( .A(n6765), .B(n6766), .C(n6767), .Y(
        \U_0/U_0/U_0/nextState [1]) );
  NOR2X1 U8432 ( .A(n6768), .B(n6769), .Y(n6767) );
  OAI21X1 U8433 ( .A(n6770), .B(n6771), .C(n6772), .Y(n6769) );
  NAND3X1 U8434 ( .A(n10592), .B(n11165), .C(n6774), .Y(n6772) );
  OAI21X1 U8436 ( .A(n6775), .B(n6383), .C(\U_0/B_READY ), .Y(n6759) );
  NAND3X1 U8437 ( .A(n11175), .B(n11176), .C(n6776), .Y(n6771) );
  NOR2X1 U8438 ( .A(\U_0/U_0/U_0/prefillCounter[0] ), .B(n6941), .Y(n6776) );
  NAND3X1 U8441 ( .A(n6777), .B(n11179), .C(n6778), .Y(n6770) );
  NOR2X1 U8442 ( .A(\U_0/U_0/U_0/prefillCounter[4] ), .B(
        \U_0/U_0/U_0/prefillCounter[3] ), .Y(n6778) );
  NOR2X1 U8444 ( .A(\U_0/U_0/U_0/prefillCounter[7] ), .B(
        \U_0/U_0/U_0/prefillCounter[6] ), .Y(n6777) );
  AOI22X1 U8446 ( .A(n6727), .B(n6781), .C(n10591), .D(n6762), .Y(n6766) );
  OAI21X1 U8448 ( .A(n11164), .B(n6782), .C(n11170), .Y(n6781) );
  NAND2X1 U8449 ( .A(n6761), .B(n10592), .Y(n6782) );
  NOR2X1 U8450 ( .A(n6784), .B(n11092), .Y(n6761) );
  NOR2X1 U8452 ( .A(n6763), .B(n6785), .Y(n6765) );
  NAND3X1 U8454 ( .A(n11159), .B(n6788), .C(n6789), .Y(n6787) );
  NOR2X1 U8455 ( .A(n6719), .B(n6785), .Y(n6789) );
  OAI21X1 U8457 ( .A(\U_0/U_0/U_0/permuteComplete ), .B(n11150), .C(n11131), 
        .Y(n6790) );
  OAI21X1 U8458 ( .A(n6725), .B(n11169), .C(n566), .Y(n3569) );
  OAI21X1 U8459 ( .A(n11169), .B(n11162), .C(n3518), .Y(n6719) );
  OAI21X1 U8461 ( .A(n6793), .B(n6794), .C(n10592), .Y(n6788) );
  NAND3X1 U8463 ( .A(n6603), .B(n10600), .C(n10593), .Y(n6748) );
  NAND3X1 U8465 ( .A(n5682), .B(n10594), .C(n6797), .Y(n6795) );
  NOR2X1 U8466 ( .A(n10601), .B(n6799), .Y(n6797) );
  NAND2X1 U8467 ( .A(n5702), .B(n5684), .Y(n6799) );
  NAND3X1 U8468 ( .A(n6800), .B(n10605), .C(\U_0/U_0/U_1/U_8/state[0] ), .Y(
        n5684) );
  NAND3X1 U8471 ( .A(\U_0/U_0/U_1/U_8/state[2] ), .B(n10607), .C(n5731), .Y(
        n5685) );
  NAND2X1 U8473 ( .A(n5633), .B(n5698), .Y(n5663) );
  NAND3X1 U8474 ( .A(\U_0/U_0/U_1/U_8/state[0] ), .B(n6800), .C(
        \U_0/U_0/U_1/U_8/state[2] ), .Y(n5698) );
  NAND3X1 U8475 ( .A(n10597), .B(n10605), .C(n6800), .Y(n5633) );
  AOI21X1 U8476 ( .A(n10607), .B(n10599), .C(n10596), .Y(n5682) );
  NAND3X1 U8478 ( .A(n6800), .B(n10597), .C(\U_0/U_0/U_1/U_8/state[2] ), .Y(
        n5701) );
  NOR2X1 U8480 ( .A(n10608), .B(\U_0/U_0/U_1/U_8/state[3] ), .Y(n6800) );
  NOR2X1 U8483 ( .A(n10607), .B(n5732), .Y(n5724) );
  NAND2X1 U8484 ( .A(n5731), .B(n10605), .Y(n5732) );
  NOR2X1 U8485 ( .A(\U_0/U_0/U_1/U_8/state[1] ), .B(\U_0/U_0/U_1/U_8/state[0] ), .Y(n5731) );
  NAND2X1 U8486 ( .A(\U_0/U_0/U_1/U_8/parityError ), .B(n5723), .Y(n6603) );
  NOR2X1 U8487 ( .A(n6801), .B(n10605), .Y(n5723) );
  NAND3X1 U8489 ( .A(n10608), .B(n10607), .C(\U_0/U_0/U_1/U_8/state[0] ), .Y(
        n6801) );
  OAI22X1 U8492 ( .A(\U_0/U_0/U_0/state[3] ), .B(n11161), .C(\U_0/B_READY ), 
        .D(n6742), .Y(n6794) );
  OAI21X1 U8493 ( .A(n11094), .B(n6803), .C(n6804), .Y(n6793) );
  NAND3X1 U8494 ( .A(n6784), .B(n11093), .C(n11152), .Y(n6804) );
  NOR2X1 U8496 ( .A(n11095), .B(n11113), .Y(n6383) );
  NAND2X1 U8497 ( .A(n11113), .B(n11095), .Y(n6784) );
  NAND2X1 U8499 ( .A(\U_0/B_READY ), .B(n6762), .Y(n6803) );
  NOR2X1 U8501 ( .A(n11095), .B(\U_0/PRGA_OPCODE[1] ), .Y(n6775) );
  NAND3X1 U8503 ( .A(n569), .B(n6625), .C(n6806), .Y(n6786) );
  NOR2X1 U8505 ( .A(n9191), .B(n6779), .Y(n6625) );
  OAI21X1 U8506 ( .A(n6808), .B(n11206), .C(n6810), .Y(
        \U_0/U_0/U_0/nextProcessedData[7] ) );
  AOI22X1 U8507 ( .A(n9191), .B(n6811), .C(\U_0/PRGA_IN [7]), .D(n6779), .Y(
        n6810) );
  XNOR2X1 U8508 ( .A(n11205), .B(\U_0/U_0/U_0/delaydata [7]), .Y(n6811) );
  OAI21X1 U8511 ( .A(n6808), .B(n11208), .C(n6813), .Y(
        \U_0/U_0/U_0/nextProcessedData[6] ) );
  AOI22X1 U8512 ( .A(n9191), .B(n6814), .C(\U_0/PRGA_IN [6]), .D(n6779), .Y(
        n6813) );
  XNOR2X1 U8513 ( .A(n11198), .B(\U_0/U_0/U_0/delaydata [6]), .Y(n6814) );
  OAI21X1 U8516 ( .A(n6808), .B(n11211), .C(n6816), .Y(
        \U_0/U_0/U_0/nextProcessedData[5] ) );
  AOI22X1 U8517 ( .A(n9191), .B(n6817), .C(\U_0/PRGA_IN [5]), .D(n6779), .Y(
        n6816) );
  XNOR2X1 U8518 ( .A(n11204), .B(\U_0/U_0/U_0/delaydata [5]), .Y(n6817) );
  OAI21X1 U8521 ( .A(n6808), .B(n11212), .C(n6819), .Y(
        \U_0/U_0/U_0/nextProcessedData[4] ) );
  AOI22X1 U8522 ( .A(n9191), .B(n6820), .C(\U_0/PRGA_IN [4]), .D(n6779), .Y(
        n6819) );
  XNOR2X1 U8523 ( .A(n11203), .B(\U_0/U_0/U_0/delaydata [4]), .Y(n6820) );
  OAI21X1 U8526 ( .A(n6808), .B(n11214), .C(n6822), .Y(
        \U_0/U_0/U_0/nextProcessedData[3] ) );
  AOI22X1 U8527 ( .A(n9191), .B(n6823), .C(\U_0/PRGA_IN [3]), .D(n6779), .Y(
        n6822) );
  XNOR2X1 U8528 ( .A(n11202), .B(\U_0/U_0/U_0/delaydata [3]), .Y(n6823) );
  OAI21X1 U8531 ( .A(n6808), .B(n11215), .C(n6825), .Y(
        \U_0/U_0/U_0/nextProcessedData[2] ) );
  AOI22X1 U8532 ( .A(n9191), .B(n6826), .C(\U_0/PRGA_IN [2]), .D(n6779), .Y(
        n6825) );
  XNOR2X1 U8533 ( .A(n11201), .B(\U_0/U_0/U_0/delaydata [2]), .Y(n6826) );
  OAI21X1 U8536 ( .A(n6808), .B(n11216), .C(n6828), .Y(
        \U_0/U_0/U_0/nextProcessedData[1] ) );
  AOI22X1 U8537 ( .A(n9191), .B(n6829), .C(\U_0/PRGA_IN [1]), .D(n6779), .Y(
        n6828) );
  XNOR2X1 U8538 ( .A(n11200), .B(\U_0/U_0/U_0/delaydata [1]), .Y(n6829) );
  OAI21X1 U8541 ( .A(n6808), .B(n11217), .C(n6831), .Y(
        \U_0/U_0/U_0/nextProcessedData[0] ) );
  AOI22X1 U8542 ( .A(n9191), .B(n6832), .C(\U_0/PRGA_IN [0]), .D(n6779), .Y(
        n6831) );
  NOR2X1 U8543 ( .A(n6833), .B(n6725), .Y(n6779) );
  XNOR2X1 U8544 ( .A(n11199), .B(\U_0/U_0/U_0/delaydata [0]), .Y(n6832) );
  NOR2X1 U8546 ( .A(n6833), .B(n11162), .Y(n6807) );
  NOR2X1 U8548 ( .A(n6834), .B(n6835), .Y(n6808) );
  NAND3X1 U8549 ( .A(n3667), .B(n6732), .C(n6836), .Y(n6835) );
  NOR2X1 U8550 ( .A(n6670), .B(n6763), .Y(n6836) );
  NAND3X1 U8551 ( .A(n569), .B(n3558), .C(n11142), .Y(n6763) );
  NAND2X1 U8553 ( .A(n3518), .B(n9190), .Y(n3585) );
  NOR2X1 U8555 ( .A(n6664), .B(n6837), .Y(n6672) );
  NAND2X1 U8556 ( .A(n6715), .B(n11168), .Y(n3518) );
  NAND3X1 U8557 ( .A(n9320), .B(n11166), .C(n6727), .Y(n3558) );
  NAND2X1 U8558 ( .A(n9320), .B(n9187), .Y(n569) );
  OAI21X1 U8559 ( .A(n6664), .B(n6662), .C(n567), .Y(n6670) );
  NAND3X1 U8560 ( .A(n9320), .B(n11166), .C(n3669), .Y(n567) );
  NOR2X1 U8561 ( .A(n6762), .B(n11152), .Y(n6732) );
  OAI21X1 U8563 ( .A(n6718), .B(n6727), .C(n11165), .Y(n6742) );
  NAND2X1 U8565 ( .A(n6751), .B(n9320), .Y(n6833) );
  NAND2X1 U8566 ( .A(n11158), .B(n6741), .Y(n6762) );
  NAND3X1 U8567 ( .A(n11168), .B(n9320), .C(n3669), .Y(n6741) );
  NOR2X1 U8570 ( .A(n11161), .B(n6664), .Y(n3655) );
  NAND2X1 U8571 ( .A(\U_0/U_0/U_0/state[3] ), .B(\U_0/U_0/U_0/state[2] ), .Y(
        n6664) );
  NOR2X1 U8572 ( .A(n6839), .B(n6840), .Y(n3667) );
  NAND3X1 U8573 ( .A(n11136), .B(n11141), .C(n11159), .Y(n6840) );
  OAI21X1 U8575 ( .A(n6661), .B(n11161), .C(n11160), .Y(n6671) );
  NOR2X1 U8577 ( .A(n11164), .B(n11161), .Y(n6631) );
  NAND2X1 U8580 ( .A(n11149), .B(n6941), .Y(n3563) );
  NAND2X1 U8581 ( .A(n6715), .B(n6764), .Y(n6941) );
  OAI21X1 U8583 ( .A(n6837), .B(n11164), .C(n11150), .Y(n6717) );
  NOR2X1 U8585 ( .A(n11164), .B(n6662), .Y(n6753) );
  OAI21X1 U8588 ( .A(n6661), .B(n6662), .C(n566), .Y(n6676) );
  NAND2X1 U8589 ( .A(n6751), .B(n6715), .Y(n566) );
  NOR2X1 U8590 ( .A(n6725), .B(n9320), .Y(n6715) );
  NOR2X1 U8591 ( .A(n11167), .B(\U_0/U_0/U_0/state[2] ), .Y(n6751) );
  NAND3X1 U8592 ( .A(n3503), .B(n11131), .C(n11148), .Y(n6839) );
  NOR2X1 U8594 ( .A(n6662), .B(n11170), .Y(n3438) );
  NAND2X1 U8595 ( .A(n6718), .B(n11171), .Y(n6662) );
  NOR2X1 U8597 ( .A(n9166), .B(n9320), .Y(n3481) );
  NAND2X1 U8600 ( .A(\U_0/U_0/U_0/state[1] ), .B(n11156), .Y(n6725) );
  NAND2X1 U8601 ( .A(n11154), .B(n11166), .Y(n3503) );
  NAND3X1 U8603 ( .A(n11155), .B(n3504), .C(n6843), .Y(n6834) );
  NOR2X1 U8604 ( .A(n3670), .B(n11147), .Y(n6843) );
  NAND3X1 U8606 ( .A(n9320), .B(n11166), .C(n6718), .Y(n3672) );
  NOR2X1 U8607 ( .A(n11156), .B(n11173), .Y(n6718) );
  NAND2X1 U8610 ( .A(\U_0/U_0/U_0/state[2] ), .B(n11167), .Y(n6661) );
  NOR2X1 U8612 ( .A(n11170), .B(n11171), .Y(n3670) );
  NAND2X1 U8613 ( .A(n6842), .B(n6764), .Y(n3504) );
  NOR2X1 U8614 ( .A(n11162), .B(n9320), .Y(n6842) );
  NOR2X1 U8616 ( .A(\U_0/U_0/U_0/state[0] ), .B(\U_0/U_0/U_0/state[1] ), .Y(
        n3669) );
  NOR2X1 U8618 ( .A(n11170), .B(n6837), .Y(n3570) );
  NAND2X1 U8619 ( .A(n6727), .B(n11171), .Y(n6837) );
  NOR2X1 U8621 ( .A(n11156), .B(\U_0/U_0/U_0/state[1] ), .Y(n6727) );
  NOR2X1 U8624 ( .A(\U_0/U_0/U_0/state[2] ), .B(\U_0/U_0/U_0/state[3] ), .Y(
        n6764) );
  NAND3X1 U8625 ( .A(n6844), .B(n6845), .C(n6846), .Y(\U_0/U_0/U_0/N479 ) );
  NOR2X1 U8626 ( .A(n6847), .B(n6848), .Y(n6846) );
  OAI22X1 U8627 ( .A(n11280), .B(n6850), .C(n11261), .D(n6851), .Y(n6848) );
  OAI22X1 U8630 ( .A(n11264), .B(n6853), .C(n11272), .D(n6855), .Y(n6847) );
  AOI22X1 U8633 ( .A(n11244), .B(\U_0/U_0/U_0/keyTable[5][0] ), .C(n11243), 
        .D(\U_0/U_0/U_0/keyTable[4][0] ), .Y(n6845) );
  AOI22X1 U8634 ( .A(n11247), .B(\U_0/U_0/U_0/keyTable[7][0] ), .C(n11246), 
        .D(\U_0/U_0/U_0/keyTable[6][0] ), .Y(n6844) );
  NAND3X1 U8635 ( .A(n6860), .B(n6861), .C(n6862), .Y(\U_0/U_0/U_0/N478 ) );
  NOR2X1 U8636 ( .A(n6863), .B(n6864), .Y(n6862) );
  OAI22X1 U8637 ( .A(n11281), .B(n6850), .C(n11260), .D(n6851), .Y(n6864) );
  OAI22X1 U8640 ( .A(n11265), .B(n6853), .C(n11273), .D(n6855), .Y(n6863) );
  AOI22X1 U8643 ( .A(n11244), .B(\U_0/U_0/U_0/keyTable[5][1] ), .C(n11243), 
        .D(\U_0/U_0/U_0/keyTable[4][1] ), .Y(n6861) );
  AOI22X1 U8644 ( .A(n11247), .B(\U_0/U_0/U_0/keyTable[7][1] ), .C(n11246), 
        .D(\U_0/U_0/U_0/keyTable[6][1] ), .Y(n6860) );
  NAND3X1 U8645 ( .A(n6868), .B(n6869), .C(n6870), .Y(\U_0/U_0/U_0/N477 ) );
  NOR2X1 U8646 ( .A(n6871), .B(n6872), .Y(n6870) );
  OAI22X1 U8647 ( .A(n11282), .B(n6850), .C(n11259), .D(n6851), .Y(n6872) );
  OAI22X1 U8650 ( .A(n11266), .B(n6853), .C(n11274), .D(n6855), .Y(n6871) );
  AOI22X1 U8653 ( .A(n11244), .B(\U_0/U_0/U_0/keyTable[5][2] ), .C(n11243), 
        .D(\U_0/U_0/U_0/keyTable[4][2] ), .Y(n6869) );
  AOI22X1 U8654 ( .A(n11247), .B(\U_0/U_0/U_0/keyTable[7][2] ), .C(n11246), 
        .D(\U_0/U_0/U_0/keyTable[6][2] ), .Y(n6868) );
  NAND3X1 U8655 ( .A(n6876), .B(n6877), .C(n6878), .Y(\U_0/U_0/U_0/N476 ) );
  NOR2X1 U8656 ( .A(n6879), .B(n6880), .Y(n6878) );
  OAI22X1 U8657 ( .A(n11283), .B(n6850), .C(n11258), .D(n6851), .Y(n6880) );
  OAI22X1 U8660 ( .A(n11267), .B(n6853), .C(n11275), .D(n6855), .Y(n6879) );
  AOI22X1 U8663 ( .A(n11244), .B(\U_0/U_0/U_0/keyTable[5][3] ), .C(n11243), 
        .D(\U_0/U_0/U_0/keyTable[4][3] ), .Y(n6877) );
  AOI22X1 U8664 ( .A(n11247), .B(\U_0/U_0/U_0/keyTable[7][3] ), .C(n11246), 
        .D(\U_0/U_0/U_0/keyTable[6][3] ), .Y(n6876) );
  NAND3X1 U8665 ( .A(n6884), .B(n6885), .C(n6886), .Y(\U_0/U_0/U_0/N475 ) );
  NOR2X1 U8666 ( .A(n6887), .B(n6888), .Y(n6886) );
  OAI22X1 U8667 ( .A(n11284), .B(n6850), .C(n11257), .D(n6851), .Y(n6888) );
  OAI22X1 U8670 ( .A(n11268), .B(n6853), .C(n11276), .D(n6855), .Y(n6887) );
  AOI22X1 U8673 ( .A(n11244), .B(\U_0/U_0/U_0/keyTable[5][4] ), .C(n11243), 
        .D(\U_0/U_0/U_0/keyTable[4][4] ), .Y(n6885) );
  AOI22X1 U8674 ( .A(n11247), .B(\U_0/U_0/U_0/keyTable[7][4] ), .C(n11246), 
        .D(\U_0/U_0/U_0/keyTable[6][4] ), .Y(n6884) );
  NAND3X1 U8675 ( .A(n6893), .B(n6894), .C(n6895), .Y(\U_0/U_0/U_0/N474 ) );
  NOR2X1 U8676 ( .A(n6896), .B(n6897), .Y(n6895) );
  OAI22X1 U8677 ( .A(n11285), .B(n6850), .C(n11256), .D(n6851), .Y(n6897) );
  OAI22X1 U8680 ( .A(n11269), .B(n6853), .C(n11277), .D(n6855), .Y(n6896) );
  AOI22X1 U8683 ( .A(n11244), .B(\U_0/U_0/U_0/keyTable[5][5] ), .C(n11243), 
        .D(\U_0/U_0/U_0/keyTable[4][5] ), .Y(n6894) );
  AOI22X1 U8684 ( .A(n11247), .B(\U_0/U_0/U_0/keyTable[7][5] ), .C(n11246), 
        .D(\U_0/U_0/U_0/keyTable[6][5] ), .Y(n6893) );
  NAND3X1 U8685 ( .A(n6902), .B(n6903), .C(n6904), .Y(\U_0/U_0/U_0/N473 ) );
  NOR2X1 U8686 ( .A(n6905), .B(n6906), .Y(n6904) );
  OAI22X1 U8687 ( .A(n11286), .B(n6850), .C(n11255), .D(n6851), .Y(n6906) );
  OAI22X1 U8690 ( .A(n11270), .B(n6853), .C(n11278), .D(n6855), .Y(n6905) );
  AOI22X1 U8693 ( .A(n11244), .B(\U_0/U_0/U_0/keyTable[5][6] ), .C(n11243), 
        .D(\U_0/U_0/U_0/keyTable[4][6] ), .Y(n6903) );
  AOI22X1 U8694 ( .A(n11247), .B(\U_0/U_0/U_0/keyTable[7][6] ), .C(n11246), 
        .D(\U_0/U_0/U_0/keyTable[6][6] ), .Y(n6902) );
  NAND3X1 U8695 ( .A(n6911), .B(n6912), .C(n6913), .Y(\U_0/U_0/U_0/N472 ) );
  NOR2X1 U8696 ( .A(n6914), .B(n6915), .Y(n6913) );
  OAI22X1 U8697 ( .A(n11262), .B(n6850), .C(n11263), .D(n6851), .Y(n6915) );
  NAND3X1 U8698 ( .A(n11245), .B(n11249), .C(n11253), .Y(n6851) );
  NAND3X1 U8700 ( .A(n11245), .B(n11249), .C(\U_0/U_0/U_0/keyi[0] ), .Y(n6850)
         );
  OAI22X1 U8702 ( .A(n11271), .B(n6853), .C(n11279), .D(n6855), .Y(n6914) );
  NAND3X1 U8703 ( .A(n11253), .B(n11249), .C(\U_0/U_0/U_0/keyi[1] ), .Y(n6855)
         );
  NAND3X1 U8705 ( .A(\U_0/U_0/U_0/keyi[1] ), .B(n11249), .C(
        \U_0/U_0/U_0/keyi[0] ), .Y(n6853) );
  AOI22X1 U8708 ( .A(n11244), .B(\U_0/U_0/U_0/keyTable[5][7] ), .C(n11243), 
        .D(\U_0/U_0/U_0/keyTable[4][7] ), .Y(n6912) );
  NAND3X1 U8710 ( .A(n11253), .B(n11245), .C(\U_0/U_0/U_0/keyi[2] ), .Y(n6920)
         );
  NAND3X1 U8712 ( .A(\U_0/U_0/U_0/keyi[2] ), .B(n11245), .C(
        \U_0/U_0/U_0/keyi[0] ), .Y(n6921) );
  AOI22X1 U8714 ( .A(n11247), .B(\U_0/U_0/U_0/keyTable[7][7] ), .C(n11246), 
        .D(\U_0/U_0/U_0/keyTable[6][7] ), .Y(n6911) );
  NAND3X1 U8716 ( .A(\U_0/U_0/U_0/keyi[2] ), .B(n11253), .C(
        \U_0/U_0/U_0/keyi[1] ), .Y(n6922) );
  NAND3X1 U8719 ( .A(\U_0/U_0/U_0/keyi[1] ), .B(\U_0/U_0/U_0/keyi[2] ), .C(
        \U_0/U_0/U_0/keyi[0] ), .Y(n6923) );
  AND2X2 U14 ( .A(n196), .B(n197), .Y(n194) );
  AND2X2 U21 ( .A(n204), .B(n205), .Y(n202) );
  AND2X2 U28 ( .A(n209), .B(n210), .Y(n207) );
  AND2X2 U35 ( .A(n214), .B(n215), .Y(n212) );
  AND2X2 U42 ( .A(n219), .B(n220), .Y(n217) );
  AND2X2 U51 ( .A(n224), .B(n225), .Y(n222) );
  AND2X2 U97 ( .A(n228), .B(n9501), .Y(n179) );
  AND2X2 U99 ( .A(n230), .B(n231), .Y(n227) );
  AND2X2 U222 ( .A(n318), .B(n11898), .Y(n317) );
  AND2X2 U223 ( .A(n9179), .B(n320), .Y(n315) );
  AND2X2 U274 ( .A(n362), .B(n9507), .Y(n326) );
  OR2X2 U423 ( .A(\U_1/U_0/U_1/SET_RBUF_FULL ), .B(\U_1/RBUF_FULL ), .Y(n7299)
         );
  AND2X2 U437 ( .A(n482), .B(n483), .Y(n480) );
  AND2X2 U444 ( .A(n490), .B(n491), .Y(n488) );
  AND2X2 U451 ( .A(n495), .B(n496), .Y(n493) );
  AND2X2 U458 ( .A(n500), .B(n501), .Y(n498) );
  AND2X2 U465 ( .A(n505), .B(n506), .Y(n503) );
  AND2X2 U472 ( .A(n510), .B(n511), .Y(n508) );
  AND2X2 U478 ( .A(n514), .B(n9506), .Y(n465) );
  AND2X2 U480 ( .A(n516), .B(n517), .Y(n513) );
  OR2X2 U541 ( .A(n560), .B(n561), .Y(n556) );
  AND2X2 U646 ( .A(n646), .B(n9505), .Y(n610) );
  OR2X2 U795 ( .A(\U_0/U_0/U_1/SET_RBUF_FULL ), .B(\U_0/RBUF_FULL ), .Y(n7691)
         );
  AND2X2 U939 ( .A(n191), .B(n11650), .Y(n875) );
  AND2X2 U975 ( .A(n9197), .B(n9276), .Y(n896) );
  OR2X2 U978 ( .A(n917), .B(n918), .Y(n916) );
  AND2X2 U1072 ( .A(n316), .B(n10520), .Y(n1009) );
  AND2X2 U1079 ( .A(n11913), .B(n1020), .Y(n1019) );
  AND2X2 U1099 ( .A(n321), .B(n1033), .Y(n1017) );
  AND2X2 U1170 ( .A(n11895), .B(n9277), .Y(n1068) );
  AND2X2 U1181 ( .A(n1098), .B(n1099), .Y(n1092) );
  OR2X2 U1320 ( .A(n1176), .B(n1177), .Y(n1175) );
  OR2X2 U1333 ( .A(n1212), .B(n1213), .Y(n1174) );
  OR2X2 U1349 ( .A(n1251), .B(n1252), .Y(n1250) );
  OR2X2 U1362 ( .A(n1271), .B(n1272), .Y(n1249) );
  OR2X2 U1378 ( .A(n1294), .B(n1295), .Y(n1293) );
  OR2X2 U1391 ( .A(n1314), .B(n1315), .Y(n1292) );
  OR2X2 U1407 ( .A(n1337), .B(n1338), .Y(n1336) );
  OR2X2 U1420 ( .A(n1357), .B(n1358), .Y(n1335) );
  OR2X2 U1436 ( .A(n1380), .B(n1381), .Y(n1379) );
  OR2X2 U1449 ( .A(n1400), .B(n1401), .Y(n1378) );
  OR2X2 U1465 ( .A(n1423), .B(n1424), .Y(n1422) );
  OR2X2 U1478 ( .A(n1443), .B(n1444), .Y(n1421) );
  OR2X2 U1494 ( .A(n1466), .B(n1467), .Y(n1465) );
  OR2X2 U1507 ( .A(n1486), .B(n1487), .Y(n1464) );
  OR2X2 U1523 ( .A(n1509), .B(n1510), .Y(n1508) );
  OR2X2 U1536 ( .A(n1529), .B(n1530), .Y(n1507) );
  OR2X2 U1552 ( .A(n1552), .B(n1553), .Y(n1551) );
  OR2X2 U1565 ( .A(n1572), .B(n1573), .Y(n1550) );
  OR2X2 U1581 ( .A(n1595), .B(n1596), .Y(n1594) );
  AND2X2 U1591 ( .A(n11665), .B(n1610), .Y(n1192) );
  AND2X2 U1592 ( .A(n11661), .B(n1610), .Y(n1191) );
  AND2X2 U1594 ( .A(n11665), .B(n1611), .Y(n1194) );
  AND2X2 U1597 ( .A(n11661), .B(n1611), .Y(n1193) );
  AND2X2 U1609 ( .A(n11666), .B(n1605), .Y(n1209) );
  AND2X2 U1610 ( .A(n11662), .B(n1605), .Y(n1208) );
  AND2X2 U1612 ( .A(n11666), .B(n1609), .Y(n1211) );
  AND2X2 U1615 ( .A(n11662), .B(n1609), .Y(n1210) );
  OR2X2 U1618 ( .A(n1629), .B(n1630), .Y(n1593) );
  AND2X2 U1628 ( .A(n11667), .B(n1605), .Y(n1228) );
  AND2X2 U1629 ( .A(n11663), .B(n1605), .Y(n1227) );
  AND2X2 U1631 ( .A(n11667), .B(n1609), .Y(n1230) );
  AND2X2 U1634 ( .A(n11663), .B(n1609), .Y(n1229) );
  AND2X2 U1642 ( .A(\U_1/U_1/U_1/readptr[2] ), .B(n9299), .Y(n1609) );
  AND2X2 U1646 ( .A(\U_1/U_1/U_1/readptr[2] ), .B(\U_1/U_1/U_1/readptr[1] ), 
        .Y(n1605) );
  AND2X2 U1648 ( .A(n11664), .B(n1611), .Y(n1245) );
  AND2X2 U1649 ( .A(n1611), .B(n11668), .Y(n1244) );
  AND2X2 U1652 ( .A(n1610), .B(n11664), .Y(n1247) );
  AND2X2 U1656 ( .A(n1610), .B(n11668), .Y(n1246) );
  AND2X2 U2451 ( .A(n1987), .B(n9504), .Y(n1902) );
  AND2X2 U2453 ( .A(n1988), .B(n9508), .Y(n1923) );
  AND2X2 U2476 ( .A(n879), .B(n1997), .Y(n882) );
  AND2X2 U2834 ( .A(n9445), .B(n2330), .Y(n2329) );
  AND2X2 U2849 ( .A(n9445), .B(n2346), .Y(n2345) );
  AND2X2 U2864 ( .A(n9446), .B(n2361), .Y(n2360) );
  AND2X2 U2879 ( .A(n9446), .B(n2376), .Y(n2375) );
  AND2X2 U2894 ( .A(n9446), .B(n2391), .Y(n2390) );
  AND2X2 U2909 ( .A(n9446), .B(n2406), .Y(n2405) );
  AND2X2 U2924 ( .A(n9446), .B(n2421), .Y(n2420) );
  AND2X2 U2933 ( .A(n2193), .B(n11508), .Y(n2320) );
  AND2X2 U2934 ( .A(n2429), .B(n2319), .Y(n2193) );
  AND2X2 U2941 ( .A(n9446), .B(n2438), .Y(n2437) );
  AND2X2 U2948 ( .A(n2319), .B(n11508), .Y(n2336) );
  AND2X2 U2957 ( .A(n9446), .B(n2454), .Y(n2453) );
  AND2X2 U2972 ( .A(n9446), .B(n2469), .Y(n2468) );
  AND2X2 U2987 ( .A(n9445), .B(n2483), .Y(n2482) );
  AND2X2 U3002 ( .A(n9445), .B(n2497), .Y(n2496) );
  AND2X2 U3017 ( .A(n9445), .B(n2511), .Y(n2510) );
  AND2X2 U3032 ( .A(n9445), .B(n2525), .Y(n2524) );
  AND2X2 U3047 ( .A(n9445), .B(n2539), .Y(n2538) );
  AND2X2 U3062 ( .A(n9445), .B(n2553), .Y(n2552) );
  AND2X2 U3069 ( .A(n2559), .B(\U_1/U_0/U_1/U_8/address[3] ), .Y(n2460) );
  AND2X2 U3078 ( .A(n9445), .B(n2569), .Y(n2568) );
  AND2X2 U3093 ( .A(n9445), .B(n2584), .Y(n2583) );
  AND2X2 U3108 ( .A(n9445), .B(n2598), .Y(n2597) );
  AND2X2 U3123 ( .A(n9445), .B(n2612), .Y(n2611) );
  AND2X2 U3138 ( .A(n9445), .B(n2626), .Y(n2625) );
  AND2X2 U3153 ( .A(n9445), .B(n2640), .Y(n2639) );
  AND2X2 U3168 ( .A(n9445), .B(n2654), .Y(n2653) );
  AND2X2 U3177 ( .A(n2444), .B(n11508), .Y(n2560) );
  AND2X2 U3178 ( .A(n2559), .B(n2429), .Y(n2444) );
  AND2X2 U3185 ( .A(n9445), .B(n2668), .Y(n2667) );
  AND2X2 U3192 ( .A(n2559), .B(n11508), .Y(n2575) );
  AND2X2 U3202 ( .A(n9445), .B(n2684), .Y(n2683) );
  AND2X2 U3217 ( .A(n9445), .B(n2699), .Y(n2698) );
  AND2X2 U3232 ( .A(n9445), .B(n2713), .Y(n2712) );
  AND2X2 U3247 ( .A(n9445), .B(n2727), .Y(n2726) );
  AND2X2 U3262 ( .A(n9445), .B(n2741), .Y(n2740) );
  AND2X2 U3277 ( .A(n9445), .B(n2755), .Y(n2754) );
  AND2X2 U3292 ( .A(n9445), .B(n2769), .Y(n2768) );
  AND2X2 U3307 ( .A(n9445), .B(n2783), .Y(n2782) );
  AND2X2 U3314 ( .A(n2789), .B(\U_1/U_0/U_1/U_8/address[3] ), .Y(n2690) );
  AND2X2 U3323 ( .A(n9445), .B(n2799), .Y(n2798) );
  AND2X2 U3338 ( .A(n9445), .B(n2814), .Y(n2813) );
  AND2X2 U3353 ( .A(n9445), .B(n2828), .Y(n2827) );
  AND2X2 U3368 ( .A(n9445), .B(n2842), .Y(n2841) );
  AND2X2 U3383 ( .A(n9445), .B(n2856), .Y(n2855) );
  AND2X2 U3398 ( .A(n9445), .B(n2870), .Y(n2869) );
  AND2X2 U3413 ( .A(n9445), .B(n2884), .Y(n2883) );
  AND2X2 U3422 ( .A(n2675), .B(n11508), .Y(n2790) );
  AND2X2 U3423 ( .A(n2789), .B(n2429), .Y(n2675) );
  AND2X2 U3430 ( .A(n9445), .B(n2898), .Y(n2897) );
  AND2X2 U3437 ( .A(n2789), .B(n11508), .Y(n2805) );
  AND2X2 U3447 ( .A(n9445), .B(n2914), .Y(n2913) );
  AND2X2 U3462 ( .A(n9445), .B(n2929), .Y(n2928) );
  AND2X2 U3477 ( .A(n9445), .B(n2943), .Y(n2942) );
  AND2X2 U3492 ( .A(n9445), .B(n2957), .Y(n2956) );
  AND2X2 U3507 ( .A(n9445), .B(n2971), .Y(n2970) );
  AND2X2 U3522 ( .A(n9446), .B(n2985), .Y(n2984) );
  AND2X2 U3537 ( .A(n9445), .B(n2999), .Y(n2998) );
  AND2X2 U3553 ( .A(n9445), .B(n3013), .Y(n3012) );
  AND2X2 U3560 ( .A(n3019), .B(\U_1/U_0/U_1/U_8/address[3] ), .Y(n2920) );
  AND2X2 U3569 ( .A(n2177), .B(n3029), .Y(n3028) );
  AND2X2 U3585 ( .A(n2177), .B(n3044), .Y(n3043) );
  AND2X2 U3601 ( .A(n2177), .B(n3059), .Y(n3058) );
  AND2X2 U3617 ( .A(n2177), .B(n3073), .Y(n3072) );
  AND2X2 U3685 ( .A(n2905), .B(n11508), .Y(n3020) );
  AND2X2 U3686 ( .A(n3019), .B(n2429), .Y(n2905) );
  AND2X2 U3718 ( .A(n3019), .B(n11508), .Y(n3035) );
  AND2X2 U3772 ( .A(n9245), .B(n3162), .Y(n3147) );
  AND2X2 U3829 ( .A(n9245), .B(n3197), .Y(n3142) );
  OR2X2 U3850 ( .A(n3224), .B(n3225), .Y(n8442) );
  AND2X2 U3879 ( .A(n3236), .B(n11320), .Y(n3251) );
  OR2X2 U3903 ( .A(\U_1/U_0/U_1/U_7/state[5] ), .B(\U_1/U_0/U_1/U_7/state[6] ), 
        .Y(n3270) );
  AND2X2 U3932 ( .A(n3279), .B(n3296), .Y(n3281) );
  OR2X2 U3935 ( .A(n3297), .B(n3298), .Y(n3296) );
  AND2X2 U4240 ( .A(n9515), .B(n569), .Y(n3565) );
  AND2X2 U4245 ( .A(n3504), .B(n3572), .Y(n3561) );
  OR2X2 U4427 ( .A(n3679), .B(n3680), .Y(n3678) );
  OR2X2 U4440 ( .A(n3715), .B(n3716), .Y(n3677) );
  OR2X2 U4456 ( .A(n3754), .B(n3755), .Y(n3753) );
  OR2X2 U4469 ( .A(n3774), .B(n3775), .Y(n3752) );
  OR2X2 U4485 ( .A(n3797), .B(n3798), .Y(n3796) );
  OR2X2 U4498 ( .A(n3817), .B(n3818), .Y(n3795) );
  OR2X2 U4514 ( .A(n3840), .B(n3841), .Y(n3839) );
  OR2X2 U4527 ( .A(n3860), .B(n3861), .Y(n3838) );
  OR2X2 U4543 ( .A(n3883), .B(n3884), .Y(n3882) );
  OR2X2 U4556 ( .A(n3903), .B(n3904), .Y(n3881) );
  OR2X2 U4572 ( .A(n3926), .B(n3927), .Y(n3925) );
  OR2X2 U4585 ( .A(n3946), .B(n3947), .Y(n3924) );
  OR2X2 U4601 ( .A(n3969), .B(n3970), .Y(n3968) );
  OR2X2 U4614 ( .A(n3989), .B(n3990), .Y(n3967) );
  OR2X2 U4630 ( .A(n4012), .B(n4013), .Y(n4011) );
  OR2X2 U4643 ( .A(n4032), .B(n4033), .Y(n4010) );
  OR2X2 U4659 ( .A(n4055), .B(n4056), .Y(n4054) );
  OR2X2 U4672 ( .A(n4075), .B(n4076), .Y(n4053) );
  OR2X2 U4688 ( .A(n4098), .B(n4099), .Y(n4097) );
  AND2X2 U4698 ( .A(n10913), .B(n4113), .Y(n3695) );
  AND2X2 U4699 ( .A(n10909), .B(n4113), .Y(n3694) );
  AND2X2 U4701 ( .A(n10913), .B(n4114), .Y(n3697) );
  AND2X2 U4704 ( .A(n10909), .B(n4114), .Y(n3696) );
  AND2X2 U4716 ( .A(n10914), .B(n4108), .Y(n3712) );
  AND2X2 U4717 ( .A(n10910), .B(n4108), .Y(n3711) );
  AND2X2 U4719 ( .A(n10914), .B(n4112), .Y(n3714) );
  AND2X2 U4722 ( .A(n10910), .B(n4112), .Y(n3713) );
  OR2X2 U4725 ( .A(n4132), .B(n4133), .Y(n4096) );
  AND2X2 U4735 ( .A(n10915), .B(n4108), .Y(n3731) );
  AND2X2 U4736 ( .A(n10911), .B(n4108), .Y(n3730) );
  AND2X2 U4738 ( .A(n10915), .B(n4112), .Y(n3733) );
  AND2X2 U4741 ( .A(n10911), .B(n4112), .Y(n3732) );
  AND2X2 U4749 ( .A(\U_0/U_1/U_1/readptr[2] ), .B(n9333), .Y(n4112) );
  AND2X2 U4753 ( .A(\U_0/U_1/U_1/readptr[2] ), .B(\U_0/U_1/U_1/readptr[1] ), 
        .Y(n4108) );
  AND2X2 U4755 ( .A(n10912), .B(n4114), .Y(n3748) );
  AND2X2 U4756 ( .A(n4114), .B(n10916), .Y(n3747) );
  AND2X2 U4759 ( .A(n4113), .B(n10912), .Y(n3750) );
  AND2X2 U4763 ( .A(n4113), .B(n10916), .Y(n3749) );
  AND2X2 U5558 ( .A(n4490), .B(n9502), .Y(n4405) );
  AND2X2 U5560 ( .A(n4491), .B(n9503), .Y(n4426) );
  AND2X2 U5583 ( .A(n3402), .B(n4500), .Y(n3405) );
  AND2X2 U5940 ( .A(n9410), .B(n4831), .Y(n4830) );
  AND2X2 U5955 ( .A(n9410), .B(n4847), .Y(n4846) );
  AND2X2 U5970 ( .A(n9411), .B(n4862), .Y(n4861) );
  AND2X2 U5985 ( .A(n9411), .B(n4877), .Y(n4876) );
  AND2X2 U6000 ( .A(n9411), .B(n4892), .Y(n4891) );
  AND2X2 U6015 ( .A(n9411), .B(n4907), .Y(n4906) );
  AND2X2 U6030 ( .A(n9411), .B(n4922), .Y(n4921) );
  AND2X2 U6039 ( .A(n4694), .B(n10756), .Y(n4821) );
  AND2X2 U6040 ( .A(n4930), .B(n4820), .Y(n4694) );
  AND2X2 U6047 ( .A(n9411), .B(n4939), .Y(n4938) );
  AND2X2 U6054 ( .A(n4820), .B(n10756), .Y(n4837) );
  AND2X2 U6063 ( .A(n9411), .B(n4955), .Y(n4954) );
  AND2X2 U6078 ( .A(n9411), .B(n4970), .Y(n4969) );
  AND2X2 U6093 ( .A(n9410), .B(n4984), .Y(n4983) );
  AND2X2 U6108 ( .A(n9410), .B(n4998), .Y(n4997) );
  AND2X2 U6123 ( .A(n9410), .B(n5012), .Y(n5011) );
  AND2X2 U6138 ( .A(n9410), .B(n5026), .Y(n5025) );
  AND2X2 U6153 ( .A(n9410), .B(n5040), .Y(n5039) );
  AND2X2 U6168 ( .A(n9410), .B(n5054), .Y(n5053) );
  AND2X2 U6175 ( .A(n5060), .B(\U_0/U_0/U_1/U_8/address[3] ), .Y(n4961) );
  AND2X2 U6184 ( .A(n9410), .B(n5070), .Y(n5069) );
  AND2X2 U6199 ( .A(n9410), .B(n5085), .Y(n5084) );
  AND2X2 U6214 ( .A(n9410), .B(n5099), .Y(n5098) );
  AND2X2 U6229 ( .A(n9410), .B(n5113), .Y(n5112) );
  AND2X2 U6244 ( .A(n9410), .B(n5127), .Y(n5126) );
  AND2X2 U6259 ( .A(n9410), .B(n5141), .Y(n5140) );
  AND2X2 U6274 ( .A(n9410), .B(n5155), .Y(n5154) );
  AND2X2 U6283 ( .A(n4945), .B(n10756), .Y(n5061) );
  AND2X2 U6284 ( .A(n5060), .B(n4930), .Y(n4945) );
  AND2X2 U6291 ( .A(n9410), .B(n5169), .Y(n5168) );
  AND2X2 U6298 ( .A(n5060), .B(n10756), .Y(n5076) );
  AND2X2 U6308 ( .A(n9410), .B(n5185), .Y(n5184) );
  AND2X2 U6323 ( .A(n9410), .B(n5200), .Y(n5199) );
  AND2X2 U6338 ( .A(n9410), .B(n5214), .Y(n5213) );
  AND2X2 U6353 ( .A(n9410), .B(n5228), .Y(n5227) );
  AND2X2 U6368 ( .A(n9410), .B(n5242), .Y(n5241) );
  AND2X2 U6383 ( .A(n9410), .B(n5256), .Y(n5255) );
  AND2X2 U6398 ( .A(n9410), .B(n5270), .Y(n5269) );
  AND2X2 U6413 ( .A(n9410), .B(n5284), .Y(n5283) );
  AND2X2 U6420 ( .A(n5290), .B(\U_0/U_0/U_1/U_8/address[3] ), .Y(n5191) );
  AND2X2 U6429 ( .A(n9410), .B(n5300), .Y(n5299) );
  AND2X2 U6444 ( .A(n9410), .B(n5315), .Y(n5314) );
  AND2X2 U6459 ( .A(n9410), .B(n5329), .Y(n5328) );
  AND2X2 U6474 ( .A(n9410), .B(n5343), .Y(n5342) );
  AND2X2 U6489 ( .A(n9410), .B(n5357), .Y(n5356) );
  AND2X2 U6504 ( .A(n9410), .B(n5371), .Y(n5370) );
  AND2X2 U6519 ( .A(n9410), .B(n5385), .Y(n5384) );
  AND2X2 U6528 ( .A(n5176), .B(n10756), .Y(n5291) );
  AND2X2 U6529 ( .A(n5290), .B(n4930), .Y(n5176) );
  AND2X2 U6536 ( .A(n9410), .B(n5399), .Y(n5398) );
  AND2X2 U6543 ( .A(n5290), .B(n10756), .Y(n5306) );
  AND2X2 U6553 ( .A(n9410), .B(n5415), .Y(n5414) );
  AND2X2 U6568 ( .A(n9410), .B(n5430), .Y(n5429) );
  AND2X2 U6583 ( .A(n9410), .B(n5444), .Y(n5443) );
  AND2X2 U6598 ( .A(n9410), .B(n5458), .Y(n5457) );
  AND2X2 U6613 ( .A(n9410), .B(n5472), .Y(n5471) );
  AND2X2 U6628 ( .A(n9411), .B(n5486), .Y(n5485) );
  AND2X2 U6643 ( .A(n9410), .B(n5500), .Y(n5499) );
  AND2X2 U6659 ( .A(n9410), .B(n5514), .Y(n5513) );
  AND2X2 U6666 ( .A(n5520), .B(\U_0/U_0/U_1/U_8/address[3] ), .Y(n5421) );
  AND2X2 U6675 ( .A(n4678), .B(n5530), .Y(n5529) );
  AND2X2 U6691 ( .A(n4678), .B(n5545), .Y(n5544) );
  AND2X2 U6707 ( .A(n4678), .B(n5560), .Y(n5559) );
  AND2X2 U6723 ( .A(n4678), .B(n5574), .Y(n5573) );
  AND2X2 U6791 ( .A(n5406), .B(n10756), .Y(n5521) );
  AND2X2 U6792 ( .A(n5520), .B(n4930), .Y(n5406) );
  AND2X2 U6824 ( .A(n5520), .B(n10756), .Y(n5536) );
  AND2X2 U6878 ( .A(n9207), .B(n5663), .Y(n5648) );
  AND2X2 U6935 ( .A(n9207), .B(n5698), .Y(n5643) );
  OR2X2 U6956 ( .A(n5725), .B(n5726), .Y(n9145) );
  AND2X2 U6985 ( .A(n5737), .B(n10568), .Y(n5752) );
  OR2X2 U7010 ( .A(\U_0/U_0/U_1/U_7/state[5] ), .B(\U_0/U_0/U_1/U_7/state[6] ), 
        .Y(n5770) );
  AND2X2 U7039 ( .A(n5779), .B(n5796), .Y(n5781) );
  OR2X2 U7042 ( .A(n5797), .B(n5798), .Y(n5796) );
  OR2X2 U7052 ( .A(PARITY_ERROR), .B(PARITY_ERROR1), .Y(c_parity_error) );
  OR2X2 U7081 ( .A(n5828), .B(n5829), .Y(\U_1/U_3/U_3/nextstate [0]) );
  AND2X2 U7083 ( .A(n237), .B(n187), .Y(n5813) );
  OR2X2 U7084 ( .A(n236), .B(\U_1/U_3/U_3/state[0] ), .Y(n187) );
  AND2X2 U7091 ( .A(n5835), .B(n5816), .Y(n5834) );
  AND2X2 U7110 ( .A(n5850), .B(\U_1/U_3/U_0/state[2] ), .Y(n5845) );
  OR2X2 U7111 ( .A(n5851), .B(n5852), .Y(\U_1/U_3/U_0/nextstate [1]) );
  OR2X2 U7136 ( .A(n5864), .B(n11621), .Y(n784) );
  AND2X2 U7148 ( .A(n5885), .B(n5886), .Y(n5884) );
  AND2X2 U7201 ( .A(n5914), .B(\U_1/U_2/U_7/state ), .Y(n5911) );
  AND2X2 U7281 ( .A(n5986), .B(n9698), .Y(\U_1/U_2/U_1/N32 ) );
  AND2X2 U7351 ( .A(\U_1/U_1/U_1/N337 ), .B(n9318), .Y(\U_1/U_1/U_1/N347 ) );
  AND2X2 U7352 ( .A(\U_1/U_1/U_1/N336 ), .B(n9318), .Y(\U_1/U_1/U_1/N346 ) );
  AND2X2 U7353 ( .A(\U_1/U_1/U_1/N335 ), .B(n9318), .Y(\U_1/U_1/U_1/N345 ) );
  AND2X2 U7354 ( .A(\U_1/U_1/U_1/N334 ), .B(n9318), .Y(\U_1/U_1/U_1/N344 ) );
  AND2X2 U7355 ( .A(\U_1/U_1/U_1/N333 ), .B(n9318), .Y(\U_1/U_1/U_1/N343 ) );
  AND2X2 U7356 ( .A(\U_1/U_1/U_1/N193 ), .B(n9318), .Y(\U_1/U_1/U_1/N342 ) );
  AND2X2 U7357 ( .A(\U_1/U_1/U_1/N192 ), .B(n9318), .Y(\U_1/U_1/U_1/N341 ) );
  AND2X2 U7358 ( .A(\U_1/U_1/U_1/N191 ), .B(n9318), .Y(\U_1/U_1/U_1/N340 ) );
  AND2X2 U7359 ( .A(\U_1/U_1/U_1/N190 ), .B(n9318), .Y(\U_1/U_1/U_1/N339 ) );
  AND2X2 U7360 ( .A(\U_1/U_1/U_1/N189 ), .B(n9318), .Y(\U_1/U_1/U_1/N338 ) );
  AND2X2 U7361 ( .A(\U_1/U_1/U_1/N194 ), .B(\U_1/U_1/R_ENABLE ), .Y(
        \U_1/U_1/U_1/N195 ) );
  AND2X2 U7403 ( .A(n6038), .B(n6039), .Y(n6037) );
  AND2X2 U7424 ( .A(n11326), .B(\U_1/U_0/U_1/U_2/state[0] ), .Y(n6050) );
  AND2X2 U7439 ( .A(\U_1/U_0/U_1/U_2/N30 ), .B(\U_1/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_1/U_0/U_1/U_2/N38 ) );
  AND2X2 U7440 ( .A(\U_1/U_0/U_1/U_2/N29 ), .B(\U_1/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_1/U_0/U_1/U_2/N37 ) );
  AND2X2 U7441 ( .A(\U_1/U_0/U_1/U_2/N28 ), .B(\U_1/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_1/U_0/U_1/U_2/N36 ) );
  AND2X2 U7442 ( .A(\U_1/U_0/U_1/U_2/N27 ), .B(\U_1/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_1/U_0/U_1/U_2/N35 ) );
  AND2X2 U7443 ( .A(\U_1/U_0/U_1/U_2/N26 ), .B(\U_1/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_1/U_0/U_1/U_2/N34 ) );
  AND2X2 U7444 ( .A(\U_1/U_0/U_1/U_2/N25 ), .B(\U_1/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_1/U_0/U_1/U_2/N33 ) );
  AND2X2 U7445 ( .A(\U_1/U_0/U_1/U_2/N24 ), .B(\U_1/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_1/U_0/U_1/U_2/N32 ) );
  OR2X2 U7446 ( .A(\U_1/U_0/U_1/U_2/N23 ), .B(n11323), .Y(
        \U_1/U_0/U_1/U_2/N31 ) );
  OR2X2 U7495 ( .A(n6099), .B(n11895), .Y(n6098) );
  AND2X2 U7552 ( .A(n1001), .B(n1018), .Y(n6153) );
  OR2X2 U7568 ( .A(n6167), .B(n6168), .Y(\U_1/U_0/U_0/nextState [4]) );
  AND2X2 U7605 ( .A(n6194), .B(n6215), .Y(n6210) );
  OR2X2 U7614 ( .A(n6223), .B(n6224), .Y(\U_1/U_0/U_0/nextState [0]) );
  OR2X2 U7631 ( .A(n6238), .B(\U_1/U_0/U_1/U_8/state[2] ), .Y(n3201) );
  AND2X2 U7708 ( .A(n6271), .B(n6215), .Y(n6243) );
  OR2X2 U7913 ( .A(n6392), .B(n6393), .Y(\U_0/U_3/U_3/nextstate [0]) );
  AND2X2 U7915 ( .A(n522), .B(n473), .Y(n6377) );
  AND2X2 U7923 ( .A(n6399), .B(n6380), .Y(n6398) );
  AND2X2 U7941 ( .A(n6414), .B(\U_0/U_3/U_0/state[2] ), .Y(n6409) );
  OR2X2 U7942 ( .A(n6415), .B(n6416), .Y(\U_0/U_3/U_0/nextstate [1]) );
  OR2X2 U7967 ( .A(n6428), .B(n10869), .Y(n3306) );
  AND2X2 U7979 ( .A(n6449), .B(n6450), .Y(n6448) );
  AND2X2 U8031 ( .A(n6478), .B(\U_0/U_2/U_7/state ), .Y(n6475) );
  AND2X2 U8111 ( .A(n6550), .B(n9690), .Y(\U_0/U_2/U_1/N32 ) );
  AND2X2 U8182 ( .A(\U_0/U_1/U_1/N337 ), .B(n9353), .Y(\U_0/U_1/U_1/N347 ) );
  AND2X2 U8183 ( .A(\U_0/U_1/U_1/N336 ), .B(n9353), .Y(\U_0/U_1/U_1/N346 ) );
  AND2X2 U8184 ( .A(\U_0/U_1/U_1/N335 ), .B(n9353), .Y(\U_0/U_1/U_1/N345 ) );
  AND2X2 U8185 ( .A(\U_0/U_1/U_1/N334 ), .B(n9353), .Y(\U_0/U_1/U_1/N344 ) );
  AND2X2 U8186 ( .A(\U_0/U_1/U_1/N333 ), .B(n9353), .Y(\U_0/U_1/U_1/N343 ) );
  AND2X2 U8187 ( .A(\U_0/U_1/U_1/N193 ), .B(n9353), .Y(\U_0/U_1/U_1/N342 ) );
  AND2X2 U8188 ( .A(\U_0/U_1/U_1/N192 ), .B(n9353), .Y(\U_0/U_1/U_1/N341 ) );
  AND2X2 U8189 ( .A(\U_0/U_1/U_1/N191 ), .B(n9353), .Y(\U_0/U_1/U_1/N340 ) );
  AND2X2 U8190 ( .A(\U_0/U_1/U_1/N190 ), .B(n9353), .Y(\U_0/U_1/U_1/N339 ) );
  AND2X2 U8191 ( .A(\U_0/U_1/U_1/N189 ), .B(n9353), .Y(\U_0/U_1/U_1/N338 ) );
  AND2X2 U8192 ( .A(\U_0/U_1/U_1/N194 ), .B(\U_0/U_1/R_ENABLE ), .Y(
        \U_0/U_1/U_1/N195 ) );
  AND2X2 U8234 ( .A(n6602), .B(n6603), .Y(n6601) );
  AND2X2 U8255 ( .A(n10574), .B(\U_0/U_0/U_1/U_2/state[0] ), .Y(n6614) );
  AND2X2 U8270 ( .A(\U_0/U_0/U_1/U_2/N30 ), .B(\U_0/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_0/U_0/U_1/U_2/N38 ) );
  AND2X2 U8271 ( .A(\U_0/U_0/U_1/U_2/N29 ), .B(\U_0/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_0/U_0/U_1/U_2/N37 ) );
  AND2X2 U8272 ( .A(\U_0/U_0/U_1/U_2/N28 ), .B(\U_0/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_0/U_0/U_1/U_2/N36 ) );
  AND2X2 U8273 ( .A(\U_0/U_0/U_1/U_2/N27 ), .B(\U_0/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_0/U_0/U_1/U_2/N35 ) );
  AND2X2 U8274 ( .A(\U_0/U_0/U_1/U_2/N26 ), .B(\U_0/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_0/U_0/U_1/U_2/N34 ) );
  AND2X2 U8275 ( .A(\U_0/U_0/U_1/U_2/N25 ), .B(\U_0/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_0/U_0/U_1/U_2/N33 ) );
  AND2X2 U8276 ( .A(\U_0/U_0/U_1/U_2/N24 ), .B(\U_0/U_0/U_1/U_2/timerRunning ), 
        .Y(\U_0/U_0/U_1/U_2/N32 ) );
  OR2X2 U8277 ( .A(\U_0/U_0/U_1/U_2/N23 ), .B(n10571), .Y(
        \U_0/U_0/U_1/U_2/N31 ) );
  AND2X2 U8338 ( .A(n9190), .B(n3583), .Y(n6663) );
  AND2X2 U8435 ( .A(n6759), .B(n6718), .Y(n6774) );
  OR2X2 U8445 ( .A(n6779), .B(n11154), .Y(n6768) );
  OR2X2 U8453 ( .A(n6786), .B(n6787), .Y(\U_0/U_0/U_0/nextState [0]) );
  OR2X2 U8456 ( .A(n3569), .B(n6790), .Y(n6785) );
  OR2X2 U8469 ( .A(n6801), .B(\U_0/U_0/U_1/U_8/state[2] ), .Y(n5702) );
  AND2X2 U8504 ( .A(n6941), .B(n567), .Y(n6806) );
  rmedt_square_DW01_inc_1 \U_1/U_0/U_1/U_7/add_39  ( .A({
        \U_1/U_0/U_1/U_7/nextState[7] , \U_1/U_0/U_1/U_7/nextState[6] , 
        \U_1/U_0/U_1/U_7/nextState[5] , \U_1/U_0/U_1/U_7/nextState[4] , 
        \U_1/U_0/U_1/U_7/nextState[3] , \U_1/U_0/U_1/U_7/nextState[2] , 
        \U_1/U_0/U_1/U_7/nextState[1] , \U_1/U_0/U_1/U_7/nextState[0] }), 
        .SUM({\U_1/U_0/U_1/U_7/N33 , \U_1/U_0/U_1/U_7/N32 , 
        \U_1/U_0/U_1/U_7/N31 , \U_1/U_0/U_1/U_7/N30 , \U_1/U_0/U_1/U_7/N29 , 
        \U_1/U_0/U_1/U_7/N28 , \U_1/U_0/U_1/U_7/N27 , \U_1/U_0/U_1/U_7/N26 })
         );
  rmedt_square_DW01_add_2 \U_1/U_0/U_0/add_377  ( .A({\U_1/U_0/U_0/temp[7] , 
        \U_1/U_0/U_0/temp[6] , \U_1/U_0/U_0/temp[5] , \U_1/U_0/U_0/temp[4] , 
        \U_1/U_0/U_0/temp[3] , \U_1/U_0/U_0/temp[2] , \U_1/U_0/U_0/temp[1] , 
        \U_1/U_0/U_0/temp[0] }), .B({\U_1/U_0/U_0/extratemp[7] , 
        \U_1/U_0/U_0/extratemp[6] , \U_1/U_0/U_0/extratemp[5] , 
        \U_1/U_0/U_0/extratemp[4] , \U_1/U_0/U_0/extratemp[3] , 
        \U_1/U_0/U_0/extratemp[2] , \U_1/U_0/U_0/extratemp[1] , 
        \U_1/U_0/U_0/extratemp[0] }), .CI(1'b0), .SUM({\U_1/U_0/U_0/N527 , 
        \U_1/U_0/U_0/N526 , \U_1/U_0/U_0/N525 , \U_1/U_0/U_0/N524 , 
        \U_1/U_0/U_0/N523 , \U_1/U_0/U_0/N522 , \U_1/U_0/U_0/N521 , 
        \U_1/U_0/U_0/N520 }) );
  rmedt_square_DW01_add_3 \U_1/U_0/U_0/add_337  ( .A({\U_1/U_0/U_0/intj[7] , 
        \U_1/U_0/U_0/intj[6] , \U_1/U_0/U_0/intj[5] , \U_1/U_0/U_0/intj[4] , 
        \U_1/U_0/U_0/intj[3] , \U_1/U_0/U_0/intj[2] , \U_1/U_0/U_0/intj[1] , 
        \U_1/U_0/U_0/intj[0] }), .B(DATA_IN_S), .CI(1'b0), .SUM({
        \U_1/U_0/U_0/N519 , \U_1/U_0/U_0/N518 , \U_1/U_0/U_0/N517 , 
        \U_1/U_0/U_0/N516 , \U_1/U_0/U_0/N515 , \U_1/U_0/U_0/N514 , 
        \U_1/U_0/U_0/N513 , \U_1/U_0/U_0/N512 }) );
  rmedt_square_DW01_inc_2 \U_1/U_0/U_0/add_289  ( .A({\U_1/U_0/U_0/si[7] , 
        \U_1/U_0/U_0/si[6] , \U_1/U_0/U_0/si[5] , \U_1/U_0/U_0/si[4] , 
        \U_1/U_0/U_0/si[3] , \U_1/U_0/U_0/si[2] , \U_1/U_0/U_0/si[1] , 
        \U_1/U_0/U_0/si[0] }), .SUM({\U_1/U_0/U_0/N431 , \U_1/U_0/U_0/N430 , 
        \U_1/U_0/U_0/N429 , \U_1/U_0/U_0/N428 , \U_1/U_0/U_0/N427 , 
        \U_1/U_0/U_0/N426 , \U_1/U_0/U_0/N425 , \U_1/U_0/U_0/N424 }) );
  rmedt_square_DW01_inc_3 \U_1/U_0/U_0/add_263  ( .A({
        \U_1/U_0/U_0/prefillCounter[7] , \U_1/U_0/U_0/prefillCounter[6] , 
        \U_1/U_0/U_0/prefillCounter[5] , \U_1/U_0/U_0/prefillCounter[4] , 
        \U_1/U_0/U_0/prefillCounter[3] , \U_1/U_0/U_0/prefillCounter[2] , 
        \U_1/U_0/U_0/prefillCounter[1] , \U_1/U_0/U_0/prefillCounter[0] }), 
        .SUM({\U_1/U_0/U_0/N414 , \U_1/U_0/U_0/N413 , \U_1/U_0/U_0/N412 , 
        \U_1/U_0/U_0/N411 , \U_1/U_0/U_0/N410 , \U_1/U_0/U_0/N409 , 
        \U_1/U_0/U_0/N408 , \U_1/U_0/U_0/N407 }) );
  rmedt_square_DW01_inc_5 \U_0/U_0/U_1/U_7/add_39  ( .A({
        \U_0/U_0/U_1/U_7/nextState[7] , \U_0/U_0/U_1/U_7/nextState[6] , 
        \U_0/U_0/U_1/U_7/nextState[5] , \U_0/U_0/U_1/U_7/nextState[4] , 
        \U_0/U_0/U_1/U_7/nextState[3] , \U_0/U_0/U_1/U_7/nextState[2] , 
        \U_0/U_0/U_1/U_7/nextState[1] , \U_0/U_0/U_1/U_7/nextState[0] }), 
        .SUM({\U_0/U_0/U_1/U_7/N33 , \U_0/U_0/U_1/U_7/N32 , 
        \U_0/U_0/U_1/U_7/N31 , \U_0/U_0/U_1/U_7/N30 , \U_0/U_0/U_1/U_7/N29 , 
        \U_0/U_0/U_1/U_7/N28 , \U_0/U_0/U_1/U_7/N27 , \U_0/U_0/U_1/U_7/N26 })
         );
  rmedt_square_DW01_add_6 \U_0/U_0/U_0/add_377  ( .A({\U_0/U_0/U_0/temp[7] , 
        \U_0/U_0/U_0/temp[6] , \U_0/U_0/U_0/temp[5] , \U_0/U_0/U_0/temp[4] , 
        \U_0/U_0/U_0/temp[3] , \U_0/U_0/U_0/temp[2] , \U_0/U_0/U_0/temp[1] , 
        \U_0/U_0/U_0/temp[0] }), .B({\U_0/U_0/U_0/extratemp[7] , 
        \U_0/U_0/U_0/extratemp[6] , \U_0/U_0/U_0/extratemp[5] , 
        \U_0/U_0/U_0/extratemp[4] , \U_0/U_0/U_0/extratemp[3] , 
        \U_0/U_0/U_0/extratemp[2] , \U_0/U_0/U_0/extratemp[1] , 
        \U_0/U_0/U_0/extratemp[0] }), .CI(1'b0), .SUM({\U_0/U_0/U_0/N527 , 
        \U_0/U_0/U_0/N526 , \U_0/U_0/U_0/N525 , \U_0/U_0/U_0/N524 , 
        \U_0/U_0/U_0/N523 , \U_0/U_0/U_0/N522 , \U_0/U_0/U_0/N521 , 
        \U_0/U_0/U_0/N520 }) );
  rmedt_square_DW01_add_7 \U_0/U_0/U_0/add_337  ( .A({\U_0/U_0/U_0/intj[7] , 
        \U_0/U_0/U_0/intj[6] , \U_0/U_0/U_0/intj[5] , \U_0/U_0/U_0/intj[4] , 
        \U_0/U_0/U_0/intj[3] , \U_0/U_0/U_0/intj[2] , \U_0/U_0/U_0/intj[1] , 
        \U_0/U_0/U_0/intj[0] }), .B(DATA_IN_H), .CI(1'b0), .SUM({
        \U_0/U_0/U_0/N519 , \U_0/U_0/U_0/N518 , \U_0/U_0/U_0/N517 , 
        \U_0/U_0/U_0/N516 , \U_0/U_0/U_0/N515 , \U_0/U_0/U_0/N514 , 
        \U_0/U_0/U_0/N513 , \U_0/U_0/U_0/N512 }) );
  rmedt_square_DW01_inc_6 \U_0/U_0/U_0/add_289  ( .A({\U_0/U_0/U_0/si[7] , 
        \U_0/U_0/U_0/si[6] , \U_0/U_0/U_0/si[5] , \U_0/U_0/U_0/si[4] , 
        \U_0/U_0/U_0/si[3] , \U_0/U_0/U_0/si[2] , \U_0/U_0/U_0/si[1] , 
        \U_0/U_0/U_0/si[0] }), .SUM({\U_0/U_0/U_0/N431 , \U_0/U_0/U_0/N430 , 
        \U_0/U_0/U_0/N429 , \U_0/U_0/U_0/N428 , \U_0/U_0/U_0/N427 , 
        \U_0/U_0/U_0/N426 , \U_0/U_0/U_0/N425 , \U_0/U_0/U_0/N424 }) );
  rmedt_square_DW01_inc_7 \U_0/U_0/U_0/add_263  ( .A({
        \U_0/U_0/U_0/prefillCounter[7] , \U_0/U_0/U_0/prefillCounter[6] , 
        \U_0/U_0/U_0/prefillCounter[5] , \U_0/U_0/U_0/prefillCounter[4] , 
        \U_0/U_0/U_0/prefillCounter[3] , \U_0/U_0/U_0/prefillCounter[2] , 
        \U_0/U_0/U_0/prefillCounter[1] , \U_0/U_0/U_0/prefillCounter[0] }), 
        .SUM({\U_0/U_0/U_0/N414 , \U_0/U_0/U_0/N413 , \U_0/U_0/U_0/N412 , 
        \U_0/U_0/U_0/N411 , \U_0/U_0/U_0/N410 , \U_0/U_0/U_0/N409 , 
        \U_0/U_0/U_0/N408 , \U_0/U_0/U_0/N407 }) );
  rmedt_square_DW01_inc_8 r2041 ( .A({\U_1/U_3/U_3/N188 , 
        \U_1/U_3/U_3/count[5] , \U_1/U_3/U_3/count[4] , \U_1/U_3/U_3/count[3] , 
        \U_1/U_3/U_3/count[2] , \U_1/U_3/U_3/count[1] , \U_1/U_3/U_3/count[0] }), .SUM({\U_1/U_3/U_3/N65 , \U_1/U_3/U_3/N64 , \U_1/U_3/U_3/N63 , 
        \U_1/U_3/U_3/N62 , \U_1/U_3/U_3/N61 , \U_1/U_3/U_3/N60 , 
        \U_1/U_3/U_3/N59 }) );
  rmedt_square_DW01_add_9 r2023 ( .A({\U_1/U_0/U_1/U_8/parityAccumulator[7] , 
        \U_1/U_0/U_1/U_8/parityAccumulator[6] , 
        \U_1/U_0/U_1/U_8/parityAccumulator[5] , 
        \U_1/U_0/U_1/U_8/parityAccumulator[4] , 
        \U_1/U_0/U_1/U_8/parityAccumulator[3] , 
        \U_1/U_0/U_1/U_8/parityAccumulator[2] , 
        \U_1/U_0/U_1/U_8/parityAccumulator[1] , 
        \U_1/U_0/U_1/U_8/parityAccumulator[0] }), .B({
        \U_1/U_0/U_1/RCV_DATA [7:3], n9474, \U_1/U_0/U_1/RCV_DATA [1], n9479}), 
        .CI(1'b0), .SUM({\U_1/U_0/U_1/U_8/N1799 , \U_1/U_0/U_1/U_8/N1798 , 
        \U_1/U_0/U_1/U_8/N1797 , \U_1/U_0/U_1/U_8/N1796 , 
        \U_1/U_0/U_1/U_8/N1795 , \U_1/U_0/U_1/U_8/N1794 , 
        \U_1/U_0/U_1/U_8/N1793 , \U_1/U_0/U_1/U_8/N1792 }) );
  rmedt_square_DW01_inc_10 r2017 ( .A({\U_1/U_0/U_0/inti[7] , 
        \U_1/U_0/U_0/inti[6] , \U_1/U_0/U_0/inti[5] , \U_1/U_0/U_0/inti[4] , 
        \U_1/U_0/U_0/inti[3] , \U_1/U_0/U_0/inti[2] , \U_1/U_0/U_0/inti[1] , 
        \U_1/U_0/U_0/inti[0] }), .SUM({\U_1/U_0/U_0/N503 , \U_1/U_0/U_0/N502 , 
        \U_1/U_0/U_0/N501 , \U_1/U_0/U_0/N500 , \U_1/U_0/U_0/N499 , 
        \U_1/U_0/U_0/N498 , \U_1/U_0/U_0/N497 , \U_1/U_0/U_0/N496 }) );
  rmedt_square_DW01_inc_11 r2007 ( .A({\U_0/U_3/U_3/N188 , 
        \U_0/U_3/U_3/count[5] , \U_0/U_3/U_3/count[4] , \U_0/U_3/U_3/count[3] , 
        \U_0/U_3/U_3/count[2] , \U_0/U_3/U_3/count[1] , \U_0/U_3/U_3/count[0] }), .SUM({\U_0/U_3/U_3/N65 , \U_0/U_3/U_3/N64 , \U_0/U_3/U_3/N63 , 
        \U_0/U_3/U_3/N62 , \U_0/U_3/U_3/N61 , \U_0/U_3/U_3/N60 , 
        \U_0/U_3/U_3/N59 }) );
  rmedt_square_DW01_add_11 r1989 ( .A({\U_0/U_0/U_1/U_8/parityAccumulator[7] , 
        \U_0/U_0/U_1/U_8/parityAccumulator[6] , 
        \U_0/U_0/U_1/U_8/parityAccumulator[5] , 
        \U_0/U_0/U_1/U_8/parityAccumulator[4] , 
        \U_0/U_0/U_1/U_8/parityAccumulator[3] , 
        \U_0/U_0/U_1/U_8/parityAccumulator[2] , 
        \U_0/U_0/U_1/U_8/parityAccumulator[1] , 
        \U_0/U_0/U_1/U_8/parityAccumulator[0] }), .B({
        \U_0/U_0/U_1/RCV_DATA [7:3], n9481, \U_0/U_0/U_1/RCV_DATA [1], n9486}), 
        .CI(1'b0), .SUM({\U_0/U_0/U_1/U_8/N1799 , \U_0/U_0/U_1/U_8/N1798 , 
        \U_0/U_0/U_1/U_8/N1797 , \U_0/U_0/U_1/U_8/N1796 , 
        \U_0/U_0/U_1/U_8/N1795 , \U_0/U_0/U_1/U_8/N1794 , 
        \U_0/U_0/U_1/U_8/N1793 , \U_0/U_0/U_1/U_8/N1792 }) );
  rmedt_square_DW01_inc_13 r1983 ( .A({\U_0/U_0/U_0/inti[7] , 
        \U_0/U_0/U_0/inti[6] , \U_0/U_0/U_0/inti[5] , \U_0/U_0/U_0/inti[4] , 
        \U_0/U_0/U_0/inti[3] , \U_0/U_0/U_0/inti[2] , \U_0/U_0/U_0/inti[1] , 
        \U_0/U_0/U_0/inti[0] }), .SUM({\U_0/U_0/U_0/N503 , \U_0/U_0/U_0/N502 , 
        \U_0/U_0/U_0/N501 , \U_0/U_0/U_0/N500 , \U_0/U_0/U_0/N499 , 
        \U_0/U_0/U_0/N498 , \U_0/U_0/U_0/N497 , \U_0/U_0/U_0/N496 }) );
  rmedt_square_DW01_add_15 \add_1_root_add_0_root_U_0/U_0/U_0/add_302_2  ( .A(
        DATA_IN_H), .B({\U_0/U_0/U_0/sj[7] , \U_0/U_0/U_0/sj[6] , 
        \U_0/U_0/U_0/sj[5] , \U_0/U_0/U_0/sj[4] , \U_0/U_0/U_0/sj[3] , 
        \U_0/U_0/U_0/sj[2] , \U_0/U_0/U_0/sj[1] , \U_0/U_0/U_0/sj[0] }), .CI(
        1'b0), .SUM({\U_0/U_0/U_0/N456 , \U_0/U_0/U_0/N455 , 
        \U_0/U_0/U_0/N454 , \U_0/U_0/U_0/N453 , \U_0/U_0/U_0/N452 , 
        \U_0/U_0/U_0/N451 , \U_0/U_0/U_0/N450 , \U_0/U_0/U_0/N449 }) );
  rmedt_square_DW01_add_14 \add_0_root_add_0_root_U_0/U_0/U_0/add_302_2  ( .A(
        {\U_0/U_0/U_0/N472 , \U_0/U_0/U_0/N473 , \U_0/U_0/U_0/N474 , 
        \U_0/U_0/U_0/N475 , \U_0/U_0/U_0/N476 , \U_0/U_0/U_0/N477 , 
        \U_0/U_0/U_0/N478 , \U_0/U_0/U_0/N479 }), .B({\U_0/U_0/U_0/N456 , 
        \U_0/U_0/U_0/N455 , \U_0/U_0/U_0/N454 , \U_0/U_0/U_0/N453 , 
        \U_0/U_0/U_0/N452 , \U_0/U_0/U_0/N451 , \U_0/U_0/U_0/N450 , 
        \U_0/U_0/U_0/N449 }), .CI(1'b0), .SUM({\U_0/U_0/U_0/N487 , 
        \U_0/U_0/U_0/N486 , \U_0/U_0/U_0/N485 , \U_0/U_0/U_0/N484 , 
        \U_0/U_0/U_0/N483 , \U_0/U_0/U_0/N482 , \U_0/U_0/U_0/N481 , 
        \U_0/U_0/U_0/N480 }) );
  rmedt_square_DW01_add_13 \add_1_root_add_0_root_U_1/U_0/U_0/add_302_2  ( .A(
        DATA_IN_S), .B({\U_1/U_0/U_0/sj[7] , \U_1/U_0/U_0/sj[6] , 
        \U_1/U_0/U_0/sj[5] , \U_1/U_0/U_0/sj[4] , \U_1/U_0/U_0/sj[3] , 
        \U_1/U_0/U_0/sj[2] , \U_1/U_0/U_0/sj[1] , \U_1/U_0/U_0/sj[0] }), .CI(
        1'b0), .SUM({\U_1/U_0/U_0/N456 , \U_1/U_0/U_0/N455 , 
        \U_1/U_0/U_0/N454 , \U_1/U_0/U_0/N453 , \U_1/U_0/U_0/N452 , 
        \U_1/U_0/U_0/N451 , \U_1/U_0/U_0/N450 , \U_1/U_0/U_0/N449 }) );
  rmedt_square_DW01_add_12 \add_0_root_add_0_root_U_1/U_0/U_0/add_302_2  ( .A(
        {\U_1/U_0/U_0/N472 , \U_1/U_0/U_0/N473 , \U_1/U_0/U_0/N474 , 
        \U_1/U_0/U_0/N475 , \U_1/U_0/U_0/N476 , \U_1/U_0/U_0/N477 , 
        \U_1/U_0/U_0/N478 , \U_1/U_0/U_0/N479 }), .B({\U_1/U_0/U_0/N456 , 
        \U_1/U_0/U_0/N455 , \U_1/U_0/U_0/N454 , \U_1/U_0/U_0/N453 , 
        \U_1/U_0/U_0/N452 , \U_1/U_0/U_0/N451 , \U_1/U_0/U_0/N450 , 
        \U_1/U_0/U_0/N449 }), .CI(1'b0), .SUM({\U_1/U_0/U_0/N487 , 
        \U_1/U_0/U_0/N486 , \U_1/U_0/U_0/N485 , \U_1/U_0/U_0/N484 , 
        \U_1/U_0/U_0/N483 , \U_1/U_0/U_0/N482 , \U_1/U_0/U_0/N481 , 
        \U_1/U_0/U_0/N480 }) );
  FAX1 \U_1/U_1/U_1/sub_72/U2_1  ( .A(n9290), .B(n9299), .C(
        \U_1/U_1/U_1/sub_72/carry[1] ), .YC(\U_1/U_1/U_1/sub_72/carry[2] ), 
        .YS(\U_1/U_1/U_1/N190 ) );
  FAX1 \U_1/U_1/U_1/sub_72/U2_2  ( .A(n9288), .B(n9298), .C(
        \U_1/U_1/U_1/sub_72/carry[2] ), .YC(\U_1/U_1/U_1/sub_72/carry[3] ), 
        .YS(\U_1/U_1/U_1/N191 ) );
  FAX1 \U_1/U_1/U_1/sub_72/U2_3  ( .A(n9292), .B(n9296), .C(
        \U_1/U_1/U_1/sub_72/carry[3] ), .YC(\U_1/U_1/U_1/sub_72/carry[4] ), 
        .YS(\U_1/U_1/U_1/N192 ) );
  FAX1 \U_1/U_1/U_1/sub_72/U2_4  ( .A(n9294), .B(n9295), .C(
        \U_1/U_1/U_1/sub_72/carry[4] ), .YS(\U_1/U_1/U_1/N193 ) );
  HAX1 \U_1/U_1/U_1/add_67/U1_1_1  ( .A(n9290), .B(\U_1/U_1/U_1/writeptr[0] ), 
        .YC(\U_1/U_1/U_1/add_67/carry[2] ), .YS(\U_1/U_1/U_1/N48 ) );
  HAX1 \U_1/U_1/U_1/add_67/U1_1_2  ( .A(\U_1/U_1/U_1/writeptr[2] ), .B(
        \U_1/U_1/U_1/add_67/carry[2] ), .YC(\U_1/U_1/U_1/add_67/carry[3] ), 
        .YS(\U_1/U_1/U_1/N49 ) );
  HAX1 \U_1/U_1/U_1/add_67/U1_1_3  ( .A(n9292), .B(
        \U_1/U_1/U_1/add_67/carry[3] ), .YC(\U_1/U_1/U_1/add_67/carry[4] ), 
        .YS(\U_1/U_1/U_1/N50 ) );
  FAX1 \U_0/U_1/U_1/sub_72/U2_1  ( .A(n9324), .B(n9333), .C(
        \U_0/U_1/U_1/sub_72/carry[1] ), .YC(\U_0/U_1/U_1/sub_72/carry[2] ), 
        .YS(\U_0/U_1/U_1/N190 ) );
  FAX1 \U_0/U_1/U_1/sub_72/U2_2  ( .A(n9322), .B(n9332), .C(
        \U_0/U_1/U_1/sub_72/carry[2] ), .YC(\U_0/U_1/U_1/sub_72/carry[3] ), 
        .YS(\U_0/U_1/U_1/N191 ) );
  FAX1 \U_0/U_1/U_1/sub_72/U2_3  ( .A(n9326), .B(n9330), .C(
        \U_0/U_1/U_1/sub_72/carry[3] ), .YC(\U_0/U_1/U_1/sub_72/carry[4] ), 
        .YS(\U_0/U_1/U_1/N192 ) );
  FAX1 \U_0/U_1/U_1/sub_72/U2_4  ( .A(n9328), .B(n9329), .C(
        \U_0/U_1/U_1/sub_72/carry[4] ), .YS(\U_0/U_1/U_1/N193 ) );
  HAX1 \U_0/U_1/U_1/add_67/U1_1_1  ( .A(n9324), .B(\U_0/U_1/U_1/writeptr[0] ), 
        .YC(\U_0/U_1/U_1/add_67/carry[2] ), .YS(\U_0/U_1/U_1/N48 ) );
  HAX1 \U_0/U_1/U_1/add_67/U1_1_2  ( .A(\U_0/U_1/U_1/writeptr[2] ), .B(
        \U_0/U_1/U_1/add_67/carry[2] ), .YC(\U_0/U_1/U_1/add_67/carry[3] ), 
        .YS(\U_0/U_1/U_1/N49 ) );
  HAX1 \U_0/U_1/U_1/add_67/U1_1_3  ( .A(n9326), .B(
        \U_0/U_1/U_1/add_67/carry[3] ), .YC(\U_0/U_1/U_1/add_67/carry[4] ), 
        .YS(\U_0/U_1/U_1/N50 ) );
  HAX1 \r2028/U1_1_1  ( .A(\U_1/U_1/U_1/writeptr[1] ), .B(
        \U_1/U_1/U_1/writeptr[0] ), .YC(\r2028/carry[2] ), .YS(
        \U_1/U_1/U_1/N32 ) );
  HAX1 \r2028/U1_1_2  ( .A(n9288), .B(\r2028/carry[2] ), .YC(\r2028/carry[3] ), 
        .YS(\U_1/U_1/U_1/N33 ) );
  HAX1 \r2028/U1_1_3  ( .A(\U_1/U_1/U_1/writeptr[3] ), .B(\r2028/carry[3] ), 
        .YC(\r2028/carry[4] ), .YS(\U_1/U_1/U_1/N34 ) );
  HAX1 \r1994/U1_1_1  ( .A(\U_0/U_1/U_1/writeptr[1] ), .B(
        \U_0/U_1/U_1/writeptr[0] ), .YC(\r1994/carry[2] ), .YS(
        \U_0/U_1/U_1/N32 ) );
  HAX1 \r1994/U1_1_2  ( .A(n9322), .B(\r1994/carry[2] ), .YC(\r1994/carry[3] ), 
        .YS(\U_0/U_1/U_1/N33 ) );
  HAX1 \r1994/U1_1_3  ( .A(\U_0/U_1/U_1/writeptr[3] ), .B(\r1994/carry[3] ), 
        .YC(\r1994/carry[4] ), .YS(\U_0/U_1/U_1/N34 ) );
  TBUFX1 \U_0/U_0/U_0/nfdata_tri[7]  ( .A(n6940), .EN(n6941), .Y(
        \U_0/U_0/U_0/nfdata[7] ) );
  TBUFX1 \U_0/U_0/U_0/nfdata_tri[6]  ( .A(n6939), .EN(n6941), .Y(
        \U_0/U_0/U_0/nfdata[6] ) );
  TBUFX1 \U_0/U_0/U_0/nfdata_tri[5]  ( .A(n6938), .EN(n6941), .Y(
        \U_0/U_0/U_0/nfdata[5] ) );
  TBUFX1 \U_0/U_0/U_0/nfdata_tri[4]  ( .A(n6937), .EN(n6941), .Y(
        \U_0/U_0/U_0/nfdata[4] ) );
  TBUFX1 \U_0/U_0/U_0/nfdata_tri[3]  ( .A(n6936), .EN(n6941), .Y(
        \U_0/U_0/U_0/nfdata[3] ) );
  TBUFX1 \U_0/U_0/U_0/nfdata_tri[2]  ( .A(n6935), .EN(n6941), .Y(
        \U_0/U_0/U_0/nfdata[2] ) );
  TBUFX1 \U_0/U_0/U_0/nfdata_tri[1]  ( .A(n6934), .EN(n6941), .Y(
        \U_0/U_0/U_0/nfdata[1] ) );
  TBUFX1 \U_0/U_0/U_0/nfdata_tri[0]  ( .A(n6933), .EN(n6941), .Y(
        \U_0/U_0/U_0/nfdata[0] ) );
  TBUFX1 \U_1/U_0/U_0/nfaddr_tri[7]  ( .A(n6949), .EN(n9201), .Y(
        \U_1/U_0/U_0/nfaddr[7] ) );
  TBUFX1 \U_1/U_0/U_0/nfaddr_tri[6]  ( .A(n6948), .EN(n9201), .Y(
        \U_1/U_0/U_0/nfaddr[6] ) );
  TBUFX1 \U_1/U_0/U_0/nfaddr_tri[5]  ( .A(n6947), .EN(n9201), .Y(
        \U_1/U_0/U_0/nfaddr[5] ) );
  TBUFX1 \U_1/U_0/U_0/nfaddr_tri[4]  ( .A(n6946), .EN(n9201), .Y(
        \U_1/U_0/U_0/nfaddr[4] ) );
  TBUFX1 \U_1/U_0/U_0/nfaddr_tri[3]  ( .A(n6945), .EN(n9201), .Y(
        \U_1/U_0/U_0/nfaddr[3] ) );
  TBUFX1 \U_1/U_0/U_0/nfaddr_tri[2]  ( .A(n6944), .EN(n9201), .Y(
        \U_1/U_0/U_0/nfaddr[2] ) );
  TBUFX1 \U_1/U_0/U_0/nfaddr_tri[1]  ( .A(n6943), .EN(n9201), .Y(
        \U_1/U_0/U_0/nfaddr[1] ) );
  TBUFX1 \U_1/U_0/U_0/nfaddr_tri[0]  ( .A(n6942), .EN(n9201), .Y(
        \U_1/U_0/U_0/nfaddr[0] ) );
  TBUFX1 \U_0/U_0/U_0/nfaddr_tri[7]  ( .A(n6931), .EN(n11144), .Y(
        \U_0/U_0/U_0/nfaddr[7] ) );
  TBUFX1 \U_0/U_0/U_0/nfaddr_tri[6]  ( .A(n6930), .EN(n11144), .Y(
        \U_0/U_0/U_0/nfaddr[6] ) );
  TBUFX1 \U_0/U_0/U_0/nfaddr_tri[5]  ( .A(n6929), .EN(n11144), .Y(
        \U_0/U_0/U_0/nfaddr[5] ) );
  TBUFX1 \U_0/U_0/U_0/nfaddr_tri[4]  ( .A(n6928), .EN(n11144), .Y(
        \U_0/U_0/U_0/nfaddr[4] ) );
  TBUFX1 \U_0/U_0/U_0/nfaddr_tri[3]  ( .A(n6927), .EN(n11144), .Y(
        \U_0/U_0/U_0/nfaddr[3] ) );
  TBUFX1 \U_0/U_0/U_0/nfaddr_tri[2]  ( .A(n6926), .EN(n11144), .Y(
        \U_0/U_0/U_0/nfaddr[2] ) );
  TBUFX1 \U_0/U_0/U_0/nfaddr_tri[1]  ( .A(n6925), .EN(n11144), .Y(
        \U_0/U_0/U_0/nfaddr[1] ) );
  TBUFX1 \U_0/U_0/U_0/nfaddr_tri[0]  ( .A(n6924), .EN(n11144), .Y(
        \U_0/U_0/U_0/nfaddr[0] ) );
  TBUFX1 \U_1/U_0/U_0/nfdata_tri[7]  ( .A(n6958), .EN(n11913), .Y(
        \U_1/U_0/U_0/nfdata[7] ) );
  TBUFX1 \U_1/U_0/U_0/nfdata_tri[6]  ( .A(n6957), .EN(n11913), .Y(
        \U_1/U_0/U_0/nfdata[6] ) );
  TBUFX1 \U_1/U_0/U_0/nfdata_tri[5]  ( .A(n6956), .EN(n11913), .Y(
        \U_1/U_0/U_0/nfdata[5] ) );
  TBUFX1 \U_1/U_0/U_0/nfdata_tri[4]  ( .A(n6955), .EN(n11913), .Y(
        \U_1/U_0/U_0/nfdata[4] ) );
  TBUFX1 \U_1/U_0/U_0/nfdata_tri[3]  ( .A(n6954), .EN(n11913), .Y(
        \U_1/U_0/U_0/nfdata[3] ) );
  TBUFX1 \U_1/U_0/U_0/nfdata_tri[2]  ( .A(n6953), .EN(n11913), .Y(
        \U_1/U_0/U_0/nfdata[2] ) );
  TBUFX1 \U_1/U_0/U_0/nfdata_tri[1]  ( .A(n6952), .EN(n11913), .Y(
        \U_1/U_0/U_0/nfdata[1] ) );
  TBUFX1 \U_1/U_0/U_0/nfdata_tri[0]  ( .A(n6951), .EN(n11913), .Y(
        \U_1/U_0/U_0/nfdata[0] ) );
  AND2X2 U9188 ( .A(n9276), .B(n1020), .Y(n9163) );
  OR2X2 U9189 ( .A(n9409), .B(n10766), .Y(n9164) );
  OR2X2 U9190 ( .A(n9444), .B(n11518), .Y(n9165) );
  OR2X2 U9191 ( .A(n6661), .B(n6725), .Y(n9166) );
  OR2X2 U9192 ( .A(n1005), .B(n1006), .Y(n9167) );
  AND2X2 U9193 ( .A(n320), .B(n1016), .Y(n9168) );
  AND2X2 U9194 ( .A(n4788), .B(n4694), .Y(n9169) );
  AND2X2 U9195 ( .A(n2287), .B(n2193), .Y(n9170) );
  AND2X2 U9196 ( .A(n9193), .B(n9211), .Y(n9171) );
  AND2X2 U9197 ( .A(n9203), .B(n9249), .Y(n9172) );
  INVX2 U9198 ( .A(n9465), .Y(n9457) );
  INVX2 U9199 ( .A(n9466), .Y(n9456) );
  INVX2 U9200 ( .A(n9464), .Y(n9458) );
  INVX2 U9201 ( .A(n9462), .Y(n9460) );
  INVX2 U9202 ( .A(n9463), .Y(n9459) );
  INVX2 U9203 ( .A(n9428), .Y(n9421) );
  INVX2 U9204 ( .A(n9425), .Y(n9423) );
  INVX2 U9205 ( .A(n9426), .Y(n9422) );
  INVX2 U9206 ( .A(n9454), .Y(n9452) );
  INVX2 U9207 ( .A(n9419), .Y(n9417) );
  BUFX2 U9208 ( .A(n9173), .Y(n9453) );
  BUFX2 U9209 ( .A(n9174), .Y(n9418) );
  INVX2 U9210 ( .A(n9265), .Y(n10198) );
  INVX2 U9211 ( .A(n9266), .Y(n10199) );
  INVX2 U9212 ( .A(n9267), .Y(n10200) );
  INVX2 U9213 ( .A(n9252), .Y(n10121) );
  INVX2 U9214 ( .A(n9253), .Y(n10122) );
  INVX2 U9215 ( .A(n9254), .Y(n10123) );
  INVX2 U9216 ( .A(n9255), .Y(n10124) );
  INVX2 U9217 ( .A(n9272), .Y(n10237) );
  INVX2 U9218 ( .A(n9273), .Y(n10238) );
  INVX2 U9219 ( .A(n9274), .Y(n10239) );
  INVX2 U9220 ( .A(n9227), .Y(n9867) );
  INVX2 U9221 ( .A(n9228), .Y(n9868) );
  INVX2 U9222 ( .A(n9229), .Y(n9869) );
  INVX2 U9223 ( .A(n9214), .Y(n9790) );
  INVX2 U9224 ( .A(n9215), .Y(n9791) );
  INVX2 U9225 ( .A(n9216), .Y(n9792) );
  INVX2 U9226 ( .A(n9217), .Y(n9793) );
  INVX2 U9227 ( .A(n9234), .Y(n9906) );
  INVX2 U9228 ( .A(n9235), .Y(n9907) );
  INVX2 U9229 ( .A(n9236), .Y(n9908) );
  INVX2 U9230 ( .A(n9264), .Y(n10197) );
  INVX2 U9231 ( .A(n9226), .Y(n9866) );
  INVX2 U9232 ( .A(n9260), .Y(n10169) );
  INVX2 U9233 ( .A(n9261), .Y(n10178) );
  INVX2 U9234 ( .A(n9262), .Y(n10187) );
  INVX2 U9235 ( .A(n9263), .Y(n10196) );
  INVX2 U9236 ( .A(n9268), .Y(n10209) );
  INVX2 U9237 ( .A(n9269), .Y(n10218) );
  INVX2 U9238 ( .A(n9257), .Y(n10142) );
  INVX2 U9239 ( .A(n9258), .Y(n10151) );
  INVX2 U9240 ( .A(n9259), .Y(n10160) );
  INVX2 U9241 ( .A(n9270), .Y(n10227) );
  INVX2 U9242 ( .A(n9271), .Y(n10236) );
  INVX2 U9243 ( .A(n9222), .Y(n9838) );
  INVX2 U9244 ( .A(n9223), .Y(n9847) );
  INVX2 U9245 ( .A(n9224), .Y(n9856) );
  INVX2 U9246 ( .A(n9225), .Y(n9865) );
  INVX2 U9247 ( .A(n9230), .Y(n9878) );
  INVX2 U9248 ( .A(n9231), .Y(n9887) );
  INVX2 U9249 ( .A(n9219), .Y(n9811) );
  INVX2 U9250 ( .A(n9220), .Y(n9820) );
  INVX2 U9251 ( .A(n9221), .Y(n9829) );
  INVX2 U9252 ( .A(n9232), .Y(n9896) );
  INVX2 U9253 ( .A(n9233), .Y(n9905) );
  INVX2 U9254 ( .A(n9256), .Y(n10133) );
  INVX2 U9255 ( .A(n9218), .Y(n9802) );
  INVX2 U9256 ( .A(n1714), .Y(n10241) );
  INVX2 U9257 ( .A(n1712), .Y(n10242) );
  INVX2 U9258 ( .A(n1710), .Y(n10243) );
  INVX2 U9259 ( .A(n1700), .Y(n10244) );
  INVX2 U9260 ( .A(n4217), .Y(n9910) );
  INVX2 U9261 ( .A(n4215), .Y(n9911) );
  INVX2 U9262 ( .A(n4213), .Y(n9912) );
  INVX2 U9263 ( .A(n4203), .Y(n9913) );
  INVX2 U9264 ( .A(n1682), .Y(n10262) );
  INVX2 U9265 ( .A(n1672), .Y(n10271) );
  INVX2 U9266 ( .A(n4185), .Y(n9931) );
  INVX2 U9267 ( .A(n4175), .Y(n9940) );
  INVX2 U9268 ( .A(n1662), .Y(n10280) );
  INVX2 U9269 ( .A(n4165), .Y(n9949) );
  INVX2 U9270 ( .A(n1692), .Y(n10253) );
  INVX2 U9271 ( .A(n4195), .Y(n9922) );
  BUFX2 U9272 ( .A(n9163), .Y(n9466) );
  BUFX2 U9273 ( .A(n9163), .Y(n9465) );
  BUFX2 U9274 ( .A(n9163), .Y(n9464) );
  BUFX2 U9275 ( .A(n9163), .Y(n9463) );
  BUFX2 U9276 ( .A(n9163), .Y(n9462) );
  BUFX2 U9277 ( .A(n9467), .Y(n9461) );
  BUFX2 U9278 ( .A(n9465), .Y(n9472) );
  BUFX2 U9279 ( .A(n9464), .Y(n9471) );
  BUFX2 U9280 ( .A(n9466), .Y(n9470) );
  BUFX2 U9281 ( .A(n9163), .Y(n9469) );
  BUFX2 U9282 ( .A(n9163), .Y(n9467) );
  BUFX2 U9283 ( .A(n9163), .Y(n9468) );
  INVX2 U9284 ( .A(n9442), .Y(n9443) );
  INVX2 U9285 ( .A(n9407), .Y(n9408) );
  INVX2 U9286 ( .A(n9444), .Y(n9446) );
  INVX2 U9287 ( .A(n9409), .Y(n9411) );
  BUFX2 U9288 ( .A(n9437), .Y(n9429) );
  BUFX2 U9289 ( .A(n9437), .Y(n9428) );
  BUFX2 U9290 ( .A(n9437), .Y(n9427) );
  BUFX2 U9291 ( .A(n9437), .Y(n9426) );
  BUFX2 U9292 ( .A(n9437), .Y(n9425) );
  BUFX2 U9293 ( .A(n9437), .Y(n9424) );
  BUFX2 U9294 ( .A(n9437), .Y(n9435) );
  BUFX2 U9295 ( .A(n9437), .Y(n9434) );
  BUFX2 U9296 ( .A(n9437), .Y(n9433) );
  BUFX2 U9297 ( .A(n9437), .Y(n9432) );
  BUFX2 U9298 ( .A(n9437), .Y(n9430) );
  BUFX2 U9299 ( .A(n9437), .Y(n9431) );
  INVX2 U9300 ( .A(n9444), .Y(n9445) );
  INVX2 U9301 ( .A(n9409), .Y(n9410) );
  BUFX2 U9302 ( .A(n9468), .Y(n9473) );
  BUFX2 U9303 ( .A(n9424), .Y(n9436) );
  BUFX2 U9304 ( .A(n9173), .Y(n9454) );
  BUFX2 U9305 ( .A(n9174), .Y(n9419) );
  INVX2 U9306 ( .A(n9175), .Y(n9284) );
  INVX2 U9307 ( .A(n9176), .Y(n9242) );
  BUFX2 U9308 ( .A(n9173), .Y(n9455) );
  BUFX2 U9309 ( .A(n9174), .Y(n9420) );
  OR2X2 U9310 ( .A(n2034), .B(n9180), .Y(n9173) );
  OR2X2 U9311 ( .A(n4535), .B(n9181), .Y(n9174) );
  BUFX2 U9312 ( .A(n1806), .Y(n9260) );
  BUFX2 U9313 ( .A(n1796), .Y(n9261) );
  BUFX2 U9314 ( .A(n1786), .Y(n9262) );
  BUFX2 U9315 ( .A(n1776), .Y(n9263) );
  BUFX2 U9316 ( .A(n1758), .Y(n9268) );
  BUFX2 U9317 ( .A(n1748), .Y(n9269) );
  BUFX2 U9318 ( .A(n1846), .Y(n9256) );
  BUFX2 U9319 ( .A(n1836), .Y(n9257) );
  BUFX2 U9320 ( .A(n1826), .Y(n9258) );
  BUFX2 U9321 ( .A(n1816), .Y(n9259) );
  BUFX2 U9322 ( .A(n1738), .Y(n9270) );
  BUFX2 U9323 ( .A(n1728), .Y(n9271) );
  BUFX2 U9324 ( .A(n4309), .Y(n9222) );
  BUFX2 U9325 ( .A(n4299), .Y(n9223) );
  BUFX2 U9326 ( .A(n4289), .Y(n9224) );
  BUFX2 U9327 ( .A(n4279), .Y(n9225) );
  BUFX2 U9328 ( .A(n4261), .Y(n9230) );
  BUFX2 U9329 ( .A(n4251), .Y(n9231) );
  BUFX2 U9330 ( .A(n4349), .Y(n9218) );
  BUFX2 U9331 ( .A(n4339), .Y(n9219) );
  BUFX2 U9332 ( .A(n4329), .Y(n9220) );
  BUFX2 U9333 ( .A(n4319), .Y(n9221) );
  BUFX2 U9334 ( .A(n4241), .Y(n9232) );
  BUFX2 U9335 ( .A(n4231), .Y(n9233) );
  BUFX2 U9336 ( .A(n1772), .Y(n9264) );
  BUFX2 U9337 ( .A(n1770), .Y(n9265) );
  BUFX2 U9338 ( .A(n1768), .Y(n9266) );
  BUFX2 U9339 ( .A(n1766), .Y(n9267) );
  BUFX2 U9340 ( .A(n1860), .Y(n9252) );
  BUFX2 U9341 ( .A(n1858), .Y(n9253) );
  BUFX2 U9342 ( .A(n1856), .Y(n9254) );
  BUFX2 U9343 ( .A(n1854), .Y(n9255) );
  BUFX2 U9344 ( .A(n1720), .Y(n9272) );
  BUFX2 U9345 ( .A(n1718), .Y(n9273) );
  BUFX2 U9346 ( .A(n1716), .Y(n9274) );
  BUFX2 U9347 ( .A(n4275), .Y(n9226) );
  BUFX2 U9348 ( .A(n4273), .Y(n9227) );
  BUFX2 U9349 ( .A(n4271), .Y(n9228) );
  BUFX2 U9350 ( .A(n4269), .Y(n9229) );
  BUFX2 U9351 ( .A(n4363), .Y(n9214) );
  BUFX2 U9352 ( .A(n4361), .Y(n9215) );
  BUFX2 U9353 ( .A(n4359), .Y(n9216) );
  BUFX2 U9354 ( .A(n4357), .Y(n9217) );
  BUFX2 U9355 ( .A(n4223), .Y(n9234) );
  BUFX2 U9356 ( .A(n4221), .Y(n9235) );
  BUFX2 U9357 ( .A(n4219), .Y(n9236) );
  BUFX2 U9358 ( .A(n1722), .Y(n9275) );
  BUFX2 U9359 ( .A(n4225), .Y(n9237) );
  BUFX2 U9360 ( .A(n10055), .Y(n9369) );
  BUFX2 U9361 ( .A(n9724), .Y(n9359) );
  BUFX2 U9362 ( .A(n10055), .Y(n9365) );
  BUFX2 U9363 ( .A(n9724), .Y(n9355) );
  BUFX2 U9364 ( .A(n10055), .Y(n9366) );
  BUFX2 U9365 ( .A(n10055), .Y(n9367) );
  BUFX2 U9366 ( .A(n10055), .Y(n9368) );
  BUFX2 U9367 ( .A(n9724), .Y(n9356) );
  BUFX2 U9368 ( .A(n9724), .Y(n9357) );
  BUFX2 U9369 ( .A(n9724), .Y(n9358) );
  BUFX2 U9370 ( .A(n9184), .Y(n9376) );
  BUFX2 U9371 ( .A(n9185), .Y(n9380) );
  BUFX2 U9372 ( .A(n9184), .Y(n9377) );
  BUFX2 U9373 ( .A(n9185), .Y(n9381) );
  BUFX2 U9374 ( .A(n9184), .Y(n9375) );
  BUFX2 U9375 ( .A(n9185), .Y(n9379) );
  INVX2 U9376 ( .A(n6170), .Y(n11914) );
  INVX2 U9377 ( .A(n3434), .Y(n10012) );
  INVX2 U9378 ( .A(n3473), .Y(n11134) );
  INVX2 U9379 ( .A(n9165), .Y(n9440) );
  INVX2 U9380 ( .A(n9165), .Y(n9439) );
  INVX2 U9381 ( .A(n9164), .Y(n9405) );
  INVX2 U9382 ( .A(n9164), .Y(n9404) );
  INVX2 U9383 ( .A(n9165), .Y(n9438) );
  INVX2 U9384 ( .A(n9164), .Y(n9403) );
  BUFX2 U9385 ( .A(n9184), .Y(n9378) );
  BUFX2 U9386 ( .A(n9185), .Y(n9382) );
  INVX2 U9387 ( .A(n9177), .Y(n9249) );
  INVX2 U9388 ( .A(n9178), .Y(n9211) );
  INVX2 U9389 ( .A(n3589), .Y(n9437) );
  INVX2 U9390 ( .A(n6188), .Y(n11896) );
  INVX2 U9391 ( .A(n3570), .Y(n11155) );
  INVX2 U9392 ( .A(n9179), .Y(n9197) );
  AND2X2 U9393 ( .A(n11642), .B(n9283), .Y(n9175) );
  INVX2 U9394 ( .A(n321), .Y(n11899) );
  INVX2 U9395 ( .A(n2237), .Y(n11467) );
  INVX2 U9396 ( .A(n4738), .Y(n10715) );
  AND2X2 U9397 ( .A(n10891), .B(n9241), .Y(n9176) );
  INVX2 U9398 ( .A(n9204), .Y(n11557) );
  INVX2 U9399 ( .A(n9194), .Y(n10805) );
  INVX2 U9400 ( .A(n9180), .Y(n9248) );
  INVX2 U9401 ( .A(n9181), .Y(n9210) );
  BUFX2 U9402 ( .A(n10056), .Y(n9370) );
  BUFX2 U9403 ( .A(n10056), .Y(n9371) );
  BUFX2 U9404 ( .A(n10056), .Y(n9372) );
  BUFX2 U9405 ( .A(n10056), .Y(n9373) );
  BUFX2 U9406 ( .A(n9725), .Y(n9360) );
  BUFX2 U9407 ( .A(n9725), .Y(n9361) );
  BUFX2 U9408 ( .A(n9725), .Y(n9362) );
  BUFX2 U9409 ( .A(n9725), .Y(n9363) );
  INVX2 U9410 ( .A(n6204), .Y(n11886) );
  INVX2 U9411 ( .A(n9442), .Y(n9441) );
  INVX2 U9412 ( .A(n2200), .Y(n9442) );
  INVX2 U9413 ( .A(n9407), .Y(n9406) );
  INVX2 U9414 ( .A(n4701), .Y(n9407) );
  INVX2 U9415 ( .A(n2177), .Y(n9444) );
  INVX2 U9416 ( .A(n4678), .Y(n9409) );
  BUFX2 U9417 ( .A(n2170), .Y(n9447) );
  BUFX2 U9418 ( .A(n4671), .Y(n9412) );
  BUFX2 U9419 ( .A(n2170), .Y(n9448) );
  BUFX2 U9420 ( .A(n2170), .Y(n9449) );
  BUFX2 U9421 ( .A(n2170), .Y(n9450) );
  BUFX2 U9422 ( .A(n4671), .Y(n9413) );
  BUFX2 U9423 ( .A(n4671), .Y(n9414) );
  BUFX2 U9424 ( .A(n4671), .Y(n9415) );
  BUFX2 U9425 ( .A(n2170), .Y(n9451) );
  BUFX2 U9426 ( .A(n4671), .Y(n9416) );
  INVX2 U9427 ( .A(n304), .Y(n11918) );
  INVX2 U9428 ( .A(n308), .Y(n11892) );
  BUFX2 U9429 ( .A(n6631), .Y(n9188) );
  BUFX2 U9430 ( .A(n6807), .Y(n9191) );
  AND2X2 U9431 ( .A(n9205), .B(n9180), .Y(n9177) );
  AND2X2 U9432 ( .A(n9195), .B(n9181), .Y(n9178) );
  BUFX2 U9433 ( .A(n10056), .Y(n9374) );
  BUFX2 U9434 ( .A(n9725), .Y(n9364) );
  INVX2 U9435 ( .A(n6110), .Y(n9198) );
  INVX2 U9436 ( .A(n9167), .Y(n9280) );
  INVX2 U9437 ( .A(n3574), .Y(n9238) );
  INVX2 U9438 ( .A(n1056), .Y(n9278) );
  INVX2 U9439 ( .A(n9182), .Y(n9247) );
  INVX2 U9440 ( .A(n9183), .Y(n9209) );
  INVX4 U9441 ( .A(n9476), .Y(n9474) );
  INVX4 U9442 ( .A(n9483), .Y(n9481) );
  INVX2 U9443 ( .A(n6205), .Y(n11913) );
  INVX2 U9444 ( .A(n3444), .Y(n11144) );
  INVX2 U9445 ( .A(n951), .Y(n11883) );
  BUFX2 U9446 ( .A(n792), .Y(n9285) );
  BUFX2 U9447 ( .A(n3314), .Y(n9243) );
  OR2X2 U9448 ( .A(n6165), .B(n11928), .Y(n9179) );
  INVX2 U9449 ( .A(n9172), .Y(n9250) );
  INVX2 U9450 ( .A(n9171), .Y(n9212) );
  INVX2 U9451 ( .A(n9168), .Y(n9199) );
  INVX2 U9452 ( .A(n2316), .Y(n11393) );
  INVX2 U9453 ( .A(n4817), .Y(n10641) );
  INVX2 U9454 ( .A(n9282), .Y(n9283) );
  INVX2 U9455 ( .A(n9240), .Y(n9241) );
  INVX2 U9456 ( .A(n9170), .Y(n9246) );
  INVX2 U9457 ( .A(n9169), .Y(n9208) );
  BUFX2 U9458 ( .A(n1888), .Y(n9204) );
  BUFX2 U9459 ( .A(n4391), .Y(n9194) );
  OR2X2 U9460 ( .A(n11547), .B(n11557), .Y(n9180) );
  OR2X2 U9461 ( .A(n10795), .B(n10805), .Y(n9181) );
  BUFX2 U9462 ( .A(n3144), .Y(n9245) );
  BUFX2 U9463 ( .A(n5645), .Y(n9207) );
  BUFX2 U9464 ( .A(n893), .Y(n9276) );
  INVX2 U9465 ( .A(n9308), .Y(n9309) );
  INVX2 U9466 ( .A(n9310), .Y(n9311) );
  INVX2 U9467 ( .A(n9302), .Y(n9303) );
  INVX2 U9468 ( .A(n9343), .Y(n9344) );
  INVX2 U9469 ( .A(n9345), .Y(n9346) );
  INVX2 U9470 ( .A(n9337), .Y(n9338) );
  INVX2 U9471 ( .A(n9314), .Y(n9315) );
  INVX2 U9472 ( .A(n9349), .Y(n9350) );
  INVX2 U9473 ( .A(n9312), .Y(n9313) );
  INVX2 U9474 ( .A(n9304), .Y(n9305) );
  INVX2 U9475 ( .A(n9347), .Y(n9348) );
  INVX2 U9476 ( .A(n9339), .Y(n9340) );
  INVX2 U9477 ( .A(n9306), .Y(n9307) );
  INVX2 U9478 ( .A(n9341), .Y(n9342) );
  INVX2 U9479 ( .A(n9316), .Y(n9317) );
  INVX2 U9480 ( .A(n9351), .Y(n9352) );
  INVX4 U9481 ( .A(n9480), .Y(n9479) );
  INVX4 U9482 ( .A(n9487), .Y(n9486) );
  BUFX2 U9483 ( .A(n1065), .Y(n9277) );
  BUFX2 U9484 ( .A(n1034), .Y(n9279) );
  OR2X2 U9485 ( .A(n2161), .B(n2155), .Y(n9182) );
  OR2X2 U9486 ( .A(n4662), .B(n4656), .Y(n9183) );
  INVX2 U9487 ( .A(n6670), .Y(n9189) );
  INVX2 U9488 ( .A(n9166), .Y(n9187) );
  INVX2 U9489 ( .A(n9184), .Y(n9251) );
  INVX2 U9490 ( .A(n9185), .Y(n9213) );
  INVX2 U9491 ( .A(n9293), .Y(n9294) );
  INVX2 U9492 ( .A(n9327), .Y(n9328) );
  INVX2 U9493 ( .A(n9287), .Y(n9288) );
  INVX2 U9494 ( .A(n9321), .Y(n9322) );
  BUFX2 U9495 ( .A(n9478), .Y(n9476) );
  BUFX2 U9496 ( .A(n9485), .Y(n9483) );
  BUFX2 U9497 ( .A(n1888), .Y(n9205) );
  BUFX2 U9498 ( .A(n4391), .Y(n9195) );
  INVX2 U9499 ( .A(n956), .Y(n9200) );
  INVX2 U9500 ( .A(n6672), .Y(n9190) );
  INVX2 U9501 ( .A(n819), .Y(n9282) );
  INVX2 U9502 ( .A(n3341), .Y(n9240) );
  INVX2 U9503 ( .A(n1659), .Y(n10282) );
  INVX2 U9504 ( .A(n4162), .Y(n9951) );
  BUFX2 U9505 ( .A(n11520), .Y(n9393) );
  BUFX2 U9506 ( .A(n10768), .Y(n9383) );
  BUFX2 U9507 ( .A(n11520), .Y(n9394) );
  BUFX2 U9508 ( .A(n11520), .Y(n9395) );
  BUFX2 U9509 ( .A(n11520), .Y(n9396) );
  BUFX2 U9510 ( .A(n10768), .Y(n9384) );
  BUFX2 U9511 ( .A(n10768), .Y(n9385) );
  BUFX2 U9512 ( .A(n10768), .Y(n9386) );
  BUFX2 U9513 ( .A(n11523), .Y(n9398) );
  BUFX2 U9514 ( .A(n10771), .Y(n9388) );
  BUFX2 U9515 ( .A(n11523), .Y(n9399) );
  BUFX2 U9516 ( .A(n11523), .Y(n9400) );
  BUFX2 U9517 ( .A(n11523), .Y(n9401) );
  BUFX2 U9518 ( .A(n10771), .Y(n9389) );
  BUFX2 U9519 ( .A(n10771), .Y(n9390) );
  BUFX2 U9520 ( .A(n10771), .Y(n9391) );
  INVX2 U9521 ( .A(n2212), .Y(n11410) );
  INVX2 U9522 ( .A(n4713), .Y(n10658) );
  INVX2 U9523 ( .A(n2302), .Y(n11445) );
  INVX2 U9524 ( .A(n2247), .Y(n11427) );
  INVX2 U9525 ( .A(n4803), .Y(n10693) );
  INVX2 U9526 ( .A(n4748), .Y(n10675) );
  INVX2 U9527 ( .A(n2197), .Y(n11461) );
  INVX2 U9528 ( .A(n4698), .Y(n10709) );
  INVX2 U9529 ( .A(n2266), .Y(n11496) );
  INVX2 U9530 ( .A(n2232), .Y(n11478) );
  INVX2 U9531 ( .A(n4767), .Y(n10744) );
  INVX2 U9532 ( .A(n4733), .Y(n10726) );
  INVX2 U9533 ( .A(n2286), .Y(n11374) );
  INVX2 U9534 ( .A(n4787), .Y(n10622) );
  BUFX2 U9535 ( .A(n11523), .Y(n9402) );
  BUFX2 U9536 ( .A(n10771), .Y(n9392) );
  BUFX2 U9537 ( .A(n776), .Y(n9239) );
  BUFX2 U9538 ( .A(n11520), .Y(n9397) );
  BUFX2 U9539 ( .A(n10768), .Y(n9387) );
  INVX2 U9540 ( .A(n9291), .Y(n9292) );
  INVX2 U9541 ( .A(n9325), .Y(n9326) );
  INVX2 U9542 ( .A(n9289), .Y(n9290) );
  INVX2 U9543 ( .A(n9323), .Y(n9324) );
  INVX2 U9544 ( .A(n9186), .Y(n9201) );
  BUFX2 U9545 ( .A(n1888), .Y(n9203) );
  BUFX2 U9546 ( .A(n4391), .Y(n9193) );
  BUFX2 U9547 ( .A(n9478), .Y(n9475) );
  BUFX2 U9548 ( .A(n9485), .Y(n9482) );
  INVX2 U9549 ( .A(n238), .Y(n10509) );
  INVX2 U9550 ( .A(n523), .Y(n10510) );
  BUFX2 U9551 ( .A(n9478), .Y(n9477) );
  BUFX2 U9552 ( .A(n9485), .Y(n9484) );
  INVX2 U9553 ( .A(n9202), .Y(n9698) );
  INVX2 U9554 ( .A(n9192), .Y(n9690) );
  INVX2 U9555 ( .A(\U_1/U_2/U_5/state[1] ), .Y(n11577) );
  INVX2 U9556 ( .A(\U_0/U_2/U_5/state[1] ), .Y(n10825) );
  INVX2 U9557 ( .A(\U_1/U_1/U_1/writeptr[1] ), .Y(n9289) );
  INVX2 U9558 ( .A(\U_0/U_1/U_1/writeptr[1] ), .Y(n9323) );
  INVX2 U9559 ( .A(\U_1/RCV_DATA [3]), .Y(n9308) );
  INVX2 U9560 ( .A(\U_1/RCV_DATA [4]), .Y(n9310) );
  INVX2 U9561 ( .A(\U_1/RCV_DATA [6]), .Y(n9314) );
  INVX2 U9562 ( .A(\U_1/RCV_DATA [5]), .Y(n9312) );
  INVX2 U9563 ( .A(\U_1/RCV_DATA [0]), .Y(n9302) );
  INVX2 U9564 ( .A(\U_1/RCV_DATA [2]), .Y(n9306) );
  INVX2 U9565 ( .A(\U_1/RCV_DATA [1]), .Y(n9304) );
  INVX2 U9566 ( .A(\U_0/RCV_DATA [3]), .Y(n9343) );
  INVX2 U9567 ( .A(\U_0/RCV_DATA [4]), .Y(n9345) );
  INVX2 U9568 ( .A(\U_0/RCV_DATA [6]), .Y(n9349) );
  INVX2 U9569 ( .A(\U_0/RCV_DATA [5]), .Y(n9347) );
  INVX2 U9570 ( .A(\U_0/RCV_DATA [0]), .Y(n9337) );
  INVX2 U9571 ( .A(\U_0/RCV_DATA [2]), .Y(n9341) );
  INVX2 U9572 ( .A(\U_0/RCV_DATA [1]), .Y(n9339) );
  INVX2 U9573 ( .A(\U_1/RCV_DATA [7]), .Y(n9316) );
  INVX2 U9574 ( .A(\U_0/RCV_DATA [7]), .Y(n9351) );
  INVX2 U9575 ( .A(\U_1/U_2/U_5/state[2] ), .Y(n9301) );
  INVX2 U9576 ( .A(\U_0/U_2/U_5/state[2] ), .Y(n9336) );
  BUFX2 U9577 ( .A(\U_0/U_0/U_0/state[4] ), .Y(n9320) );
  INVX2 U9578 ( .A(\U_1/U_0/U_1/RCV_DATA [0]), .Y(n9480) );
  INVX2 U9579 ( .A(\U_0/U_0/U_1/RCV_DATA [0]), .Y(n9487) );
  BUFX2 U9580 ( .A(n6105), .Y(n9196) );
  OR2X2 U9581 ( .A(n9249), .B(RST), .Y(n9184) );
  OR2X2 U9582 ( .A(n9211), .B(RST), .Y(n9185) );
  BUFX2 U9583 ( .A(\U_1/U_0/U_0/state[4] ), .Y(n9286) );
  INVX2 U9584 ( .A(\U_1/U_1/U_1/writeptr[2] ), .Y(n9287) );
  INVX2 U9585 ( .A(\U_0/U_1/U_1/writeptr[2] ), .Y(n9321) );
  INVX2 U9586 ( .A(\U_1/U_1/U_1/writeptr[3] ), .Y(n9291) );
  INVX2 U9587 ( .A(\U_1/U_1/U_1/writeptr[4] ), .Y(n9293) );
  INVX2 U9588 ( .A(\U_0/U_1/U_1/writeptr[3] ), .Y(n9325) );
  INVX2 U9589 ( .A(\U_0/U_1/U_1/writeptr[4] ), .Y(n9327) );
  INVX2 U9590 ( .A(\U_1/U_1/U_1/readptr[1] ), .Y(n9299) );
  INVX2 U9591 ( .A(\U_0/U_1/U_1/readptr[1] ), .Y(n9333) );
  INVX2 U9592 ( .A(\U_1/U_1/U_1/readptr[0] ), .Y(n9300) );
  INVX2 U9593 ( .A(\U_0/U_1/U_1/readptr[0] ), .Y(n9334) );
  INVX2 U9594 ( .A(\U_1/U_1/U_1/readptr[2] ), .Y(n9298) );
  INVX2 U9595 ( .A(\U_0/U_1/U_1/readptr[2] ), .Y(n9332) );
  INVX2 U9596 ( .A(n9296), .Y(n9297) );
  INVX2 U9597 ( .A(\U_1/U_1/U_1/readptr[3] ), .Y(n9296) );
  INVX2 U9598 ( .A(n9330), .Y(n9331) );
  INVX2 U9599 ( .A(\U_0/U_1/U_1/readptr[3] ), .Y(n9330) );
  INVX2 U9600 ( .A(\U_1/U_1/U_1/readptr[4] ), .Y(n9295) );
  INVX2 U9601 ( .A(\U_0/U_1/U_1/readptr[4] ), .Y(n9329) );
  INVX2 U9602 ( .A(\U_0/U_3/U_3/N188 ), .Y(n9335) );
  INVX2 U9603 ( .A(\U_1/U_0/U_1/RCV_DATA [2]), .Y(n9478) );
  INVX2 U9604 ( .A(\U_0/U_0/U_1/RCV_DATA [2]), .Y(n9485) );
  INVX2 U9605 ( .A(\U_1/U_0/U_1/U_8/address[3] ), .Y(n11508) );
  INVX2 U9606 ( .A(\U_0/U_0/U_1/U_8/address[3] ), .Y(n10756) );
  OR2X2 U9607 ( .A(n1004), .B(n6150), .Y(n9186) );
  INVX2 U9608 ( .A(n777), .Y(n9281) );
  BUFX2 U9609 ( .A(\U_1/U_1/U_1/state ), .Y(n9318) );
  BUFX2 U9610 ( .A(\U_0/U_1/U_1/state ), .Y(n9353) );
  INVX2 U9611 ( .A(n5665), .Y(n9206) );
  INVX2 U9612 ( .A(n3164), .Y(n9244) );
  INVX2 U9613 ( .A(\U_1/U_0/U_1/RBUF_LOAD ), .Y(n9319) );
  INVX2 U9614 ( .A(\U_0/U_0/U_1/RBUF_LOAD ), .Y(n9354) );
  BUFX2 U9615 ( .A(n2159), .Y(n9202) );
  BUFX2 U9616 ( .A(n4660), .Y(n9192) );
  INVX2 U9617 ( .A(RST), .Y(n9527) );
  INVX2 U9618 ( .A(RST), .Y(n9526) );
  INVX2 U9619 ( .A(RST), .Y(n9524) );
  INVX2 U9620 ( .A(RST), .Y(n9523) );
  INVX2 U9621 ( .A(RST), .Y(n9525) );
  INVX2 U9622 ( .A(RST), .Y(n9530) );
  INVX2 U9623 ( .A(RST), .Y(n9529) );
  INVX2 U9624 ( .A(RST), .Y(n9528) );
  INVX2 U9625 ( .A(RST), .Y(n9534) );
  INVX2 U9626 ( .A(RST), .Y(n9531) );
  INVX2 U9627 ( .A(RST), .Y(n9522) );
  INVX2 U9628 ( .A(RST), .Y(n9532) );
  INVX2 U9629 ( .A(RST), .Y(n9533) );
  INVX2 U9630 ( .A(RST), .Y(n9488) );
  INVX2 U9631 ( .A(RST), .Y(n9489) );
  INVX2 U9632 ( .A(RST), .Y(n9490) );
  INVX2 U9633 ( .A(RST), .Y(n9491) );
  INVX2 U9634 ( .A(RST), .Y(n9492) );
  INVX2 U9635 ( .A(RST), .Y(n9493) );
  INVX2 U9636 ( .A(RST), .Y(n9494) );
  INVX2 U9637 ( .A(RST), .Y(n9495) );
  INVX2 U9638 ( .A(RST), .Y(n9496) );
  INVX2 U9639 ( .A(RST), .Y(n9497) );
  INVX2 U9640 ( .A(RST), .Y(n9498) );
  INVX2 U9641 ( .A(RST), .Y(n9499) );
  INVX2 U9642 ( .A(RST), .Y(n9500) );
  INVX2 U9643 ( .A(RST), .Y(n9501) );
  INVX2 U9644 ( .A(RST), .Y(n9502) );
  INVX2 U9645 ( .A(RST), .Y(n9503) );
  INVX2 U9646 ( .A(RST), .Y(n9504) );
  INVX2 U9647 ( .A(RST), .Y(n9505) );
  INVX2 U9648 ( .A(RST), .Y(n9506) );
  INVX2 U9649 ( .A(RST), .Y(n9507) );
  INVX2 U9650 ( .A(RST), .Y(n9508) );
  INVX2 U9651 ( .A(RST), .Y(n9509) );
  INVX2 U9652 ( .A(RST), .Y(n9510) );
  INVX2 U9653 ( .A(RST), .Y(n9511) );
  INVX2 U9654 ( .A(RST), .Y(n9512) );
  INVX2 U9655 ( .A(RST), .Y(n9513) );
  INVX2 U9656 ( .A(RST), .Y(n9514) );
  INVX2 U9657 ( .A(RST), .Y(n9515) );
  INVX2 U9658 ( .A(RST), .Y(n9516) );
  INVX2 U9659 ( .A(RST), .Y(n9517) );
  INVX2 U9660 ( .A(RST), .Y(n9518) );
  INVX2 U9661 ( .A(RST), .Y(n9519) );
  INVX2 U9662 ( .A(RST), .Y(n9520) );
  INVX2 U9663 ( .A(RST), .Y(n9521) );
  OR2X1 U9664 ( .A(n9300), .B(\U_1/U_1/U_1/writeptr[0] ), .Y(
        \U_1/U_1/U_1/sub_72/carry[1] ) );
  XNOR2X1 U9665 ( .A(\U_1/U_1/U_1/writeptr[0] ), .B(n9300), .Y(
        \U_1/U_1/U_1/N189 ) );
  XOR2X1 U9666 ( .A(\U_1/U_1/U_1/readptr[4] ), .B(
        \U_1/U_1/U_1/add_76_aco/carry[4] ), .Y(\U_1/U_1/U_1/N337 ) );
  AND2X1 U9667 ( .A(n9297), .B(\U_1/U_1/U_1/add_76_aco/carry[3] ), .Y(
        \U_1/U_1/U_1/add_76_aco/carry[4] ) );
  XOR2X1 U9668 ( .A(\U_1/U_1/U_1/add_76_aco/carry[3] ), .B(n9297), .Y(
        \U_1/U_1/U_1/N336 ) );
  AND2X1 U9669 ( .A(\U_1/U_1/U_1/readptr[2] ), .B(
        \U_1/U_1/U_1/add_76_aco/carry[2] ), .Y(
        \U_1/U_1/U_1/add_76_aco/carry[3] ) );
  XOR2X1 U9670 ( .A(\U_1/U_1/U_1/add_76_aco/carry[2] ), .B(
        \U_1/U_1/U_1/readptr[2] ), .Y(\U_1/U_1/U_1/N335 ) );
  AND2X1 U9671 ( .A(\U_1/U_1/U_1/readptr[1] ), .B(
        \U_1/U_1/U_1/add_76_aco/carry[1] ), .Y(
        \U_1/U_1/U_1/add_76_aco/carry[2] ) );
  XOR2X1 U9672 ( .A(\U_1/U_1/U_1/add_76_aco/carry[1] ), .B(
        \U_1/U_1/U_1/readptr[1] ), .Y(\U_1/U_1/U_1/N334 ) );
  AND2X1 U9673 ( .A(\U_1/U_1/U_1/readptr[0] ), .B(\U_1/U_1/U_1/N195 ), .Y(
        \U_1/U_1/U_1/add_76_aco/carry[1] ) );
  XOR2X1 U9674 ( .A(\U_1/U_1/U_1/N195 ), .B(\U_1/U_1/U_1/readptr[0] ), .Y(
        \U_1/U_1/U_1/N333 ) );
  XOR2X1 U9675 ( .A(\U_1/U_3/U_3/N188 ), .B(\r2042/carry[6] ), .Y(
        \U_1/U_3/U_3/N90 ) );
  AND2X1 U9676 ( .A(\U_1/U_3/U_3/count[5] ), .B(\r2042/carry[5] ), .Y(
        \r2042/carry[6] ) );
  XOR2X1 U9677 ( .A(\r2042/carry[5] ), .B(\U_1/U_3/U_3/count[5] ), .Y(
        \U_1/U_3/U_3/N89 ) );
  AND2X1 U9678 ( .A(\U_1/U_3/U_3/count[4] ), .B(\r2042/carry[4] ), .Y(
        \r2042/carry[5] ) );
  XOR2X1 U9679 ( .A(\r2042/carry[4] ), .B(\U_1/U_3/U_3/count[4] ), .Y(
        \U_1/U_3/U_3/N88 ) );
  AND2X1 U9680 ( .A(\U_1/U_3/U_3/count[3] ), .B(\r2042/carry[3] ), .Y(
        \r2042/carry[4] ) );
  XOR2X1 U9681 ( .A(\r2042/carry[3] ), .B(\U_1/U_3/U_3/count[3] ), .Y(
        \U_1/U_3/U_3/N87 ) );
  AND2X1 U9682 ( .A(\U_1/U_3/U_3/count[2] ), .B(\r2042/carry[2] ), .Y(
        \r2042/carry[3] ) );
  XOR2X1 U9683 ( .A(\r2042/carry[2] ), .B(\U_1/U_3/U_3/count[2] ), .Y(
        \U_1/U_3/U_3/N86 ) );
  AND2X1 U9684 ( .A(\U_1/U_3/U_3/count[1] ), .B(\r2042/carry[1] ), .Y(
        \r2042/carry[2] ) );
  XOR2X1 U9685 ( .A(\r2042/carry[1] ), .B(\U_1/U_3/U_3/count[1] ), .Y(
        \U_1/U_3/U_3/N85 ) );
  AND2X1 U9686 ( .A(\U_1/U_3/U_3/count[0] ), .B(\U_1/U_3/U_0/N59 ), .Y(
        \r2042/carry[1] ) );
  XOR2X1 U9687 ( .A(\U_1/U_3/U_0/N59 ), .B(\U_1/U_3/U_3/count[0] ), .Y(
        \U_1/U_3/U_3/N84 ) );
  XOR2X1 U9688 ( .A(\U_1/U_0/U_1/U_2/count[7] ), .B(
        \U_1/U_0/U_1/U_2/add_46/carry[7] ), .Y(\U_1/U_0/U_1/U_2/N30 ) );
  AND2X1 U9689 ( .A(\U_1/U_0/U_1/U_2/count[6] ), .B(
        \U_1/U_0/U_1/U_2/add_46/carry[6] ), .Y(
        \U_1/U_0/U_1/U_2/add_46/carry[7] ) );
  XOR2X1 U9690 ( .A(\U_1/U_0/U_1/U_2/add_46/carry[6] ), .B(
        \U_1/U_0/U_1/U_2/count[6] ), .Y(\U_1/U_0/U_1/U_2/N29 ) );
  AND2X1 U9691 ( .A(\U_1/U_0/U_1/U_2/count[5] ), .B(
        \U_1/U_0/U_1/U_2/add_46/carry[5] ), .Y(
        \U_1/U_0/U_1/U_2/add_46/carry[6] ) );
  XOR2X1 U9692 ( .A(\U_1/U_0/U_1/U_2/add_46/carry[5] ), .B(
        \U_1/U_0/U_1/U_2/count[5] ), .Y(\U_1/U_0/U_1/U_2/N28 ) );
  AND2X1 U9693 ( .A(\U_1/U_0/U_1/U_2/count[4] ), .B(
        \U_1/U_0/U_1/U_2/add_46/carry[4] ), .Y(
        \U_1/U_0/U_1/U_2/add_46/carry[5] ) );
  XOR2X1 U9694 ( .A(\U_1/U_0/U_1/U_2/add_46/carry[4] ), .B(
        \U_1/U_0/U_1/U_2/count[4] ), .Y(\U_1/U_0/U_1/U_2/N27 ) );
  AND2X1 U9695 ( .A(\U_1/U_0/U_1/U_2/count[3] ), .B(
        \U_1/U_0/U_1/U_2/add_46/carry[3] ), .Y(
        \U_1/U_0/U_1/U_2/add_46/carry[4] ) );
  XOR2X1 U9696 ( .A(\U_1/U_0/U_1/U_2/add_46/carry[3] ), .B(
        \U_1/U_0/U_1/U_2/count[3] ), .Y(\U_1/U_0/U_1/U_2/N26 ) );
  AND2X1 U9697 ( .A(\U_1/U_0/U_1/U_2/count[2] ), .B(\U_1/U_0/U_1/U_2/count[1] ), .Y(\U_1/U_0/U_1/U_2/add_46/carry[3] ) );
  XOR2X1 U9698 ( .A(\U_1/U_0/U_1/U_2/count[1] ), .B(\U_1/U_0/U_1/U_2/count[2] ), .Y(\U_1/U_0/U_1/U_2/N25 ) );
  OR2X1 U9699 ( .A(n9334), .B(\U_0/U_1/U_1/writeptr[0] ), .Y(
        \U_0/U_1/U_1/sub_72/carry[1] ) );
  XNOR2X1 U9700 ( .A(\U_0/U_1/U_1/writeptr[0] ), .B(n9334), .Y(
        \U_0/U_1/U_1/N189 ) );
  XOR2X1 U9701 ( .A(\U_0/U_1/U_1/readptr[4] ), .B(
        \U_0/U_1/U_1/add_76_aco/carry[4] ), .Y(\U_0/U_1/U_1/N337 ) );
  AND2X1 U9702 ( .A(n9331), .B(\U_0/U_1/U_1/add_76_aco/carry[3] ), .Y(
        \U_0/U_1/U_1/add_76_aco/carry[4] ) );
  XOR2X1 U9703 ( .A(\U_0/U_1/U_1/add_76_aco/carry[3] ), .B(n9331), .Y(
        \U_0/U_1/U_1/N336 ) );
  AND2X1 U9704 ( .A(\U_0/U_1/U_1/readptr[2] ), .B(
        \U_0/U_1/U_1/add_76_aco/carry[2] ), .Y(
        \U_0/U_1/U_1/add_76_aco/carry[3] ) );
  XOR2X1 U9705 ( .A(\U_0/U_1/U_1/add_76_aco/carry[2] ), .B(
        \U_0/U_1/U_1/readptr[2] ), .Y(\U_0/U_1/U_1/N335 ) );
  AND2X1 U9706 ( .A(\U_0/U_1/U_1/readptr[1] ), .B(
        \U_0/U_1/U_1/add_76_aco/carry[1] ), .Y(
        \U_0/U_1/U_1/add_76_aco/carry[2] ) );
  XOR2X1 U9707 ( .A(\U_0/U_1/U_1/add_76_aco/carry[1] ), .B(
        \U_0/U_1/U_1/readptr[1] ), .Y(\U_0/U_1/U_1/N334 ) );
  AND2X1 U9708 ( .A(\U_0/U_1/U_1/readptr[0] ), .B(\U_0/U_1/U_1/N195 ), .Y(
        \U_0/U_1/U_1/add_76_aco/carry[1] ) );
  XOR2X1 U9709 ( .A(\U_0/U_1/U_1/N195 ), .B(\U_0/U_1/U_1/readptr[0] ), .Y(
        \U_0/U_1/U_1/N333 ) );
  XOR2X1 U9710 ( .A(\U_0/U_3/U_3/N188 ), .B(\r2008/carry[6] ), .Y(
        \U_0/U_3/U_3/N90 ) );
  AND2X1 U9711 ( .A(\U_0/U_3/U_3/count[5] ), .B(\r2008/carry[5] ), .Y(
        \r2008/carry[6] ) );
  XOR2X1 U9712 ( .A(\r2008/carry[5] ), .B(\U_0/U_3/U_3/count[5] ), .Y(
        \U_0/U_3/U_3/N89 ) );
  AND2X1 U9713 ( .A(\U_0/U_3/U_3/count[4] ), .B(\r2008/carry[4] ), .Y(
        \r2008/carry[5] ) );
  XOR2X1 U9714 ( .A(\r2008/carry[4] ), .B(\U_0/U_3/U_3/count[4] ), .Y(
        \U_0/U_3/U_3/N88 ) );
  AND2X1 U9715 ( .A(\U_0/U_3/U_3/count[3] ), .B(\r2008/carry[3] ), .Y(
        \r2008/carry[4] ) );
  XOR2X1 U9716 ( .A(\r2008/carry[3] ), .B(\U_0/U_3/U_3/count[3] ), .Y(
        \U_0/U_3/U_3/N87 ) );
  AND2X1 U9717 ( .A(\U_0/U_3/U_3/count[2] ), .B(\r2008/carry[2] ), .Y(
        \r2008/carry[3] ) );
  XOR2X1 U9718 ( .A(\r2008/carry[2] ), .B(\U_0/U_3/U_3/count[2] ), .Y(
        \U_0/U_3/U_3/N86 ) );
  AND2X1 U9719 ( .A(\U_0/U_3/U_3/count[1] ), .B(\r2008/carry[1] ), .Y(
        \r2008/carry[2] ) );
  XOR2X1 U9720 ( .A(\r2008/carry[1] ), .B(\U_0/U_3/U_3/count[1] ), .Y(
        \U_0/U_3/U_3/N85 ) );
  AND2X1 U9721 ( .A(\U_0/U_3/U_3/count[0] ), .B(\U_0/U_3/U_0/N59 ), .Y(
        \r2008/carry[1] ) );
  XOR2X1 U9722 ( .A(\U_0/U_3/U_0/N59 ), .B(\U_0/U_3/U_3/count[0] ), .Y(
        \U_0/U_3/U_3/N84 ) );
  XOR2X1 U9723 ( .A(\U_0/U_0/U_1/U_2/count[7] ), .B(
        \U_0/U_0/U_1/U_2/add_46/carry[7] ), .Y(\U_0/U_0/U_1/U_2/N30 ) );
  AND2X1 U9724 ( .A(\U_0/U_0/U_1/U_2/count[6] ), .B(
        \U_0/U_0/U_1/U_2/add_46/carry[6] ), .Y(
        \U_0/U_0/U_1/U_2/add_46/carry[7] ) );
  XOR2X1 U9725 ( .A(\U_0/U_0/U_1/U_2/add_46/carry[6] ), .B(
        \U_0/U_0/U_1/U_2/count[6] ), .Y(\U_0/U_0/U_1/U_2/N29 ) );
  AND2X1 U9726 ( .A(\U_0/U_0/U_1/U_2/count[5] ), .B(
        \U_0/U_0/U_1/U_2/add_46/carry[5] ), .Y(
        \U_0/U_0/U_1/U_2/add_46/carry[6] ) );
  XOR2X1 U9727 ( .A(\U_0/U_0/U_1/U_2/add_46/carry[5] ), .B(
        \U_0/U_0/U_1/U_2/count[5] ), .Y(\U_0/U_0/U_1/U_2/N28 ) );
  AND2X1 U9728 ( .A(\U_0/U_0/U_1/U_2/count[4] ), .B(
        \U_0/U_0/U_1/U_2/add_46/carry[4] ), .Y(
        \U_0/U_0/U_1/U_2/add_46/carry[5] ) );
  XOR2X1 U9729 ( .A(\U_0/U_0/U_1/U_2/add_46/carry[4] ), .B(
        \U_0/U_0/U_1/U_2/count[4] ), .Y(\U_0/U_0/U_1/U_2/N27 ) );
  AND2X1 U9730 ( .A(\U_0/U_0/U_1/U_2/count[3] ), .B(
        \U_0/U_0/U_1/U_2/add_46/carry[3] ), .Y(
        \U_0/U_0/U_1/U_2/add_46/carry[4] ) );
  XOR2X1 U9731 ( .A(\U_0/U_0/U_1/U_2/add_46/carry[3] ), .B(
        \U_0/U_0/U_1/U_2/count[3] ), .Y(\U_0/U_0/U_1/U_2/N26 ) );
  AND2X1 U9732 ( .A(\U_0/U_0/U_1/U_2/count[2] ), .B(\U_0/U_0/U_1/U_2/count[1] ), .Y(\U_0/U_0/U_1/U_2/add_46/carry[3] ) );
  XOR2X1 U9733 ( .A(\U_0/U_0/U_1/U_2/count[1] ), .B(\U_0/U_0/U_1/U_2/count[2] ), .Y(\U_0/U_0/U_1/U_2/N25 ) );
  NAND2X1 U9734 ( .A(n9544), .B(n11242), .Y(n9535) );
  OAI21X1 U9735 ( .A(n11242), .B(n9544), .C(n9535), .Y(\U_0/U_0/U_0/N442 ) );
  NOR2X1 U9736 ( .A(n9535), .B(\U_0/U_0/U_0/si[2] ), .Y(n9537) );
  AOI21X1 U9737 ( .A(n9535), .B(\U_0/U_0/U_0/si[2] ), .C(n9537), .Y(n9536) );
  NAND2X1 U9738 ( .A(n9537), .B(n9543), .Y(n9538) );
  OAI21X1 U9739 ( .A(n9537), .B(n9543), .C(n9538), .Y(\U_0/U_0/U_0/N444 ) );
  NOR2X1 U9740 ( .A(n9538), .B(\U_0/U_0/U_0/si[4] ), .Y(n9540) );
  AOI21X1 U9741 ( .A(n9538), .B(\U_0/U_0/U_0/si[4] ), .C(n9540), .Y(n9539) );
  NAND2X1 U9742 ( .A(n9540), .B(n11251), .Y(n9541) );
  OAI21X1 U9743 ( .A(n9540), .B(n11251), .C(n9541), .Y(\U_0/U_0/U_0/N446 ) );
  XNOR2X1 U9744 ( .A(\U_0/U_0/U_0/si[6] ), .B(n9541), .Y(\U_0/U_0/U_0/N447 )
         );
  NOR2X1 U9745 ( .A(\U_0/U_0/U_0/si[6] ), .B(n9541), .Y(n9542) );
  XOR2X1 U9746 ( .A(\U_0/U_0/U_0/si[7] ), .B(n9542), .Y(\U_0/U_0/U_0/N448 ) );
  INVX2 U9747 ( .A(\U_0/U_0/U_0/si[3] ), .Y(n9543) );
  INVX2 U9748 ( .A(\U_0/U_0/U_0/si[1] ), .Y(n9544) );
  INVX2 U9749 ( .A(n9539), .Y(\U_0/U_0/U_0/N445 ) );
  INVX2 U9750 ( .A(n9536), .Y(\U_0/U_0/U_0/N443 ) );
  XOR2X1 U9751 ( .A(\r1994/carry[4] ), .B(n9328), .Y(\U_0/U_1/U_1/N35 ) );
  NAND2X1 U9752 ( .A(n9554), .B(n11923), .Y(n9545) );
  OAI21X1 U9753 ( .A(n11923), .B(n9554), .C(n9545), .Y(\U_1/U_0/U_0/N442 ) );
  NOR2X1 U9754 ( .A(n9545), .B(\U_1/U_0/U_0/si[2] ), .Y(n9547) );
  AOI21X1 U9755 ( .A(n9545), .B(\U_1/U_0/U_0/si[2] ), .C(n9547), .Y(n9546) );
  NAND2X1 U9756 ( .A(n9547), .B(n9553), .Y(n9548) );
  OAI21X1 U9757 ( .A(n9547), .B(n9553), .C(n9548), .Y(\U_1/U_0/U_0/N444 ) );
  NOR2X1 U9758 ( .A(n9548), .B(\U_1/U_0/U_0/si[4] ), .Y(n9550) );
  AOI21X1 U9759 ( .A(n9548), .B(\U_1/U_0/U_0/si[4] ), .C(n9550), .Y(n9549) );
  NAND2X1 U9760 ( .A(n9550), .B(n11977), .Y(n9551) );
  OAI21X1 U9761 ( .A(n9550), .B(n11977), .C(n9551), .Y(\U_1/U_0/U_0/N446 ) );
  XNOR2X1 U9762 ( .A(\U_1/U_0/U_0/si[6] ), .B(n9551), .Y(\U_1/U_0/U_0/N447 )
         );
  NOR2X1 U9763 ( .A(\U_1/U_0/U_0/si[6] ), .B(n9551), .Y(n9552) );
  XOR2X1 U9764 ( .A(\U_1/U_0/U_0/si[7] ), .B(n9552), .Y(\U_1/U_0/U_0/N448 ) );
  INVX2 U9765 ( .A(\U_1/U_0/U_0/si[3] ), .Y(n9553) );
  INVX2 U9766 ( .A(\U_1/U_0/U_0/si[1] ), .Y(n9554) );
  INVX2 U9767 ( .A(n9549), .Y(\U_1/U_0/U_0/N445 ) );
  INVX2 U9768 ( .A(n9546), .Y(\U_1/U_0/U_0/N443 ) );
  XOR2X1 U9769 ( .A(\r2028/carry[4] ), .B(n9294), .Y(\U_1/U_1/U_1/N35 ) );
  INVX2 U9770 ( .A(\U_0/U_0/U_1/U_2/count[1] ), .Y(\U_0/U_0/U_1/U_2/N24 ) );
  NOR2X1 U9771 ( .A(n9324), .B(\U_0/U_1/U_1/writeptr[0] ), .Y(n9556) );
  AOI21X1 U9772 ( .A(\U_0/U_1/U_1/writeptr[0] ), .B(n9324), .C(n9556), .Y(
        n9555) );
  NAND2X1 U9773 ( .A(n9556), .B(n9321), .Y(n9557) );
  OAI21X1 U9774 ( .A(n9556), .B(n9321), .C(n9557), .Y(\U_0/U_1/U_1/N44 ) );
  XNOR2X1 U9775 ( .A(n9326), .B(n9557), .Y(\U_0/U_1/U_1/N45 ) );
  NOR2X1 U9776 ( .A(n9326), .B(n9557), .Y(n9558) );
  XOR2X1 U9777 ( .A(\U_0/U_1/U_1/writeptr[4] ), .B(n9558), .Y(
        \U_0/U_1/U_1/N46 ) );
  INVX2 U9778 ( .A(n9555), .Y(\U_0/U_1/U_1/N43 ) );
  XOR2X1 U9779 ( .A(\U_0/U_1/U_1/add_67/carry[4] ), .B(
        \U_0/U_1/U_1/writeptr[4] ), .Y(\U_0/U_1/U_1/N51 ) );
  INVX2 U9780 ( .A(\U_1/U_0/U_1/U_2/count[1] ), .Y(\U_1/U_0/U_1/U_2/N24 ) );
  NOR2X1 U9781 ( .A(n9290), .B(\U_1/U_1/U_1/writeptr[0] ), .Y(n9561) );
  AOI21X1 U9782 ( .A(\U_1/U_1/U_1/writeptr[0] ), .B(n9290), .C(n9561), .Y(
        n9560) );
  NAND2X1 U9783 ( .A(n9561), .B(n9287), .Y(n9562) );
  OAI21X1 U9784 ( .A(n9561), .B(n9287), .C(n9562), .Y(\U_1/U_1/U_1/N44 ) );
  XNOR2X1 U9785 ( .A(n9292), .B(n9562), .Y(\U_1/U_1/U_1/N45 ) );
  NOR2X1 U9786 ( .A(n9292), .B(n9562), .Y(n9563) );
  XOR2X1 U9787 ( .A(\U_1/U_1/U_1/writeptr[4] ), .B(n9563), .Y(
        \U_1/U_1/U_1/N46 ) );
  INVX2 U9788 ( .A(n9560), .Y(\U_1/U_1/U_1/N43 ) );
  XOR2X1 U9789 ( .A(\U_1/U_1/U_1/add_67/carry[4] ), .B(
        \U_1/U_1/U_1/writeptr[4] ), .Y(\U_1/U_1/U_1/N51 ) );
  OAI21X1 U9790 ( .A(\U_0/U_0/U_1/U_2/N23 ), .B(\U_0/U_0/U_1/U_2/count[1] ), 
        .C(\U_0/U_0/U_1/U_2/count[2] ), .Y(n9565) );
  NOR2X1 U9791 ( .A(n9570), .B(n9565), .Y(n9566) );
  OAI21X1 U9792 ( .A(n9566), .B(\U_0/U_0/U_1/U_2/count[4] ), .C(
        \U_0/U_0/U_1/U_2/count[6] ), .Y(n9567) );
  OAI21X1 U9793 ( .A(n9569), .B(n9567), .C(n9568), .Y(\U_0/U_0/U_1/U_2/N99 )
         );
  INVX2 U9794 ( .A(\U_0/U_0/U_1/U_2/count[7] ), .Y(n9568) );
  INVX2 U9795 ( .A(\U_0/U_0/U_1/U_2/count[5] ), .Y(n9569) );
  INVX2 U9796 ( .A(\U_0/U_0/U_1/U_2/count[3] ), .Y(n9570) );
  XNOR2X1 U9797 ( .A(\U_0/U_2/rx_CHECK_CRC [10]), .B(\U_0/U_2/RX_CRC [10]), 
        .Y(n9575) );
  XNOR2X1 U9798 ( .A(\U_0/U_2/rx_CHECK_CRC [9]), .B(\U_0/U_2/RX_CRC [9]), .Y(
        n9574) );
  XOR2X1 U9799 ( .A(\U_0/U_2/rx_CHECK_CRC [7]), .B(\U_0/U_2/RX_CRC [7]), .Y(
        n9572) );
  XOR2X1 U9800 ( .A(\U_0/U_2/rx_CHECK_CRC [8]), .B(\U_0/U_2/RX_CRC [8]), .Y(
        n9571) );
  NOR2X1 U9801 ( .A(n9572), .B(n9571), .Y(n9573) );
  NAND3X1 U9802 ( .A(n9575), .B(n9574), .C(n9573), .Y(n9582) );
  XNOR2X1 U9803 ( .A(\U_0/U_2/rx_CHECK_CRC [14]), .B(\U_0/U_2/RX_CRC [14]), 
        .Y(n9580) );
  XNOR2X1 U9804 ( .A(\U_0/U_2/rx_CHECK_CRC [13]), .B(\U_0/U_2/RX_CRC [13]), 
        .Y(n9579) );
  XOR2X1 U9805 ( .A(\U_0/U_2/rx_CHECK_CRC [11]), .B(\U_0/U_2/RX_CRC [11]), .Y(
        n9577) );
  XOR2X1 U9806 ( .A(\U_0/U_2/rx_CHECK_CRC [12]), .B(\U_0/U_2/RX_CRC [12]), .Y(
        n9576) );
  NOR2X1 U9807 ( .A(n9577), .B(n9576), .Y(n9578) );
  NAND3X1 U9808 ( .A(n9580), .B(n9579), .C(n9578), .Y(n9581) );
  NOR2X1 U9809 ( .A(n9582), .B(n9581), .Y(n9598) );
  NOR2X1 U9810 ( .A(n9601), .B(\U_0/U_2/rx_CHECK_CRC [0]), .Y(n9583) );
  OAI22X1 U9811 ( .A(\U_0/U_2/RX_CRC [1]), .B(n9583), .C(n9583), .D(n9599), 
        .Y(n9589) );
  AND2X1 U9812 ( .A(\U_0/U_2/rx_CHECK_CRC [0]), .B(n9601), .Y(n9584) );
  OAI22X1 U9813 ( .A(n9584), .B(n9600), .C(\U_0/U_2/rx_CHECK_CRC [1]), .D(
        n9584), .Y(n9588) );
  XOR2X1 U9814 ( .A(\U_0/U_2/rx_CHECK_CRC [15]), .B(\U_0/U_2/RX_CRC [15]), .Y(
        n9586) );
  XOR2X1 U9815 ( .A(\U_0/U_2/rx_CHECK_CRC [2]), .B(\U_0/U_2/RX_CRC [2]), .Y(
        n9585) );
  NOR2X1 U9816 ( .A(n9586), .B(n9585), .Y(n9587) );
  NAND3X1 U9817 ( .A(n9589), .B(n9588), .C(n9587), .Y(n9596) );
  XNOR2X1 U9818 ( .A(\U_0/U_2/rx_CHECK_CRC [6]), .B(\U_0/U_2/RX_CRC [6]), .Y(
        n9594) );
  XNOR2X1 U9819 ( .A(\U_0/U_2/rx_CHECK_CRC [5]), .B(\U_0/U_2/RX_CRC [5]), .Y(
        n9593) );
  XOR2X1 U9820 ( .A(\U_0/U_2/rx_CHECK_CRC [3]), .B(\U_0/U_2/RX_CRC [3]), .Y(
        n9591) );
  XOR2X1 U9821 ( .A(\U_0/U_2/rx_CHECK_CRC [4]), .B(\U_0/U_2/RX_CRC [4]), .Y(
        n9590) );
  NOR2X1 U9822 ( .A(n9591), .B(n9590), .Y(n9592) );
  NAND3X1 U9823 ( .A(n9594), .B(n9593), .C(n9592), .Y(n9595) );
  NOR2X1 U9824 ( .A(n9596), .B(n9595), .Y(n9597) );
  AND2X1 U9825 ( .A(n9598), .B(n9597), .Y(\U_0/U_2/U_5/N170 ) );
  INVX2 U9826 ( .A(\U_0/U_2/rx_CHECK_CRC [1]), .Y(n9599) );
  INVX2 U9827 ( .A(\U_0/U_2/RX_CRC [1]), .Y(n9600) );
  INVX2 U9828 ( .A(\U_0/U_2/RX_CRC [0]), .Y(n9601) );
  OAI21X1 U9829 ( .A(\U_1/U_0/U_1/U_2/N23 ), .B(\U_1/U_0/U_1/U_2/count[1] ), 
        .C(\U_1/U_0/U_1/U_2/count[2] ), .Y(n9602) );
  NOR2X1 U9830 ( .A(n9607), .B(n9602), .Y(n9603) );
  OAI21X1 U9831 ( .A(n9603), .B(\U_1/U_0/U_1/U_2/count[4] ), .C(
        \U_1/U_0/U_1/U_2/count[6] ), .Y(n9604) );
  OAI21X1 U9832 ( .A(n9606), .B(n9604), .C(n9605), .Y(\U_1/U_0/U_1/U_2/N99 )
         );
  INVX2 U9833 ( .A(\U_1/U_0/U_1/U_2/count[7] ), .Y(n9605) );
  INVX2 U9834 ( .A(\U_1/U_0/U_1/U_2/count[5] ), .Y(n9606) );
  INVX2 U9835 ( .A(\U_1/U_0/U_1/U_2/count[3] ), .Y(n9607) );
  XNOR2X1 U9836 ( .A(\U_1/U_2/rx_CHECK_CRC [10]), .B(\U_1/U_2/RX_CRC [10]), 
        .Y(n9612) );
  XNOR2X1 U9837 ( .A(\U_1/U_2/rx_CHECK_CRC [9]), .B(\U_1/U_2/RX_CRC [9]), .Y(
        n9611) );
  XOR2X1 U9838 ( .A(\U_1/U_2/rx_CHECK_CRC [7]), .B(\U_1/U_2/RX_CRC [7]), .Y(
        n9609) );
  XOR2X1 U9839 ( .A(\U_1/U_2/rx_CHECK_CRC [8]), .B(\U_1/U_2/RX_CRC [8]), .Y(
        n9608) );
  NOR2X1 U9840 ( .A(n9609), .B(n9608), .Y(n9610) );
  NAND3X1 U9841 ( .A(n9612), .B(n9611), .C(n9610), .Y(n9619) );
  XNOR2X1 U9842 ( .A(\U_1/U_2/rx_CHECK_CRC [14]), .B(\U_1/U_2/RX_CRC [14]), 
        .Y(n9617) );
  XNOR2X1 U9843 ( .A(\U_1/U_2/rx_CHECK_CRC [13]), .B(\U_1/U_2/RX_CRC [13]), 
        .Y(n9616) );
  XOR2X1 U9844 ( .A(\U_1/U_2/rx_CHECK_CRC [11]), .B(\U_1/U_2/RX_CRC [11]), .Y(
        n9614) );
  XOR2X1 U9845 ( .A(\U_1/U_2/rx_CHECK_CRC [12]), .B(\U_1/U_2/RX_CRC [12]), .Y(
        n9613) );
  NOR2X1 U9846 ( .A(n9614), .B(n9613), .Y(n9615) );
  NAND3X1 U9847 ( .A(n9617), .B(n9616), .C(n9615), .Y(n9618) );
  NOR2X1 U9848 ( .A(n9619), .B(n9618), .Y(n9635) );
  NOR2X1 U9849 ( .A(n9638), .B(\U_1/U_2/rx_CHECK_CRC [0]), .Y(n9620) );
  OAI22X1 U9850 ( .A(\U_1/U_2/RX_CRC [1]), .B(n9620), .C(n9620), .D(n9636), 
        .Y(n9626) );
  AND2X1 U9851 ( .A(\U_1/U_2/rx_CHECK_CRC [0]), .B(n9638), .Y(n9621) );
  OAI22X1 U9852 ( .A(n9621), .B(n9637), .C(\U_1/U_2/rx_CHECK_CRC [1]), .D(
        n9621), .Y(n9625) );
  XOR2X1 U9853 ( .A(\U_1/U_2/rx_CHECK_CRC [15]), .B(\U_1/U_2/RX_CRC [15]), .Y(
        n9623) );
  XOR2X1 U9854 ( .A(\U_1/U_2/rx_CHECK_CRC [2]), .B(\U_1/U_2/RX_CRC [2]), .Y(
        n9622) );
  NOR2X1 U9855 ( .A(n9623), .B(n9622), .Y(n9624) );
  NAND3X1 U9856 ( .A(n9626), .B(n9625), .C(n9624), .Y(n9633) );
  XNOR2X1 U9857 ( .A(\U_1/U_2/rx_CHECK_CRC [6]), .B(\U_1/U_2/RX_CRC [6]), .Y(
        n9631) );
  XNOR2X1 U9858 ( .A(\U_1/U_2/rx_CHECK_CRC [5]), .B(\U_1/U_2/RX_CRC [5]), .Y(
        n9630) );
  XOR2X1 U9859 ( .A(\U_1/U_2/rx_CHECK_CRC [3]), .B(\U_1/U_2/RX_CRC [3]), .Y(
        n9628) );
  XOR2X1 U9860 ( .A(\U_1/U_2/rx_CHECK_CRC [4]), .B(\U_1/U_2/RX_CRC [4]), .Y(
        n9627) );
  NOR2X1 U9861 ( .A(n9628), .B(n9627), .Y(n9629) );
  NAND3X1 U9862 ( .A(n9631), .B(n9630), .C(n9629), .Y(n9632) );
  NOR2X1 U9863 ( .A(n9633), .B(n9632), .Y(n9634) );
  AND2X1 U9864 ( .A(n9635), .B(n9634), .Y(\U_1/U_2/U_5/N170 ) );
  INVX2 U9865 ( .A(\U_1/U_2/rx_CHECK_CRC [1]), .Y(n9636) );
  INVX2 U9866 ( .A(\U_1/U_2/RX_CRC [1]), .Y(n9637) );
  INVX2 U9867 ( .A(\U_1/U_2/RX_CRC [0]), .Y(n9638) );
  NOR2X1 U9868 ( .A(\U_1/U_3/U_3/count[3] ), .B(\U_1/U_3/U_3/count[2] ), .Y(
        n9640) );
  NOR2X1 U9869 ( .A(\U_1/U_3/U_3/count[5] ), .B(\U_1/U_3/U_3/count[4] ), .Y(
        n9639) );
  AOI21X1 U9870 ( .A(n9640), .B(n9639), .C(n11644), .Y(\U_1/U_3/U_3/N187 ) );
  NOR2X1 U9871 ( .A(\U_1/U_1/U_0/N39 ), .B(\U_1/U_1/BYTE_COUNT [3]), .Y(n9642)
         );
  NOR2X1 U9872 ( .A(\U_1/U_1/BYTE_COUNT [1]), .B(\U_1/U_1/BYTE_COUNT [0]), .Y(
        n9641) );
  NAND3X1 U9873 ( .A(n9642), .B(n9643), .C(n9641), .Y(\U_1/U_1/U_0/N40 ) );
  INVX2 U9874 ( .A(\U_1/U_1/BYTE_COUNT [2]), .Y(n9643) );
  NOR2X1 U9875 ( .A(\U_0/U_3/U_3/count[3] ), .B(\U_0/U_3/U_3/count[2] ), .Y(
        n9645) );
  NOR2X1 U9876 ( .A(\U_0/U_3/U_3/count[5] ), .B(\U_0/U_3/U_3/count[4] ), .Y(
        n9644) );
  AOI21X1 U9877 ( .A(n9645), .B(n9644), .C(n9335), .Y(\U_0/U_3/U_3/N187 ) );
  NOR2X1 U9878 ( .A(\U_0/U_1/U_0/N39 ), .B(\U_0/U_1/BYTE_COUNT [3]), .Y(n9647)
         );
  NOR2X1 U9879 ( .A(\U_0/U_1/BYTE_COUNT [1]), .B(\U_0/U_1/BYTE_COUNT [0]), .Y(
        n9646) );
  NAND3X1 U9880 ( .A(n9647), .B(n9648), .C(n9646), .Y(\U_0/U_1/U_0/N40 ) );
  INVX2 U9881 ( .A(\U_0/U_1/BYTE_COUNT [2]), .Y(n9648) );
  XNOR2X1 U9882 ( .A(\U_1/U_1/U_1/readptr[4] ), .B(n9294), .Y(n9657) );
  XNOR2X1 U9883 ( .A(n9297), .B(n9292), .Y(n9656) );
  XOR2X1 U9884 ( .A(\U_1/U_1/U_1/readptr[2] ), .B(n9288), .Y(n9654) );
  NOR2X1 U9885 ( .A(n9300), .B(\U_1/U_1/U_1/writeptr[0] ), .Y(n9649) );
  OAI22X1 U9886 ( .A(n9649), .B(n9289), .C(\U_1/U_1/U_1/readptr[1] ), .D(n9649), .Y(n9652) );
  AND2X1 U9887 ( .A(\U_1/U_1/U_1/writeptr[0] ), .B(n9300), .Y(n9650) );
  OAI22X1 U9888 ( .A(n9290), .B(n9650), .C(n9650), .D(n9299), .Y(n9651) );
  NAND2X1 U9889 ( .A(n9652), .B(n9651), .Y(n9653) );
  NOR2X1 U9890 ( .A(n9654), .B(n9653), .Y(n9655) );
  NAND3X1 U9891 ( .A(n9657), .B(n9656), .C(n9655), .Y(\U_1/U_1/U_1/N194 ) );
  INVX2 U9892 ( .A(\U_1/U_1/U_1/N194 ), .Y(\U_1/U_1/U_1/N349 ) );
  XNOR2X1 U9893 ( .A(\U_1/U_1/U_1/readptr[4] ), .B(\U_1/U_1/U_1/N35 ), .Y(
        n9666) );
  XNOR2X1 U9894 ( .A(n9297), .B(\U_1/U_1/U_1/N34 ), .Y(n9665) );
  XOR2X1 U9895 ( .A(\U_1/U_1/U_1/readptr[2] ), .B(\U_1/U_1/U_1/N33 ), .Y(n9663) );
  NOR2X1 U9896 ( .A(n9300), .B(n11669), .Y(n9658) );
  OAI22X1 U9897 ( .A(n9658), .B(n9667), .C(\U_1/U_1/U_1/readptr[1] ), .D(n9658), .Y(n9661) );
  AND2X1 U9898 ( .A(n11669), .B(n9300), .Y(n9659) );
  OAI22X1 U9899 ( .A(\U_1/U_1/U_1/N32 ), .B(n9659), .C(n9659), .D(n9299), .Y(
        n9660) );
  NAND2X1 U9900 ( .A(n9661), .B(n9660), .Y(n9662) );
  NOR2X1 U9901 ( .A(n9663), .B(n9662), .Y(n9664) );
  NAND3X1 U9902 ( .A(n9666), .B(n9665), .C(n9664), .Y(\U_1/U_1/U_1/N36 ) );
  INVX2 U9903 ( .A(\U_1/U_1/U_1/N32 ), .Y(n9667) );
  INVX2 U9904 ( .A(\U_1/U_1/U_1/N36 ), .Y(\U_1/U_1/U_1/N355 ) );
  XNOR2X1 U9905 ( .A(\U_0/U_1/U_1/readptr[4] ), .B(n9328), .Y(n9676) );
  XNOR2X1 U9906 ( .A(n9331), .B(n9326), .Y(n9675) );
  XOR2X1 U9907 ( .A(\U_0/U_1/U_1/readptr[2] ), .B(n9322), .Y(n9673) );
  NOR2X1 U9908 ( .A(n9334), .B(\U_0/U_1/U_1/writeptr[0] ), .Y(n9668) );
  OAI22X1 U9909 ( .A(n9668), .B(n9323), .C(\U_0/U_1/U_1/readptr[1] ), .D(n9668), .Y(n9671) );
  AND2X1 U9910 ( .A(\U_0/U_1/U_1/writeptr[0] ), .B(n9334), .Y(n9669) );
  OAI22X1 U9911 ( .A(n9324), .B(n9669), .C(n9669), .D(n9333), .Y(n9670) );
  NAND2X1 U9912 ( .A(n9671), .B(n9670), .Y(n9672) );
  NOR2X1 U9913 ( .A(n9673), .B(n9672), .Y(n9674) );
  NAND3X1 U9914 ( .A(n9676), .B(n9675), .C(n9674), .Y(\U_0/U_1/U_1/N194 ) );
  INVX2 U9915 ( .A(\U_0/U_1/U_1/N194 ), .Y(\U_0/U_1/U_1/N349 ) );
  XNOR2X1 U9916 ( .A(\U_0/U_1/U_1/readptr[4] ), .B(\U_0/U_1/U_1/N35 ), .Y(
        n9685) );
  XNOR2X1 U9917 ( .A(n9331), .B(\U_0/U_1/U_1/N34 ), .Y(n9684) );
  XOR2X1 U9918 ( .A(\U_0/U_1/U_1/readptr[2] ), .B(\U_0/U_1/U_1/N33 ), .Y(n9682) );
  NOR2X1 U9919 ( .A(n9334), .B(n10917), .Y(n9677) );
  OAI22X1 U9920 ( .A(n9677), .B(n9686), .C(\U_0/U_1/U_1/readptr[1] ), .D(n9677), .Y(n9680) );
  AND2X1 U9921 ( .A(n10917), .B(n9334), .Y(n9678) );
  OAI22X1 U9922 ( .A(\U_0/U_1/U_1/N32 ), .B(n9678), .C(n9678), .D(n9333), .Y(
        n9679) );
  NAND2X1 U9923 ( .A(n9680), .B(n9679), .Y(n9681) );
  NOR2X1 U9924 ( .A(n9682), .B(n9681), .Y(n9683) );
  NAND3X1 U9925 ( .A(n9685), .B(n9684), .C(n9683), .Y(\U_0/U_1/U_1/N36 ) );
  INVX2 U9926 ( .A(\U_0/U_1/U_1/N32 ), .Y(n9686) );
  INVX2 U9927 ( .A(\U_0/U_1/U_1/N36 ), .Y(\U_0/U_1/U_1/N355 ) );
  INVX2 U9928 ( .A(n748), .Y(n9687) );
  INVX2 U9929 ( .A(n747), .Y(n9688) );
  INVX2 U9930 ( .A(n6542), .Y(n9689) );
  INVX2 U9931 ( .A(n4636), .Y(n9691) );
  INVX2 U9932 ( .A(n4628), .Y(n9692) );
  INVX2 U9933 ( .A(n4623), .Y(n9693) );
  INVX2 U9934 ( .A(n4654), .Y(n9694) );
  INVX2 U9935 ( .A(n762), .Y(n9695) );
  INVX2 U9936 ( .A(n761), .Y(n9696) );
  INVX2 U9937 ( .A(n5978), .Y(n9697) );
  INVX2 U9938 ( .A(n2135), .Y(n9699) );
  INVX2 U9939 ( .A(n2127), .Y(n9700) );
  INVX2 U9940 ( .A(n2122), .Y(n9701) );
  INVX2 U9941 ( .A(n2153), .Y(n9702) );
  INVX2 U9942 ( .A(n6555), .Y(n9703) );
  INVX2 U9943 ( .A(n758), .Y(n9704) );
  INVX2 U9944 ( .A(n6560), .Y(n9705) );
  INVX2 U9945 ( .A(n5991), .Y(n9706) );
  INVX2 U9946 ( .A(n772), .Y(n9707) );
  INVX2 U9947 ( .A(n5996), .Y(n9708) );
  INVX2 U9948 ( .A(n6478), .Y(n9709) );
  INVX2 U9949 ( .A(n4662), .Y(n9710) );
  INVX2 U9950 ( .A(n4641), .Y(n9711) );
  INVX2 U9951 ( .A(n6468), .Y(n9712) );
  INVX2 U9952 ( .A(n4513), .Y(n9713) );
  INVX2 U9953 ( .A(n4612), .Y(n9714) );
  INVX2 U9954 ( .A(n5914), .Y(n9715) );
  INVX2 U9955 ( .A(n2161), .Y(n9716) );
  INVX2 U9956 ( .A(n2140), .Y(n9717) );
  INVX2 U9957 ( .A(n5904), .Y(n9718) );
  INVX2 U9958 ( .A(n2012), .Y(n9719) );
  INVX2 U9959 ( .A(n2111), .Y(n9720) );
  INVX2 U9960 ( .A(n5687), .Y(n9721) );
  INVX2 U9961 ( .A(n5694), .Y(n9722) );
  INVX2 U9962 ( .A(n4721), .Y(n9723) );
  INVX2 U9963 ( .A(n4743), .Y(n9724) );
  INVX2 U9964 ( .A(n4676), .Y(n9725) );
  INVX2 U9965 ( .A(n4703), .Y(n9726) );
  INVX2 U9966 ( .A(n4489), .Y(n9727) );
  INVX2 U9967 ( .A(n4487), .Y(n9728) );
  INVX2 U9968 ( .A(n4396), .Y(n9729) );
  INVX2 U9969 ( .A(n4392), .Y(n9730) );
  INVX2 U9970 ( .A(n4385), .Y(n9731) );
  INVX2 U9971 ( .A(n4388), .Y(n9732) );
  INVX2 U9972 ( .A(n4386), .Y(n9733) );
  INVX2 U9973 ( .A(n4380), .Y(n9734) );
  INVX2 U9974 ( .A(n4383), .Y(n9735) );
  INVX2 U9975 ( .A(n4381), .Y(n9736) );
  INVX2 U9976 ( .A(n4375), .Y(n9737) );
  INVX2 U9977 ( .A(n4378), .Y(n9738) );
  INVX2 U9978 ( .A(n4376), .Y(n9739) );
  INVX2 U9979 ( .A(n4365), .Y(n9740) );
  INVX2 U9980 ( .A(n4369), .Y(n9741) );
  INVX2 U9981 ( .A(n4366), .Y(n9742) );
  INVX2 U9982 ( .A(n4485), .Y(n9743) );
  INVX2 U9983 ( .A(n4482), .Y(n9744) );
  INVX2 U9984 ( .A(n4477), .Y(n9745) );
  INVX2 U9985 ( .A(n4480), .Y(n9746) );
  INVX2 U9986 ( .A(n4478), .Y(n9747) );
  INVX2 U9987 ( .A(n4471), .Y(n9748) );
  INVX2 U9988 ( .A(n4474), .Y(n9749) );
  INVX2 U9989 ( .A(n4472), .Y(n9750) );
  INVX2 U9990 ( .A(n4467), .Y(n9751) );
  INVX2 U9991 ( .A(n4470), .Y(n9752) );
  INVX2 U9992 ( .A(n4468), .Y(n9753) );
  INVX2 U9993 ( .A(n4462), .Y(n9754) );
  INVX2 U9994 ( .A(n4465), .Y(n9755) );
  INVX2 U9995 ( .A(n4463), .Y(n9756) );
  INVX2 U9996 ( .A(n4458), .Y(n9757) );
  INVX2 U9997 ( .A(n4461), .Y(n9758) );
  INVX2 U9998 ( .A(n4459), .Y(n9759) );
  INVX2 U9999 ( .A(n4453), .Y(n9760) );
  INVX2 U10000 ( .A(n4456), .Y(n9761) );
  INVX2 U10001 ( .A(n4454), .Y(n9762) );
  INVX2 U10002 ( .A(n4449), .Y(n9763) );
  INVX2 U10003 ( .A(n4452), .Y(n9764) );
  INVX2 U10004 ( .A(n4450), .Y(n9765) );
  INVX2 U10005 ( .A(n4445), .Y(n9766) );
  INVX2 U10006 ( .A(n4448), .Y(n9767) );
  INVX2 U10007 ( .A(n4446), .Y(n9768) );
  INVX2 U10008 ( .A(n4444), .Y(n9769) );
  INVX2 U10009 ( .A(n4442), .Y(n9770) );
  INVX2 U10010 ( .A(n4440), .Y(n9771) );
  INVX2 U10011 ( .A(n4437), .Y(n9772) );
  INVX2 U10012 ( .A(n4432), .Y(n9773) );
  INVX2 U10013 ( .A(n4435), .Y(n9774) );
  INVX2 U10014 ( .A(n4433), .Y(n9775) );
  INVX2 U10015 ( .A(n4427), .Y(n9776) );
  INVX2 U10016 ( .A(n4430), .Y(n9777) );
  INVX2 U10017 ( .A(n4428), .Y(n9778) );
  INVX2 U10018 ( .A(n4422), .Y(n9779) );
  INVX2 U10019 ( .A(n4425), .Y(n9780) );
  INVX2 U10020 ( .A(n4423), .Y(n9781) );
  INVX2 U10021 ( .A(n4418), .Y(n9782) );
  INVX2 U10022 ( .A(n4421), .Y(n9783) );
  INVX2 U10023 ( .A(n4419), .Y(n9784) );
  INVX2 U10024 ( .A(n4411), .Y(n9785) );
  INVX2 U10025 ( .A(n4409), .Y(n9786) );
  INVX2 U10026 ( .A(n4407), .Y(n9787) );
  INVX2 U10027 ( .A(n4402), .Y(n9788) );
  INVX2 U10028 ( .A(n4399), .Y(n9789) );
  INVX2 U10029 ( .A(n4347), .Y(n9794) );
  INVX2 U10030 ( .A(n4350), .Y(n9795) );
  INVX2 U10031 ( .A(n4351), .Y(n9796) );
  INVX2 U10032 ( .A(n4352), .Y(n9797) );
  INVX2 U10033 ( .A(n4353), .Y(n9798) );
  INVX2 U10034 ( .A(n4354), .Y(n9799) );
  INVX2 U10035 ( .A(n4355), .Y(n9800) );
  INVX2 U10036 ( .A(n4356), .Y(n9801) );
  INVX2 U10037 ( .A(n4337), .Y(n9803) );
  INVX2 U10038 ( .A(n4340), .Y(n9804) );
  INVX2 U10039 ( .A(n4341), .Y(n9805) );
  INVX2 U10040 ( .A(n4342), .Y(n9806) );
  INVX2 U10041 ( .A(n4343), .Y(n9807) );
  INVX2 U10042 ( .A(n4344), .Y(n9808) );
  INVX2 U10043 ( .A(n4345), .Y(n9809) );
  INVX2 U10044 ( .A(n4346), .Y(n9810) );
  INVX2 U10045 ( .A(n4327), .Y(n9812) );
  INVX2 U10046 ( .A(n4330), .Y(n9813) );
  INVX2 U10047 ( .A(n4331), .Y(n9814) );
  INVX2 U10048 ( .A(n4332), .Y(n9815) );
  INVX2 U10049 ( .A(n4333), .Y(n9816) );
  INVX2 U10050 ( .A(n4334), .Y(n9817) );
  INVX2 U10051 ( .A(n4335), .Y(n9818) );
  INVX2 U10052 ( .A(n4336), .Y(n9819) );
  INVX2 U10053 ( .A(n4317), .Y(n9821) );
  INVX2 U10054 ( .A(n4320), .Y(n9822) );
  INVX2 U10055 ( .A(n4321), .Y(n9823) );
  INVX2 U10056 ( .A(n4322), .Y(n9824) );
  INVX2 U10057 ( .A(n4323), .Y(n9825) );
  INVX2 U10058 ( .A(n4324), .Y(n9826) );
  INVX2 U10059 ( .A(n4325), .Y(n9827) );
  INVX2 U10060 ( .A(n4326), .Y(n9828) );
  INVX2 U10061 ( .A(n4307), .Y(n9830) );
  INVX2 U10062 ( .A(n4310), .Y(n9831) );
  INVX2 U10063 ( .A(n4311), .Y(n9832) );
  INVX2 U10064 ( .A(n4312), .Y(n9833) );
  INVX2 U10065 ( .A(n4313), .Y(n9834) );
  INVX2 U10066 ( .A(n4314), .Y(n9835) );
  INVX2 U10067 ( .A(n4315), .Y(n9836) );
  INVX2 U10068 ( .A(n4316), .Y(n9837) );
  INVX2 U10069 ( .A(n4297), .Y(n9839) );
  INVX2 U10070 ( .A(n4300), .Y(n9840) );
  INVX2 U10071 ( .A(n4301), .Y(n9841) );
  INVX2 U10072 ( .A(n4302), .Y(n9842) );
  INVX2 U10073 ( .A(n4303), .Y(n9843) );
  INVX2 U10074 ( .A(n4304), .Y(n9844) );
  INVX2 U10075 ( .A(n4305), .Y(n9845) );
  INVX2 U10076 ( .A(n4306), .Y(n9846) );
  INVX2 U10077 ( .A(n4287), .Y(n9848) );
  INVX2 U10078 ( .A(n4290), .Y(n9849) );
  INVX2 U10079 ( .A(n4291), .Y(n9850) );
  INVX2 U10080 ( .A(n4292), .Y(n9851) );
  INVX2 U10081 ( .A(n4293), .Y(n9852) );
  INVX2 U10082 ( .A(n4294), .Y(n9853) );
  INVX2 U10083 ( .A(n4295), .Y(n9854) );
  INVX2 U10084 ( .A(n4296), .Y(n9855) );
  INVX2 U10085 ( .A(n4277), .Y(n9857) );
  INVX2 U10086 ( .A(n4280), .Y(n9858) );
  INVX2 U10087 ( .A(n4281), .Y(n9859) );
  INVX2 U10088 ( .A(n4282), .Y(n9860) );
  INVX2 U10089 ( .A(n4283), .Y(n9861) );
  INVX2 U10090 ( .A(n4284), .Y(n9862) );
  INVX2 U10091 ( .A(n4285), .Y(n9863) );
  INVX2 U10092 ( .A(n4286), .Y(n9864) );
  INVX2 U10093 ( .A(n4259), .Y(n9870) );
  INVX2 U10094 ( .A(n4262), .Y(n9871) );
  INVX2 U10095 ( .A(n4263), .Y(n9872) );
  INVX2 U10096 ( .A(n4264), .Y(n9873) );
  INVX2 U10097 ( .A(n4265), .Y(n9874) );
  INVX2 U10098 ( .A(n4266), .Y(n9875) );
  INVX2 U10099 ( .A(n4267), .Y(n9876) );
  INVX2 U10100 ( .A(n4268), .Y(n9877) );
  INVX2 U10101 ( .A(n4249), .Y(n9879) );
  INVX2 U10102 ( .A(n4252), .Y(n9880) );
  INVX2 U10103 ( .A(n4253), .Y(n9881) );
  INVX2 U10104 ( .A(n4254), .Y(n9882) );
  INVX2 U10105 ( .A(n4255), .Y(n9883) );
  INVX2 U10106 ( .A(n4256), .Y(n9884) );
  INVX2 U10107 ( .A(n4257), .Y(n9885) );
  INVX2 U10108 ( .A(n4258), .Y(n9886) );
  INVX2 U10109 ( .A(n4239), .Y(n9888) );
  INVX2 U10110 ( .A(n4242), .Y(n9889) );
  INVX2 U10111 ( .A(n4243), .Y(n9890) );
  INVX2 U10112 ( .A(n4244), .Y(n9891) );
  INVX2 U10113 ( .A(n4245), .Y(n9892) );
  INVX2 U10114 ( .A(n4246), .Y(n9893) );
  INVX2 U10115 ( .A(n4247), .Y(n9894) );
  INVX2 U10116 ( .A(n4248), .Y(n9895) );
  INVX2 U10117 ( .A(n4229), .Y(n9897) );
  INVX2 U10118 ( .A(n4232), .Y(n9898) );
  INVX2 U10119 ( .A(n4233), .Y(n9899) );
  INVX2 U10120 ( .A(n4234), .Y(n9900) );
  INVX2 U10121 ( .A(n4235), .Y(n9901) );
  INVX2 U10122 ( .A(n4236), .Y(n9902) );
  INVX2 U10123 ( .A(n4237), .Y(n9903) );
  INVX2 U10124 ( .A(n4238), .Y(n9904) );
  INVX2 U10125 ( .A(n9237), .Y(n9909) );
  INVX2 U10126 ( .A(n4193), .Y(n9914) );
  INVX2 U10127 ( .A(n4196), .Y(n9915) );
  INVX2 U10128 ( .A(n4197), .Y(n9916) );
  INVX2 U10129 ( .A(n4198), .Y(n9917) );
  INVX2 U10130 ( .A(n4199), .Y(n9918) );
  INVX2 U10131 ( .A(n4200), .Y(n9919) );
  INVX2 U10132 ( .A(n4201), .Y(n9920) );
  INVX2 U10133 ( .A(n4202), .Y(n9921) );
  INVX2 U10134 ( .A(n4183), .Y(n9923) );
  INVX2 U10135 ( .A(n4186), .Y(n9924) );
  INVX2 U10136 ( .A(n4187), .Y(n9925) );
  INVX2 U10137 ( .A(n4188), .Y(n9926) );
  INVX2 U10138 ( .A(n4189), .Y(n9927) );
  INVX2 U10139 ( .A(n4190), .Y(n9928) );
  INVX2 U10140 ( .A(n4191), .Y(n9929) );
  INVX2 U10141 ( .A(n4192), .Y(n9930) );
  INVX2 U10142 ( .A(n4173), .Y(n9932) );
  INVX2 U10143 ( .A(n4176), .Y(n9933) );
  INVX2 U10144 ( .A(n4177), .Y(n9934) );
  INVX2 U10145 ( .A(n4178), .Y(n9935) );
  INVX2 U10146 ( .A(n4179), .Y(n9936) );
  INVX2 U10147 ( .A(n4180), .Y(n9937) );
  INVX2 U10148 ( .A(n4181), .Y(n9938) );
  INVX2 U10149 ( .A(n4182), .Y(n9939) );
  INVX2 U10150 ( .A(n4163), .Y(n9941) );
  INVX2 U10151 ( .A(n4166), .Y(n9942) );
  INVX2 U10152 ( .A(n4167), .Y(n9943) );
  INVX2 U10153 ( .A(n4168), .Y(n9944) );
  INVX2 U10154 ( .A(n4169), .Y(n9945) );
  INVX2 U10155 ( .A(n4170), .Y(n9946) );
  INVX2 U10156 ( .A(n4171), .Y(n9947) );
  INVX2 U10157 ( .A(n4172), .Y(n9948) );
  INVX2 U10158 ( .A(n4413), .Y(n9950) );
  INVX2 U10159 ( .A(n3587), .Y(n9952) );
  INVX2 U10160 ( .A(n3590), .Y(n9953) );
  INVX2 U10161 ( .A(n3591), .Y(n9954) );
  INVX2 U10162 ( .A(n3596), .Y(n9955) );
  INVX2 U10163 ( .A(n3597), .Y(n9956) );
  INVX2 U10164 ( .A(n3598), .Y(n9957) );
  INVX2 U10165 ( .A(n3599), .Y(n9958) );
  INVX2 U10166 ( .A(n3600), .Y(n9959) );
  INVX2 U10167 ( .A(n3601), .Y(n9960) );
  INVX2 U10168 ( .A(n3602), .Y(n9961) );
  INVX2 U10169 ( .A(n3603), .Y(n9962) );
  INVX2 U10170 ( .A(n3604), .Y(n9963) );
  INVX2 U10171 ( .A(n3605), .Y(n9964) );
  INVX2 U10172 ( .A(n3606), .Y(n9965) );
  INVX2 U10173 ( .A(n3607), .Y(n9966) );
  INVX2 U10174 ( .A(n3608), .Y(n9967) );
  INVX2 U10175 ( .A(n3609), .Y(n9968) );
  INVX2 U10176 ( .A(n3610), .Y(n9969) );
  INVX2 U10177 ( .A(n3611), .Y(n9970) );
  INVX2 U10178 ( .A(n3612), .Y(n9971) );
  INVX2 U10179 ( .A(n3613), .Y(n9972) );
  INVX2 U10180 ( .A(n3614), .Y(n9973) );
  INVX2 U10181 ( .A(n3615), .Y(n9974) );
  INVX2 U10182 ( .A(n3616), .Y(n9975) );
  INVX2 U10183 ( .A(n3617), .Y(n9976) );
  INVX2 U10184 ( .A(n3618), .Y(n9977) );
  INVX2 U10185 ( .A(n3619), .Y(n9978) );
  INVX2 U10186 ( .A(n3620), .Y(n9979) );
  INVX2 U10187 ( .A(n3621), .Y(n9980) );
  INVX2 U10188 ( .A(n3622), .Y(n9981) );
  INVX2 U10189 ( .A(n3623), .Y(n9982) );
  INVX2 U10190 ( .A(n3624), .Y(n9983) );
  INVX2 U10191 ( .A(n3625), .Y(n9984) );
  INVX2 U10192 ( .A(n3626), .Y(n9985) );
  INVX2 U10193 ( .A(n3627), .Y(n9986) );
  INVX2 U10194 ( .A(n3628), .Y(n9987) );
  INVX2 U10195 ( .A(n3629), .Y(n9988) );
  INVX2 U10196 ( .A(n3630), .Y(n9989) );
  INVX2 U10197 ( .A(n3631), .Y(n9990) );
  INVX2 U10198 ( .A(n3632), .Y(n9991) );
  INVX2 U10199 ( .A(n3633), .Y(n9992) );
  INVX2 U10200 ( .A(n3634), .Y(n9993) );
  INVX2 U10201 ( .A(n3635), .Y(n9994) );
  INVX2 U10202 ( .A(n3636), .Y(n9995) );
  INVX2 U10203 ( .A(n3637), .Y(n9996) );
  INVX2 U10204 ( .A(n3638), .Y(n9997) );
  INVX2 U10205 ( .A(n3639), .Y(n9998) );
  INVX2 U10206 ( .A(n3640), .Y(n9999) );
  INVX2 U10207 ( .A(n3641), .Y(n10000) );
  INVX2 U10208 ( .A(n3642), .Y(n10001) );
  INVX2 U10209 ( .A(n3643), .Y(n10002) );
  INVX2 U10210 ( .A(n3644), .Y(n10003) );
  INVX2 U10211 ( .A(n3645), .Y(n10004) );
  INVX2 U10212 ( .A(n3646), .Y(n10005) );
  INVX2 U10213 ( .A(n3647), .Y(n10006) );
  INVX2 U10214 ( .A(n3648), .Y(n10007) );
  INVX2 U10215 ( .A(n3649), .Y(n10008) );
  INVX2 U10216 ( .A(n3650), .Y(n10009) );
  INVX2 U10217 ( .A(n3651), .Y(n10010) );
  INVX2 U10218 ( .A(n3652), .Y(n10011) );
  INVX2 U10219 ( .A(n3515), .Y(n10013) );
  INVX2 U10220 ( .A(n3514), .Y(n10014) );
  INVX2 U10221 ( .A(n3513), .Y(n10015) );
  INVX2 U10222 ( .A(n3512), .Y(n10016) );
  INVX2 U10223 ( .A(n3511), .Y(n10017) );
  INVX2 U10224 ( .A(n3510), .Y(n10018) );
  INVX2 U10225 ( .A(n3509), .Y(n10019) );
  INVX2 U10226 ( .A(n3506), .Y(n10020) );
  INVX2 U10227 ( .A(n3538), .Y(n10021) );
  INVX2 U10228 ( .A(n3656), .Y(n10022) );
  INVX2 U10229 ( .A(n3659), .Y(n10023) );
  INVX2 U10230 ( .A(n3660), .Y(n10024) );
  INVX2 U10231 ( .A(n3661), .Y(n10025) );
  INVX2 U10232 ( .A(n3662), .Y(n10026) );
  INVX2 U10233 ( .A(n3663), .Y(n10027) );
  INVX2 U10234 ( .A(n3664), .Y(n10028) );
  INVX2 U10235 ( .A(n3665), .Y(n10029) );
  INVX2 U10236 ( .A(n3658), .Y(n10030) );
  INVX2 U10237 ( .A(n3586), .Y(n10031) );
  INVX2 U10238 ( .A(n3573), .Y(n10032) );
  INVX2 U10239 ( .A(n3576), .Y(n10033) );
  INVX2 U10240 ( .A(n3577), .Y(n10034) );
  INVX2 U10241 ( .A(n3578), .Y(n10035) );
  INVX2 U10242 ( .A(n3579), .Y(n10036) );
  INVX2 U10243 ( .A(n3580), .Y(n10037) );
  INVX2 U10244 ( .A(n3581), .Y(n10038) );
  INVX2 U10245 ( .A(n3582), .Y(n10039) );
  INVX2 U10246 ( .A(n3666), .Y(n10040) );
  INVX2 U10247 ( .A(n3559), .Y(n10041) );
  INVX2 U10248 ( .A(n3440), .Y(n10042) );
  INVX2 U10249 ( .A(n3460), .Y(n10043) );
  INVX2 U10250 ( .A(n3389), .Y(n10044) );
  INVX2 U10251 ( .A(n3390), .Y(n10045) );
  INVX2 U10252 ( .A(n3391), .Y(n10046) );
  INVX2 U10253 ( .A(n3392), .Y(n10047) );
  INVX2 U10254 ( .A(n3393), .Y(n10048) );
  INVX2 U10255 ( .A(n3394), .Y(n10049) );
  INVX2 U10256 ( .A(n3395), .Y(n10050) );
  INVX2 U10257 ( .A(n9239), .Y(n10051) );
  INVX2 U10258 ( .A(n3186), .Y(n10052) );
  INVX2 U10259 ( .A(n3193), .Y(n10053) );
  INVX2 U10260 ( .A(n2220), .Y(n10054) );
  INVX2 U10261 ( .A(n2242), .Y(n10055) );
  INVX2 U10262 ( .A(n2175), .Y(n10056) );
  INVX2 U10263 ( .A(n2202), .Y(n10057) );
  INVX2 U10264 ( .A(n1986), .Y(n10058) );
  INVX2 U10265 ( .A(n1984), .Y(n10059) );
  INVX2 U10266 ( .A(n1893), .Y(n10060) );
  INVX2 U10267 ( .A(n1889), .Y(n10061) );
  INVX2 U10268 ( .A(n1882), .Y(n10062) );
  INVX2 U10269 ( .A(n1885), .Y(n10063) );
  INVX2 U10270 ( .A(n1883), .Y(n10064) );
  INVX2 U10271 ( .A(n1877), .Y(n10065) );
  INVX2 U10272 ( .A(n1880), .Y(n10066) );
  INVX2 U10273 ( .A(n1878), .Y(n10067) );
  INVX2 U10274 ( .A(n1872), .Y(n10068) );
  INVX2 U10275 ( .A(n1875), .Y(n10069) );
  INVX2 U10276 ( .A(n1873), .Y(n10070) );
  INVX2 U10277 ( .A(n1862), .Y(n10071) );
  INVX2 U10278 ( .A(n1866), .Y(n10072) );
  INVX2 U10279 ( .A(n1863), .Y(n10073) );
  INVX2 U10280 ( .A(n1982), .Y(n10074) );
  INVX2 U10281 ( .A(n1979), .Y(n10075) );
  INVX2 U10282 ( .A(n1974), .Y(n10076) );
  INVX2 U10283 ( .A(n1977), .Y(n10077) );
  INVX2 U10284 ( .A(n1975), .Y(n10078) );
  INVX2 U10285 ( .A(n1968), .Y(n10079) );
  INVX2 U10286 ( .A(n1971), .Y(n10080) );
  INVX2 U10287 ( .A(n1969), .Y(n10081) );
  INVX2 U10288 ( .A(n1964), .Y(n10082) );
  INVX2 U10289 ( .A(n1967), .Y(n10083) );
  INVX2 U10290 ( .A(n1965), .Y(n10084) );
  INVX2 U10291 ( .A(n1959), .Y(n10085) );
  INVX2 U10292 ( .A(n1962), .Y(n10086) );
  INVX2 U10293 ( .A(n1960), .Y(n10087) );
  INVX2 U10294 ( .A(n1955), .Y(n10088) );
  INVX2 U10295 ( .A(n1958), .Y(n10089) );
  INVX2 U10296 ( .A(n1956), .Y(n10090) );
  INVX2 U10297 ( .A(n1950), .Y(n10091) );
  INVX2 U10298 ( .A(n1953), .Y(n10092) );
  INVX2 U10299 ( .A(n1951), .Y(n10093) );
  INVX2 U10300 ( .A(n1946), .Y(n10094) );
  INVX2 U10301 ( .A(n1949), .Y(n10095) );
  INVX2 U10302 ( .A(n1947), .Y(n10096) );
  INVX2 U10303 ( .A(n1942), .Y(n10097) );
  INVX2 U10304 ( .A(n1945), .Y(n10098) );
  INVX2 U10305 ( .A(n1943), .Y(n10099) );
  INVX2 U10306 ( .A(n1941), .Y(n10100) );
  INVX2 U10307 ( .A(n1939), .Y(n10101) );
  INVX2 U10308 ( .A(n1937), .Y(n10102) );
  INVX2 U10309 ( .A(n1934), .Y(n10103) );
  INVX2 U10310 ( .A(n1929), .Y(n10104) );
  INVX2 U10311 ( .A(n1932), .Y(n10105) );
  INVX2 U10312 ( .A(n1930), .Y(n10106) );
  INVX2 U10313 ( .A(n1924), .Y(n10107) );
  INVX2 U10314 ( .A(n1927), .Y(n10108) );
  INVX2 U10315 ( .A(n1925), .Y(n10109) );
  INVX2 U10316 ( .A(n1919), .Y(n10110) );
  INVX2 U10317 ( .A(n1922), .Y(n10111) );
  INVX2 U10318 ( .A(n1920), .Y(n10112) );
  INVX2 U10319 ( .A(n1915), .Y(n10113) );
  INVX2 U10320 ( .A(n1918), .Y(n10114) );
  INVX2 U10321 ( .A(n1916), .Y(n10115) );
  INVX2 U10322 ( .A(n1908), .Y(n10116) );
  INVX2 U10323 ( .A(n1906), .Y(n10117) );
  INVX2 U10324 ( .A(n1904), .Y(n10118) );
  INVX2 U10325 ( .A(n1899), .Y(n10119) );
  INVX2 U10326 ( .A(n1896), .Y(n10120) );
  INVX2 U10327 ( .A(n1844), .Y(n10125) );
  INVX2 U10328 ( .A(n1847), .Y(n10126) );
  INVX2 U10329 ( .A(n1848), .Y(n10127) );
  INVX2 U10330 ( .A(n1849), .Y(n10128) );
  INVX2 U10331 ( .A(n1850), .Y(n10129) );
  INVX2 U10332 ( .A(n1851), .Y(n10130) );
  INVX2 U10333 ( .A(n1852), .Y(n10131) );
  INVX2 U10334 ( .A(n1853), .Y(n10132) );
  INVX2 U10335 ( .A(n1834), .Y(n10134) );
  INVX2 U10336 ( .A(n1837), .Y(n10135) );
  INVX2 U10337 ( .A(n1838), .Y(n10136) );
  INVX2 U10338 ( .A(n1839), .Y(n10137) );
  INVX2 U10339 ( .A(n1840), .Y(n10138) );
  INVX2 U10340 ( .A(n1841), .Y(n10139) );
  INVX2 U10341 ( .A(n1842), .Y(n10140) );
  INVX2 U10342 ( .A(n1843), .Y(n10141) );
  INVX2 U10343 ( .A(n1824), .Y(n10143) );
  INVX2 U10344 ( .A(n1827), .Y(n10144) );
  INVX2 U10345 ( .A(n1828), .Y(n10145) );
  INVX2 U10346 ( .A(n1829), .Y(n10146) );
  INVX2 U10347 ( .A(n1830), .Y(n10147) );
  INVX2 U10348 ( .A(n1831), .Y(n10148) );
  INVX2 U10349 ( .A(n1832), .Y(n10149) );
  INVX2 U10350 ( .A(n1833), .Y(n10150) );
  INVX2 U10351 ( .A(n1814), .Y(n10152) );
  INVX2 U10352 ( .A(n1817), .Y(n10153) );
  INVX2 U10353 ( .A(n1818), .Y(n10154) );
  INVX2 U10354 ( .A(n1819), .Y(n10155) );
  INVX2 U10355 ( .A(n1820), .Y(n10156) );
  INVX2 U10356 ( .A(n1821), .Y(n10157) );
  INVX2 U10357 ( .A(n1822), .Y(n10158) );
  INVX2 U10358 ( .A(n1823), .Y(n10159) );
  INVX2 U10359 ( .A(n1804), .Y(n10161) );
  INVX2 U10360 ( .A(n1807), .Y(n10162) );
  INVX2 U10361 ( .A(n1808), .Y(n10163) );
  INVX2 U10362 ( .A(n1809), .Y(n10164) );
  INVX2 U10363 ( .A(n1810), .Y(n10165) );
  INVX2 U10364 ( .A(n1811), .Y(n10166) );
  INVX2 U10365 ( .A(n1812), .Y(n10167) );
  INVX2 U10366 ( .A(n1813), .Y(n10168) );
  INVX2 U10367 ( .A(n1794), .Y(n10170) );
  INVX2 U10368 ( .A(n1797), .Y(n10171) );
  INVX2 U10369 ( .A(n1798), .Y(n10172) );
  INVX2 U10370 ( .A(n1799), .Y(n10173) );
  INVX2 U10371 ( .A(n1800), .Y(n10174) );
  INVX2 U10372 ( .A(n1801), .Y(n10175) );
  INVX2 U10373 ( .A(n1802), .Y(n10176) );
  INVX2 U10374 ( .A(n1803), .Y(n10177) );
  INVX2 U10375 ( .A(n1784), .Y(n10179) );
  INVX2 U10376 ( .A(n1787), .Y(n10180) );
  INVX2 U10377 ( .A(n1788), .Y(n10181) );
  INVX2 U10378 ( .A(n1789), .Y(n10182) );
  INVX2 U10379 ( .A(n1790), .Y(n10183) );
  INVX2 U10380 ( .A(n1791), .Y(n10184) );
  INVX2 U10381 ( .A(n1792), .Y(n10185) );
  INVX2 U10382 ( .A(n1793), .Y(n10186) );
  INVX2 U10383 ( .A(n1774), .Y(n10188) );
  INVX2 U10384 ( .A(n1777), .Y(n10189) );
  INVX2 U10385 ( .A(n1778), .Y(n10190) );
  INVX2 U10386 ( .A(n1779), .Y(n10191) );
  INVX2 U10387 ( .A(n1780), .Y(n10192) );
  INVX2 U10388 ( .A(n1781), .Y(n10193) );
  INVX2 U10389 ( .A(n1782), .Y(n10194) );
  INVX2 U10390 ( .A(n1783), .Y(n10195) );
  INVX2 U10391 ( .A(n1756), .Y(n10201) );
  INVX2 U10392 ( .A(n1759), .Y(n10202) );
  INVX2 U10393 ( .A(n1760), .Y(n10203) );
  INVX2 U10394 ( .A(n1761), .Y(n10204) );
  INVX2 U10395 ( .A(n1762), .Y(n10205) );
  INVX2 U10396 ( .A(n1763), .Y(n10206) );
  INVX2 U10397 ( .A(n1764), .Y(n10207) );
  INVX2 U10398 ( .A(n1765), .Y(n10208) );
  INVX2 U10399 ( .A(n1746), .Y(n10210) );
  INVX2 U10400 ( .A(n1749), .Y(n10211) );
  INVX2 U10401 ( .A(n1750), .Y(n10212) );
  INVX2 U10402 ( .A(n1751), .Y(n10213) );
  INVX2 U10403 ( .A(n1752), .Y(n10214) );
  INVX2 U10404 ( .A(n1753), .Y(n10215) );
  INVX2 U10405 ( .A(n1754), .Y(n10216) );
  INVX2 U10406 ( .A(n1755), .Y(n10217) );
  INVX2 U10407 ( .A(n1736), .Y(n10219) );
  INVX2 U10408 ( .A(n1739), .Y(n10220) );
  INVX2 U10409 ( .A(n1740), .Y(n10221) );
  INVX2 U10410 ( .A(n1741), .Y(n10222) );
  INVX2 U10411 ( .A(n1742), .Y(n10223) );
  INVX2 U10412 ( .A(n1743), .Y(n10224) );
  INVX2 U10413 ( .A(n1744), .Y(n10225) );
  INVX2 U10414 ( .A(n1745), .Y(n10226) );
  INVX2 U10415 ( .A(n1726), .Y(n10228) );
  INVX2 U10416 ( .A(n1729), .Y(n10229) );
  INVX2 U10417 ( .A(n1730), .Y(n10230) );
  INVX2 U10418 ( .A(n1731), .Y(n10231) );
  INVX2 U10419 ( .A(n1732), .Y(n10232) );
  INVX2 U10420 ( .A(n1733), .Y(n10233) );
  INVX2 U10421 ( .A(n1734), .Y(n10234) );
  INVX2 U10422 ( .A(n1735), .Y(n10235) );
  INVX2 U10423 ( .A(n9275), .Y(n10240) );
  INVX2 U10424 ( .A(n1690), .Y(n10245) );
  INVX2 U10425 ( .A(n1693), .Y(n10246) );
  INVX2 U10426 ( .A(n1694), .Y(n10247) );
  INVX2 U10427 ( .A(n1695), .Y(n10248) );
  INVX2 U10428 ( .A(n1696), .Y(n10249) );
  INVX2 U10429 ( .A(n1697), .Y(n10250) );
  INVX2 U10430 ( .A(n1698), .Y(n10251) );
  INVX2 U10431 ( .A(n1699), .Y(n10252) );
  INVX2 U10432 ( .A(n1680), .Y(n10254) );
  INVX2 U10433 ( .A(n1683), .Y(n10255) );
  INVX2 U10434 ( .A(n1684), .Y(n10256) );
  INVX2 U10435 ( .A(n1685), .Y(n10257) );
  INVX2 U10436 ( .A(n1686), .Y(n10258) );
  INVX2 U10437 ( .A(n1687), .Y(n10259) );
  INVX2 U10438 ( .A(n1688), .Y(n10260) );
  INVX2 U10439 ( .A(n1689), .Y(n10261) );
  INVX2 U10440 ( .A(n1670), .Y(n10263) );
  INVX2 U10441 ( .A(n1673), .Y(n10264) );
  INVX2 U10442 ( .A(n1674), .Y(n10265) );
  INVX2 U10443 ( .A(n1675), .Y(n10266) );
  INVX2 U10444 ( .A(n1676), .Y(n10267) );
  INVX2 U10445 ( .A(n1677), .Y(n10268) );
  INVX2 U10446 ( .A(n1678), .Y(n10269) );
  INVX2 U10447 ( .A(n1679), .Y(n10270) );
  INVX2 U10448 ( .A(n1660), .Y(n10272) );
  INVX2 U10449 ( .A(n1663), .Y(n10273) );
  INVX2 U10450 ( .A(n1664), .Y(n10274) );
  INVX2 U10451 ( .A(n1665), .Y(n10275) );
  INVX2 U10452 ( .A(n1666), .Y(n10276) );
  INVX2 U10453 ( .A(n1667), .Y(n10277) );
  INVX2 U10454 ( .A(n1668), .Y(n10278) );
  INVX2 U10455 ( .A(n1669), .Y(n10279) );
  INVX2 U10456 ( .A(n1910), .Y(n10281) );
  INVX2 U10457 ( .A(n1102), .Y(n10283) );
  INVX2 U10458 ( .A(n1105), .Y(n10284) );
  INVX2 U10459 ( .A(n1106), .Y(n10285) );
  INVX2 U10460 ( .A(n1111), .Y(n10286) );
  INVX2 U10461 ( .A(n1112), .Y(n10287) );
  INVX2 U10462 ( .A(n1113), .Y(n10288) );
  INVX2 U10463 ( .A(n1114), .Y(n10289) );
  INVX2 U10464 ( .A(n1115), .Y(n10290) );
  INVX2 U10465 ( .A(n1116), .Y(n10291) );
  INVX2 U10466 ( .A(n1117), .Y(n10292) );
  INVX2 U10467 ( .A(n1118), .Y(n10293) );
  INVX2 U10468 ( .A(n1119), .Y(n10294) );
  INVX2 U10469 ( .A(n1120), .Y(n10295) );
  INVX2 U10470 ( .A(n1121), .Y(n10296) );
  INVX2 U10471 ( .A(n1122), .Y(n10297) );
  INVX2 U10472 ( .A(n1123), .Y(n10298) );
  INVX2 U10473 ( .A(n1124), .Y(n10299) );
  INVX2 U10474 ( .A(n1125), .Y(n10300) );
  INVX2 U10475 ( .A(n1126), .Y(n10301) );
  INVX2 U10476 ( .A(n1127), .Y(n10302) );
  INVX2 U10477 ( .A(n1128), .Y(n10303) );
  INVX2 U10478 ( .A(n1129), .Y(n10304) );
  INVX2 U10479 ( .A(n1130), .Y(n10305) );
  INVX2 U10480 ( .A(n1131), .Y(n10306) );
  INVX2 U10481 ( .A(n1132), .Y(n10307) );
  INVX2 U10482 ( .A(n1133), .Y(n10308) );
  INVX2 U10483 ( .A(n1134), .Y(n10309) );
  INVX2 U10484 ( .A(n1135), .Y(n10310) );
  INVX2 U10485 ( .A(n1136), .Y(n10311) );
  INVX2 U10486 ( .A(n1137), .Y(n10312) );
  INVX2 U10487 ( .A(n1138), .Y(n10313) );
  INVX2 U10488 ( .A(n1139), .Y(n10314) );
  INVX2 U10489 ( .A(n1140), .Y(n10315) );
  INVX2 U10490 ( .A(n1141), .Y(n10316) );
  INVX2 U10491 ( .A(n1142), .Y(n10317) );
  INVX2 U10492 ( .A(n1143), .Y(n10318) );
  INVX2 U10493 ( .A(n1144), .Y(n10319) );
  INVX2 U10494 ( .A(n1145), .Y(n10320) );
  INVX2 U10495 ( .A(n1146), .Y(n10321) );
  INVX2 U10496 ( .A(n1147), .Y(n10322) );
  INVX2 U10497 ( .A(n1148), .Y(n10323) );
  INVX2 U10498 ( .A(n1149), .Y(n10324) );
  INVX2 U10499 ( .A(n1150), .Y(n10325) );
  INVX2 U10500 ( .A(n1151), .Y(n10326) );
  INVX2 U10501 ( .A(n1152), .Y(n10327) );
  INVX2 U10502 ( .A(n1153), .Y(n10328) );
  INVX2 U10503 ( .A(n1154), .Y(n10329) );
  INVX2 U10504 ( .A(n1155), .Y(n10330) );
  INVX2 U10505 ( .A(n1156), .Y(n10331) );
  INVX2 U10506 ( .A(n1157), .Y(n10332) );
  INVX2 U10507 ( .A(n1158), .Y(n10333) );
  INVX2 U10508 ( .A(n1159), .Y(n10334) );
  INVX2 U10509 ( .A(n1160), .Y(n10335) );
  INVX2 U10510 ( .A(n1161), .Y(n10336) );
  INVX2 U10511 ( .A(n1162), .Y(n10337) );
  INVX2 U10512 ( .A(n1163), .Y(n10338) );
  INVX2 U10513 ( .A(n1164), .Y(n10339) );
  INVX2 U10514 ( .A(n1165), .Y(n10340) );
  INVX2 U10515 ( .A(n1166), .Y(n10341) );
  INVX2 U10516 ( .A(n1167), .Y(n10342) );
  INVX2 U10517 ( .A(n926), .Y(n10343) );
  INVX2 U10518 ( .A(n722), .Y(n10344) );
  INVX2 U10519 ( .A(n721), .Y(n10345) );
  INVX2 U10520 ( .A(n720), .Y(n10346) );
  INVX2 U10521 ( .A(n719), .Y(n10347) );
  INVX2 U10522 ( .A(n718), .Y(n10348) );
  INVX2 U10523 ( .A(n717), .Y(n10349) );
  INVX2 U10524 ( .A(n716), .Y(n10350) );
  INVX2 U10525 ( .A(n715), .Y(n10351) );
  INVX2 U10526 ( .A(n714), .Y(n10352) );
  INVX2 U10527 ( .A(n713), .Y(n10353) );
  INVX2 U10528 ( .A(n712), .Y(n10354) );
  INVX2 U10529 ( .A(n711), .Y(n10355) );
  INVX2 U10530 ( .A(n710), .Y(n10356) );
  INVX2 U10531 ( .A(n709), .Y(n10357) );
  INVX2 U10532 ( .A(n708), .Y(n10358) );
  INVX2 U10533 ( .A(n707), .Y(n10359) );
  INVX2 U10534 ( .A(n706), .Y(n10360) );
  INVX2 U10535 ( .A(n705), .Y(n10361) );
  INVX2 U10536 ( .A(n704), .Y(n10362) );
  INVX2 U10537 ( .A(n703), .Y(n10363) );
  INVX2 U10538 ( .A(n702), .Y(n10364) );
  INVX2 U10539 ( .A(n701), .Y(n10365) );
  INVX2 U10540 ( .A(n700), .Y(n10366) );
  INVX2 U10541 ( .A(n699), .Y(n10367) );
  INVX2 U10542 ( .A(n698), .Y(n10368) );
  INVX2 U10543 ( .A(n697), .Y(n10369) );
  INVX2 U10544 ( .A(n696), .Y(n10370) );
  INVX2 U10545 ( .A(n695), .Y(n10371) );
  INVX2 U10546 ( .A(n694), .Y(n10372) );
  INVX2 U10547 ( .A(n693), .Y(n10373) );
  INVX2 U10548 ( .A(n692), .Y(n10374) );
  INVX2 U10549 ( .A(n691), .Y(n10375) );
  INVX2 U10550 ( .A(n690), .Y(n10376) );
  INVX2 U10551 ( .A(n689), .Y(n10377) );
  INVX2 U10552 ( .A(n688), .Y(n10378) );
  INVX2 U10553 ( .A(n687), .Y(n10379) );
  INVX2 U10554 ( .A(n686), .Y(n10380) );
  INVX2 U10555 ( .A(n685), .Y(n10381) );
  INVX2 U10556 ( .A(n684), .Y(n10382) );
  INVX2 U10557 ( .A(n683), .Y(n10383) );
  INVX2 U10558 ( .A(n682), .Y(n10384) );
  INVX2 U10559 ( .A(n681), .Y(n10385) );
  INVX2 U10560 ( .A(n680), .Y(n10386) );
  INVX2 U10561 ( .A(n679), .Y(n10387) );
  INVX2 U10562 ( .A(n678), .Y(n10388) );
  INVX2 U10563 ( .A(n677), .Y(n10389) );
  INVX2 U10564 ( .A(n676), .Y(n10390) );
  INVX2 U10565 ( .A(n675), .Y(n10391) );
  INVX2 U10566 ( .A(n674), .Y(n10392) );
  INVX2 U10567 ( .A(n673), .Y(n10393) );
  INVX2 U10568 ( .A(n672), .Y(n10394) );
  INVX2 U10569 ( .A(n671), .Y(n10395) );
  INVX2 U10570 ( .A(n670), .Y(n10396) );
  INVX2 U10571 ( .A(n669), .Y(n10397) );
  INVX2 U10572 ( .A(n668), .Y(n10398) );
  INVX2 U10573 ( .A(n667), .Y(n10399) );
  INVX2 U10574 ( .A(n666), .Y(n10400) );
  INVX2 U10575 ( .A(n665), .Y(n10401) );
  INVX2 U10576 ( .A(n664), .Y(n10402) );
  INVX2 U10577 ( .A(n656), .Y(n10403) );
  INVX2 U10578 ( .A(n655), .Y(n10404) );
  INVX2 U10579 ( .A(n598), .Y(n10405) );
  INVX2 U10580 ( .A(n597), .Y(n10406) );
  INVX2 U10581 ( .A(n596), .Y(n10407) );
  INVX2 U10582 ( .A(n595), .Y(n10408) );
  INVX2 U10583 ( .A(n594), .Y(n10409) );
  INVX2 U10584 ( .A(n593), .Y(n10410) );
  INVX2 U10585 ( .A(n592), .Y(n10411) );
  INVX2 U10586 ( .A(n591), .Y(n10412) );
  INVX2 U10587 ( .A(n551), .Y(n10413) );
  INVX2 U10588 ( .A(n548), .Y(n10414) );
  INVX2 U10589 ( .A(n545), .Y(n10415) );
  INVX2 U10590 ( .A(n542), .Y(n10416) );
  INVX2 U10591 ( .A(n539), .Y(n10417) );
  INVX2 U10592 ( .A(n536), .Y(n10418) );
  INVX2 U10593 ( .A(n533), .Y(n10419) );
  INVX2 U10594 ( .A(n530), .Y(n10420) );
  INVX2 U10595 ( .A(n470), .Y(n10421) );
  INVX2 U10596 ( .A(n438), .Y(n10422) );
  INVX2 U10597 ( .A(n437), .Y(n10423) );
  INVX2 U10598 ( .A(n436), .Y(n10424) );
  INVX2 U10599 ( .A(n435), .Y(n10425) );
  INVX2 U10600 ( .A(n434), .Y(n10426) );
  INVX2 U10601 ( .A(n433), .Y(n10427) );
  INVX2 U10602 ( .A(n432), .Y(n10428) );
  INVX2 U10603 ( .A(n431), .Y(n10429) );
  INVX2 U10604 ( .A(n430), .Y(n10430) );
  INVX2 U10605 ( .A(n429), .Y(n10431) );
  INVX2 U10606 ( .A(n428), .Y(n10432) );
  INVX2 U10607 ( .A(n427), .Y(n10433) );
  INVX2 U10608 ( .A(n426), .Y(n10434) );
  INVX2 U10609 ( .A(n425), .Y(n10435) );
  INVX2 U10610 ( .A(n424), .Y(n10436) );
  INVX2 U10611 ( .A(n423), .Y(n10437) );
  INVX2 U10612 ( .A(n422), .Y(n10438) );
  INVX2 U10613 ( .A(n421), .Y(n10439) );
  INVX2 U10614 ( .A(n420), .Y(n10440) );
  INVX2 U10615 ( .A(n419), .Y(n10441) );
  INVX2 U10616 ( .A(n418), .Y(n10442) );
  INVX2 U10617 ( .A(n417), .Y(n10443) );
  INVX2 U10618 ( .A(n416), .Y(n10444) );
  INVX2 U10619 ( .A(n415), .Y(n10445) );
  INVX2 U10620 ( .A(n414), .Y(n10446) );
  INVX2 U10621 ( .A(n413), .Y(n10447) );
  INVX2 U10622 ( .A(n412), .Y(n10448) );
  INVX2 U10623 ( .A(n411), .Y(n10449) );
  INVX2 U10624 ( .A(n410), .Y(n10450) );
  INVX2 U10625 ( .A(n409), .Y(n10451) );
  INVX2 U10626 ( .A(n408), .Y(n10452) );
  INVX2 U10627 ( .A(n407), .Y(n10453) );
  INVX2 U10628 ( .A(n406), .Y(n10454) );
  INVX2 U10629 ( .A(n405), .Y(n10455) );
  INVX2 U10630 ( .A(n404), .Y(n10456) );
  INVX2 U10631 ( .A(n403), .Y(n10457) );
  INVX2 U10632 ( .A(n402), .Y(n10458) );
  INVX2 U10633 ( .A(n401), .Y(n10459) );
  INVX2 U10634 ( .A(n400), .Y(n10460) );
  INVX2 U10635 ( .A(n399), .Y(n10461) );
  INVX2 U10636 ( .A(n398), .Y(n10462) );
  INVX2 U10637 ( .A(n397), .Y(n10463) );
  INVX2 U10638 ( .A(n396), .Y(n10464) );
  INVX2 U10639 ( .A(n395), .Y(n10465) );
  INVX2 U10640 ( .A(n394), .Y(n10466) );
  INVX2 U10641 ( .A(n393), .Y(n10467) );
  INVX2 U10642 ( .A(n392), .Y(n10468) );
  INVX2 U10643 ( .A(n391), .Y(n10469) );
  INVX2 U10644 ( .A(n390), .Y(n10470) );
  INVX2 U10645 ( .A(n389), .Y(n10471) );
  INVX2 U10646 ( .A(n388), .Y(n10472) );
  INVX2 U10647 ( .A(n387), .Y(n10473) );
  INVX2 U10648 ( .A(n386), .Y(n10474) );
  INVX2 U10649 ( .A(n385), .Y(n10475) );
  INVX2 U10650 ( .A(n384), .Y(n10476) );
  INVX2 U10651 ( .A(n383), .Y(n10477) );
  INVX2 U10652 ( .A(n382), .Y(n10478) );
  INVX2 U10653 ( .A(n381), .Y(n10479) );
  INVX2 U10654 ( .A(n380), .Y(n10480) );
  INVX2 U10655 ( .A(n372), .Y(n10481) );
  INVX2 U10656 ( .A(n371), .Y(n10482) );
  INVX2 U10657 ( .A(n297), .Y(n10483) );
  INVX2 U10658 ( .A(n294), .Y(n10484) );
  INVX2 U10659 ( .A(n293), .Y(n10485) );
  INVX2 U10660 ( .A(n290), .Y(n10486) );
  INVX2 U10661 ( .A(n287), .Y(n10487) );
  INVX2 U10662 ( .A(n286), .Y(n10488) );
  INVX2 U10663 ( .A(n283), .Y(n10489) );
  INVX2 U10664 ( .A(n280), .Y(n10490) );
  INVX2 U10665 ( .A(n279), .Y(n10491) );
  INVX2 U10666 ( .A(n276), .Y(n10492) );
  INVX2 U10667 ( .A(n273), .Y(n10493) );
  INVX2 U10668 ( .A(n272), .Y(n10494) );
  INVX2 U10669 ( .A(n269), .Y(n10495) );
  INVX2 U10670 ( .A(n266), .Y(n10496) );
  INVX2 U10671 ( .A(n265), .Y(n10497) );
  INVX2 U10672 ( .A(n262), .Y(n10498) );
  INVX2 U10673 ( .A(n259), .Y(n10499) );
  INVX2 U10674 ( .A(n258), .Y(n10500) );
  INVX2 U10675 ( .A(n255), .Y(n10501) );
  INVX2 U10676 ( .A(n252), .Y(n10502) );
  INVX2 U10677 ( .A(n251), .Y(n10503) );
  INVX2 U10678 ( .A(n248), .Y(n10504) );
  INVX2 U10679 ( .A(n245), .Y(n10505) );
  INVX2 U10680 ( .A(n244), .Y(n10506) );
  INVX2 U10681 ( .A(n232), .Y(n10507) );
  INVX2 U10682 ( .A(n184), .Y(n10508) );
  INVX2 U10683 ( .A(n867), .Y(n10511) );
  INVX2 U10684 ( .A(n868), .Y(n10512) );
  INVX2 U10685 ( .A(n869), .Y(n10513) );
  INVX2 U10686 ( .A(n870), .Y(n10514) );
  INVX2 U10687 ( .A(n871), .Y(n10515) );
  INVX2 U10688 ( .A(n872), .Y(n10516) );
  INVX2 U10689 ( .A(n873), .Y(n10517) );
  INVX2 U10690 ( .A(n917), .Y(n10518) );
  INVX2 U10691 ( .A(n1003), .Y(n10519) );
  INVX2 U10692 ( .A(n1010), .Y(n10520) );
  INVX2 U10693 ( .A(n1021), .Y(n10521) );
  INVX2 U10694 ( .A(n1024), .Y(n10522) );
  INVX2 U10695 ( .A(n1025), .Y(n10523) );
  INVX2 U10696 ( .A(n1026), .Y(n10524) );
  INVX2 U10697 ( .A(n1027), .Y(n10525) );
  INVX2 U10698 ( .A(n1028), .Y(n10526) );
  INVX2 U10699 ( .A(n1029), .Y(n10527) );
  INVX2 U10700 ( .A(n1030), .Y(n10528) );
  INVX2 U10701 ( .A(n1022), .Y(n10529) );
  INVX2 U10702 ( .A(n1032), .Y(n10530) );
  INVX2 U10703 ( .A(n1055), .Y(n10531) );
  INVX2 U10704 ( .A(n1058), .Y(n10532) );
  INVX2 U10705 ( .A(n1059), .Y(n10533) );
  INVX2 U10706 ( .A(n1060), .Y(n10534) );
  INVX2 U10707 ( .A(n1061), .Y(n10535) );
  INVX2 U10708 ( .A(n1062), .Y(n10536) );
  INVX2 U10709 ( .A(n1063), .Y(n10537) );
  INVX2 U10710 ( .A(n1064), .Y(n10538) );
  INVX2 U10711 ( .A(n3167), .Y(n10539) );
  INVX2 U10712 ( .A(n3168), .Y(n10540) );
  INVX2 U10713 ( .A(n5668), .Y(n10541) );
  INVX2 U10714 ( .A(n5669), .Y(n10542) );
  INVX2 U10715 ( .A(SERIAL_IN), .Y(n10543) );
  INVX2 U10716 ( .A(\U_0/U_0/U_0/nfdata[7] ), .Y(n10544) );
  INVX2 U10717 ( .A(\U_0/U_0/U_0/nfdata[6] ), .Y(n10545) );
  INVX2 U10718 ( .A(\U_0/U_0/U_0/nfdata[5] ), .Y(n10546) );
  INVX2 U10719 ( .A(\U_0/U_0/U_0/nfdata[4] ), .Y(n10547) );
  INVX2 U10720 ( .A(\U_0/U_0/U_0/nfdata[3] ), .Y(n10548) );
  INVX2 U10721 ( .A(\U_0/U_0/U_0/nfdata[2] ), .Y(n10549) );
  INVX2 U10722 ( .A(\U_0/U_0/U_0/nfdata[1] ), .Y(n10550) );
  INVX2 U10723 ( .A(\U_0/U_0/U_0/nfdata[0] ), .Y(n10551) );
  INVX2 U10724 ( .A(\U_1/U_0/U_0/nfdata[7] ), .Y(n10552) );
  INVX2 U10725 ( .A(\U_1/U_0/U_0/nfdata[6] ), .Y(n10553) );
  INVX2 U10726 ( .A(\U_1/U_0/U_0/nfdata[5] ), .Y(n10554) );
  INVX2 U10727 ( .A(\U_1/U_0/U_0/nfdata[4] ), .Y(n10555) );
  INVX2 U10728 ( .A(\U_1/U_0/U_0/nfdata[3] ), .Y(n10556) );
  INVX2 U10729 ( .A(\U_1/U_0/U_0/nfdata[2] ), .Y(n10557) );
  INVX2 U10730 ( .A(\U_1/U_0/U_0/nfdata[1] ), .Y(n10558) );
  INVX2 U10731 ( .A(\U_1/U_0/U_0/nfdata[0] ), .Y(n10559) );
  INVX2 U10732 ( .A(\U_0/U_0/U_1/U_2/nextState[0] ), .Y(n10560) );
  INVX2 U10733 ( .A(\U_0/U_0/U_1/U_7/nextState[7] ), .Y(n10561) );
  INVX2 U10734 ( .A(\U_0/U_0/U_1/U_7/nextState[6] ), .Y(n10562) );
  INVX2 U10735 ( .A(n5766), .Y(n10563) );
  INVX2 U10736 ( .A(\U_0/U_0/U_1/U_7/nextState[5] ), .Y(n10564) );
  INVX2 U10737 ( .A(\U_0/U_0/U_1/U_7/state[5] ), .Y(n10565) );
  INVX2 U10738 ( .A(\U_0/U_0/U_1/STOP_DATA [1]), .Y(n10566) );
  INVX2 U10739 ( .A(\U_0/U_0/U_1/STOP_DATA [0]), .Y(n10567) );
  INVX2 U10740 ( .A(\U_0/U_0/U_1/U_2/nextState[2] ), .Y(n10568) );
  INVX2 U10741 ( .A(n6619), .Y(n10569) );
  INVX2 U10742 ( .A(\U_0/U_0/U_1/U_2/nextState[1] ), .Y(n10570) );
  INVX2 U10743 ( .A(\U_0/U_0/U_1/U_2/timerRunning ), .Y(n10571) );
  INVX2 U10744 ( .A(\U_0/U_0/U_1/U_2/N99 ), .Y(n10572) );
  INVX2 U10745 ( .A(\U_0/U_0/U_1/U_2/state[1] ), .Y(n10573) );
  INVX2 U10746 ( .A(\U_0/U_0/U_1/U_2/state[2] ), .Y(n10574) );
  INVX2 U10747 ( .A(n744), .Y(n10575) );
  INVX2 U10748 ( .A(\U_0/U_0/U_1/CHK_ERROR ), .Y(n10576) );
  INVX2 U10749 ( .A(\U_0/U_0/U_1/SBC_CLR ), .Y(n10577) );
  INVX2 U10750 ( .A(\U_0/U_0/U_1/TIMER_TRIG ), .Y(n10578) );
  INVX2 U10751 ( .A(\U_0/U_0/U_1/U_7/nextState[0] ), .Y(n10579) );
  INVX2 U10752 ( .A(\U_0/U_0/U_1/U_7/nextState[1] ), .Y(n10580) );
  INVX2 U10753 ( .A(\U_0/U_0/U_1/U_7/state[1] ), .Y(n10581) );
  INVX2 U10754 ( .A(\U_0/U_0/U_1/U_7/nextState[2] ), .Y(n10582) );
  INVX2 U10755 ( .A(\U_0/U_0/U_1/U_7/state[2] ), .Y(n10583) );
  INVX2 U10756 ( .A(\U_0/U_0/U_1/U_7/nextState[3] ), .Y(n10584) );
  INVX2 U10757 ( .A(\U_0/U_0/U_1/U_7/nextState[4] ), .Y(n10585) );
  INVX2 U10758 ( .A(\U_0/U_0/U_1/U_7/state[4] ), .Y(n10586) );
  INVX2 U10759 ( .A(\U_0/U_0/U_1/SBC_EN ), .Y(n10587) );
  INVX2 U10760 ( .A(n5704), .Y(n10588) );
  INVX2 U10761 ( .A(\U_0/U_0/U_1/SBE ), .Y(n10589) );
  INVX2 U10762 ( .A(n5633), .Y(n10590) );
  INVX2 U10763 ( .A(n6782), .Y(n10591) );
  INVX2 U10764 ( .A(n6748), .Y(n10592) );
  INVX2 U10765 ( .A(n6795), .Y(n10593) );
  INVX2 U10766 ( .A(n5663), .Y(n10594) );
  INVX2 U10767 ( .A(n5728), .Y(n10595) );
  INVX2 U10768 ( .A(n5701), .Y(n10596) );
  INVX2 U10769 ( .A(\U_0/U_0/U_1/U_8/state[0] ), .Y(n10597) );
  INVX2 U10770 ( .A(n5684), .Y(n10598) );
  INVX2 U10771 ( .A(n5732), .Y(n10599) );
  INVX2 U10772 ( .A(n5724), .Y(n10600) );
  INVX2 U10773 ( .A(n5685), .Y(n10601) );
  INVX2 U10774 ( .A(n5723), .Y(n10602) );
  INVX2 U10775 ( .A(\U_0/U_0/U_1/U_8/keyCount[1] ), .Y(n10603) );
  INVX2 U10776 ( .A(\U_0/U_0/U_1/U_8/keyCount[2] ), .Y(n10604) );
  INVX2 U10777 ( .A(\U_0/U_0/U_1/U_8/state[2] ), .Y(n10605) );
  INVX2 U10778 ( .A(\U_0/U_0/U_1/U_8/keyCount[0] ), .Y(n10606) );
  INVX2 U10779 ( .A(\U_0/U_0/U_1/U_8/state[3] ), .Y(n10607) );
  INVX2 U10780 ( .A(\U_0/U_0/U_1/U_8/state[1] ), .Y(n10608) );
  INVX2 U10781 ( .A(\U_0/RBUF_FULL ), .Y(n10609) );
  INVX2 U10782 ( .A(\U_0/U_0/U_1/OE ), .Y(n10610) );
  INVX2 U10783 ( .A(n4828), .Y(n10611) );
  INVX2 U10784 ( .A(n4912), .Y(n10612) );
  INVX2 U10785 ( .A(n5031), .Y(n10613) );
  INVX2 U10786 ( .A(n5067), .Y(n10614) );
  INVX2 U10787 ( .A(n5146), .Y(n10615) );
  INVX2 U10788 ( .A(n5261), .Y(n10616) );
  INVX2 U10789 ( .A(n5297), .Y(n10617) );
  INVX2 U10790 ( .A(n5376), .Y(n10618) );
  INVX2 U10791 ( .A(n5491), .Y(n10619) );
  INVX2 U10792 ( .A(n5527), .Y(n10620) );
  INVX2 U10793 ( .A(n5610), .Y(n10621) );
  INVX2 U10794 ( .A(n5613), .Y(n10623) );
  INVX2 U10795 ( .A(n5412), .Y(n10624) );
  INVX2 U10796 ( .A(n5182), .Y(n10625) );
  INVX2 U10797 ( .A(n4952), .Y(n10626) );
  INVX2 U10798 ( .A(n4677), .Y(n10627) );
  INVX2 U10799 ( .A(n4717), .Y(n10628) );
  INVX2 U10800 ( .A(n4785), .Y(n10629) );
  INVX2 U10801 ( .A(n4859), .Y(n10630) );
  INVX2 U10802 ( .A(n4944), .Y(n10631) );
  INVX2 U10803 ( .A(n5059), .Y(n10632) );
  INVX2 U10804 ( .A(n5096), .Y(n10633) );
  INVX2 U10805 ( .A(n5174), .Y(n10634) );
  INVX2 U10806 ( .A(n5289), .Y(n10635) );
  INVX2 U10807 ( .A(n5326), .Y(n10636) );
  INVX2 U10808 ( .A(n5404), .Y(n10637) );
  INVX2 U10809 ( .A(n5519), .Y(n10638) );
  INVX2 U10810 ( .A(n5557), .Y(n10639) );
  INVX2 U10811 ( .A(n5641), .Y(n10640) );
  INVX2 U10812 ( .A(n5441), .Y(n10642) );
  INVX2 U10813 ( .A(n5211), .Y(n10643) );
  INVX2 U10814 ( .A(n4981), .Y(n10644) );
  INVX2 U10815 ( .A(n4670), .Y(n10645) );
  INVX2 U10816 ( .A(n4800), .Y(n10646) );
  INVX2 U10817 ( .A(n4757), .Y(n10647) );
  INVX2 U10818 ( .A(n4852), .Y(n10648) );
  INVX2 U10819 ( .A(n4975), .Y(n10649) );
  INVX2 U10820 ( .A(n5009), .Y(n10650) );
  INVX2 U10821 ( .A(n5090), .Y(n10651) );
  INVX2 U10822 ( .A(n5205), .Y(n10652) );
  INVX2 U10823 ( .A(n5239), .Y(n10653) );
  INVX2 U10824 ( .A(n5320), .Y(n10654) );
  INVX2 U10825 ( .A(n5435), .Y(n10655) );
  INVX2 U10826 ( .A(n5469), .Y(n10656) );
  INVX2 U10827 ( .A(n5550), .Y(n10657) );
  INVX2 U10828 ( .A(n5596), .Y(n10659) );
  INVX2 U10829 ( .A(n5354), .Y(n10660) );
  INVX2 U10830 ( .A(n5124), .Y(n10661) );
  INVX2 U10831 ( .A(n4889), .Y(n10662) );
  INVX2 U10832 ( .A(n4692), .Y(n10663) );
  INVX2 U10833 ( .A(n4794), .Y(n10664) );
  INVX2 U10834 ( .A(n4882), .Y(n10665) );
  INVX2 U10835 ( .A(n5003), .Y(n10666) );
  INVX2 U10836 ( .A(n5037), .Y(n10667) );
  INVX2 U10837 ( .A(n5118), .Y(n10668) );
  INVX2 U10838 ( .A(n5233), .Y(n10669) );
  INVX2 U10839 ( .A(n5267), .Y(n10670) );
  INVX2 U10840 ( .A(n5348), .Y(n10671) );
  INVX2 U10841 ( .A(n5463), .Y(n10672) );
  INVX2 U10842 ( .A(n5497), .Y(n10673) );
  INVX2 U10843 ( .A(n5579), .Y(n10674) );
  INVX2 U10844 ( .A(n5582), .Y(n10676) );
  INVX2 U10845 ( .A(n5382), .Y(n10677) );
  INVX2 U10846 ( .A(n5152), .Y(n10678) );
  INVX2 U10847 ( .A(n4919), .Y(n10679) );
  INVX2 U10848 ( .A(n4684), .Y(n10680) );
  INVX2 U10849 ( .A(\U_0/U_0/U_1/U_8/address[0] ), .Y(n10681) );
  INVX2 U10850 ( .A(n4844), .Y(n10682) );
  INVX2 U10851 ( .A(n4927), .Y(n10683) );
  INVX2 U10852 ( .A(n5045), .Y(n10684) );
  INVX2 U10853 ( .A(n5082), .Y(n10685) );
  INVX2 U10854 ( .A(n5160), .Y(n10686) );
  INVX2 U10855 ( .A(n5275), .Y(n10687) );
  INVX2 U10856 ( .A(n5312), .Y(n10688) );
  INVX2 U10857 ( .A(n5390), .Y(n10689) );
  INVX2 U10858 ( .A(n5505), .Y(n10690) );
  INVX2 U10859 ( .A(n5542), .Y(n10691) );
  INVX2 U10860 ( .A(n5623), .Y(n10692) );
  INVX2 U10861 ( .A(n5626), .Y(n10694) );
  INVX2 U10862 ( .A(n5427), .Y(n10695) );
  INVX2 U10863 ( .A(n5197), .Y(n10696) );
  INVX2 U10864 ( .A(n4967), .Y(n10697) );
  INVX2 U10865 ( .A(n4718), .Y(n10698) );
  INVX2 U10866 ( .A(n4836), .Y(n10699) );
  INVX2 U10867 ( .A(n4960), .Y(n10700) );
  INVX2 U10868 ( .A(n4995), .Y(n10701) );
  INVX2 U10869 ( .A(n5075), .Y(n10702) );
  INVX2 U10870 ( .A(n5190), .Y(n10703) );
  INVX2 U10871 ( .A(n5225), .Y(n10704) );
  INVX2 U10872 ( .A(n5305), .Y(n10705) );
  INVX2 U10873 ( .A(n5420), .Y(n10706) );
  INVX2 U10874 ( .A(n5455), .Y(n10707) );
  INVX2 U10875 ( .A(n5535), .Y(n10708) );
  INVX2 U10876 ( .A(n5571), .Y(n10710) );
  INVX2 U10877 ( .A(n5340), .Y(n10711) );
  INVX2 U10878 ( .A(n5110), .Y(n10712) );
  INVX2 U10879 ( .A(n4874), .Y(n10713) );
  INVX2 U10880 ( .A(n4695), .Y(n10714) );
  INVX2 U10881 ( .A(n4867), .Y(n10716) );
  INVX2 U10882 ( .A(n4989), .Y(n10717) );
  INVX2 U10883 ( .A(n5023), .Y(n10718) );
  INVX2 U10884 ( .A(n5104), .Y(n10719) );
  INVX2 U10885 ( .A(n5219), .Y(n10720) );
  INVX2 U10886 ( .A(n5253), .Y(n10721) );
  INVX2 U10887 ( .A(n5334), .Y(n10722) );
  INVX2 U10888 ( .A(n5449), .Y(n10723) );
  INVX2 U10889 ( .A(n5483), .Y(n10724) );
  INVX2 U10890 ( .A(n5565), .Y(n10725) );
  INVX2 U10891 ( .A(n5584), .Y(n10727) );
  INVX2 U10892 ( .A(n5368), .Y(n10728) );
  INVX2 U10893 ( .A(n5138), .Y(n10729) );
  INVX2 U10894 ( .A(n4904), .Y(n10730) );
  INVX2 U10895 ( .A(n4688), .Y(n10731) );
  INVX2 U10896 ( .A(n4731), .Y(n10732) );
  INVX2 U10897 ( .A(n4810), .Y(n10733) );
  INVX2 U10898 ( .A(n4897), .Y(n10734) );
  INVX2 U10899 ( .A(n5017), .Y(n10735) );
  INVX2 U10900 ( .A(n5051), .Y(n10736) );
  INVX2 U10901 ( .A(n5132), .Y(n10737) );
  INVX2 U10902 ( .A(n5247), .Y(n10738) );
  INVX2 U10903 ( .A(n5281), .Y(n10739) );
  INVX2 U10904 ( .A(n5362), .Y(n10740) );
  INVX2 U10905 ( .A(n5477), .Y(n10741) );
  INVX2 U10906 ( .A(n5511), .Y(n10742) );
  INVX2 U10907 ( .A(n5595), .Y(n10743) );
  INVX2 U10908 ( .A(n5599), .Y(n10745) );
  INVX2 U10909 ( .A(n5396), .Y(n10746) );
  INVX2 U10910 ( .A(n5166), .Y(n10747) );
  INVX2 U10911 ( .A(n4936), .Y(n10748) );
  INVX2 U10912 ( .A(n4682), .Y(n10749) );
  INVX2 U10913 ( .A(n4765), .Y(n10750) );
  INVX2 U10914 ( .A(\U_0/U_0/U_1/U_8/address[1] ), .Y(n10751) );
  INVX2 U10915 ( .A(\U_0/U_0/U_1/U_8/address[2] ), .Y(n10752) );
  INVX2 U10916 ( .A(\U_0/U_0/U_1/U_8/address[6] ), .Y(n10753) );
  INVX2 U10917 ( .A(n5642), .Y(n10754) );
  INVX2 U10918 ( .A(\U_0/U_0/U_1/U_8/address[7] ), .Y(n10755) );
  INVX2 U10919 ( .A(n4697), .Y(n10757) );
  INVX2 U10920 ( .A(\U_0/U_0/U_1/U_8/address[5] ), .Y(n10758) );
  INVX2 U10921 ( .A(\U_0/U_0/U_1/U_8/address[4] ), .Y(n10759) );
  INVX2 U10922 ( .A(\U_0/U_0/U_1/LOAD_DATA [7]), .Y(n10760) );
  INVX2 U10923 ( .A(\U_0/U_0/U_1/RCV_DATA [7]), .Y(n10761) );
  INVX2 U10924 ( .A(\U_0/U_0/U_1/LOAD_DATA [6]), .Y(n10762) );
  INVX2 U10925 ( .A(\U_0/U_0/U_1/LOAD_DATA [5]), .Y(n10763) );
  INVX2 U10926 ( .A(\U_0/U_0/U_1/RCV_DATA [5]), .Y(n10764) );
  INVX2 U10927 ( .A(\U_0/U_0/U_1/LOAD_DATA [4]), .Y(n10765) );
  INVX2 U10928 ( .A(\U_0/U_0/U_1/RCV_DATA [4]), .Y(n10766) );
  INVX2 U10929 ( .A(\U_0/U_0/U_1/LOAD_DATA [3]), .Y(n10767) );
  INVX2 U10930 ( .A(\U_0/U_0/U_1/RCV_DATA [3]), .Y(n10768) );
  INVX2 U10931 ( .A(\U_0/U_0/U_1/LOAD_DATA [2]), .Y(n10769) );
  INVX2 U10932 ( .A(\U_0/U_0/U_1/LOAD_DATA [1]), .Y(n10770) );
  INVX2 U10933 ( .A(\U_0/U_0/U_1/RCV_DATA [1]), .Y(n10771) );
  INVX2 U10934 ( .A(\U_0/U_0/U_1/LOAD_DATA [0]), .Y(n10772) );
  INVX2 U10935 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[0] ), .Y(n10773) );
  INVX2 U10936 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[1] ), .Y(n10774) );
  INVX2 U10937 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[2] ), .Y(n10775) );
  INVX2 U10938 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[3] ), .Y(n10776) );
  INVX2 U10939 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[4] ), .Y(n10777) );
  INVX2 U10940 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[5] ), .Y(n10778) );
  INVX2 U10941 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[6] ), .Y(n10779) );
  INVX2 U10942 ( .A(\U_0/U_0/U_1/U_8/parityAccumulator[7] ), .Y(n10780) );
  INVX2 U10943 ( .A(\U_0/U_0/U_1/U_8/parityError ), .Y(n10781) );
  INVX2 U10944 ( .A(\U_0/U_0/U_1/U_8/currentPlainKey[0] ), .Y(n10782) );
  INVX2 U10945 ( .A(\U_0/U_0/PLAINKEY [0]), .Y(n10783) );
  INVX2 U10946 ( .A(\U_0/U_0/U_1/U_8/currentPlainKey[1] ), .Y(n10784) );
  INVX2 U10947 ( .A(\U_0/U_0/PLAINKEY [1]), .Y(n10785) );
  INVX2 U10948 ( .A(\U_0/U_0/U_1/U_8/currentPlainKey[2] ), .Y(n10786) );
  INVX2 U10949 ( .A(\U_0/U_0/PLAINKEY [2]), .Y(n10787) );
  INVX2 U10950 ( .A(\U_0/U_0/U_1/U_8/currentPlainKey[3] ), .Y(n10788) );
  INVX2 U10951 ( .A(\U_0/U_0/PLAINKEY [3]), .Y(n10789) );
  INVX2 U10952 ( .A(\U_0/U_0/U_1/U_8/currentPlainKey[63] ), .Y(n10790) );
  INVX2 U10953 ( .A(\U_0/U_0/PLAINKEY [63]), .Y(n10791) );
  INVX2 U10954 ( .A(n6496), .Y(n10792) );
  INVX2 U10955 ( .A(n4417), .Y(n10793) );
  INVX2 U10956 ( .A(n6477), .Y(n10794) );
  INVX2 U10957 ( .A(n6572), .Y(n10795) );
  INVX2 U10958 ( .A(n4629), .Y(n10796) );
  INVX2 U10959 ( .A(n6512), .Y(n10797) );
  INVX2 U10960 ( .A(n6571), .Y(n10798) );
  INVX2 U10961 ( .A(n6511), .Y(n10799) );
  INVX2 U10962 ( .A(\U_0/U_2/U_5/state[0] ), .Y(n10800) );
  INVX2 U10963 ( .A(n6570), .Y(n10801) );
  INVX2 U10964 ( .A(n6515), .Y(n10802) );
  INVX2 U10965 ( .A(n4616), .Y(n10803) );
  INVX2 U10966 ( .A(n4611), .Y(n10804) );
  INVX2 U10967 ( .A(\U_0/U_2/U_5/state[3] ), .Y(n10806) );
  INVX2 U10968 ( .A(n6471), .Y(n10807) );
  INVX2 U10969 ( .A(\U_0/U_2/U_7/count[2] ), .Y(n10808) );
  INVX2 U10970 ( .A(n6493), .Y(BSE_H) );
  INVX2 U10971 ( .A(n760), .Y(n10810) );
  INVX2 U10972 ( .A(n4663), .Y(n10811) );
  INVX2 U10973 ( .A(\U_0/U_2/U_1/state[0] ), .Y(n10812) );
  INVX2 U10974 ( .A(n4656), .Y(n10813) );
  INVX2 U10975 ( .A(\U_0/U_2/U_1/DP_hold2 ), .Y(n10814) );
  INVX2 U10976 ( .A(\U_0/U_2/U_1/state[3] ), .Y(n10815) );
  INVX2 U10977 ( .A(\U_0/U_2/U_1/state[1] ), .Y(n10816) );
  INVX2 U10978 ( .A(n6517), .Y(n10817) );
  INVX2 U10979 ( .A(\U_0/U_2/U_5/N170 ), .Y(n10818) );
  INVX2 U10980 ( .A(\U_0/U_2/rx_CHECK_CRC [7]), .Y(n10819) );
  INVX2 U10981 ( .A(n4643), .Y(n10820) );
  INVX2 U10982 ( .A(\U_0/U_2/U_5/count[0] ), .Y(n10821) );
  INVX2 U10983 ( .A(\U_0/U_2/U_5/count[1] ), .Y(n10822) );
  INVX2 U10984 ( .A(\U_0/U_2/U_5/count[2] ), .Y(n10823) );
  INVX2 U10985 ( .A(\U_0/U_2/U_5/count[3] ), .Y(n10824) );
  INVX2 U10986 ( .A(\U_0/U_2/U_2/current_crc[15] ), .Y(n10826) );
  INVX2 U10987 ( .A(\U_0/U_2/U_2/current_crc[0] ), .Y(n10827) );
  INVX2 U10988 ( .A(\U_0/U_2/U_2/cache_1 [0]), .Y(n10828) );
  INVX2 U10989 ( .A(\U_0/U_2/U_2/current_crc[8] ), .Y(n10829) );
  INVX2 U10990 ( .A(\U_0/U_2/U_2/current_crc[2] ), .Y(n10830) );
  INVX2 U10991 ( .A(\U_0/U_2/U_2/cache_1 [2]), .Y(n10831) );
  INVX2 U10992 ( .A(\U_0/U_2/U_2/current_crc[10] ), .Y(n10832) );
  INVX2 U10993 ( .A(\U_0/U_2/U_2/current_crc[3] ), .Y(n10833) );
  INVX2 U10994 ( .A(\U_0/U_2/U_2/cache_1 [3]), .Y(n10834) );
  INVX2 U10995 ( .A(\U_0/U_2/U_2/current_crc[11] ), .Y(n10835) );
  INVX2 U10996 ( .A(\U_0/U_2/U_2/current_crc[4] ), .Y(n10836) );
  INVX2 U10997 ( .A(\U_0/U_2/U_2/cache_1 [4]), .Y(n10837) );
  INVX2 U10998 ( .A(\U_0/U_2/U_2/current_crc[12] ), .Y(n10838) );
  INVX2 U10999 ( .A(\U_0/U_2/U_2/cache_1 [12]), .Y(n10839) );
  INVX2 U11000 ( .A(\U_0/U_2/U_2/current_crc[5] ), .Y(n10840) );
  INVX2 U11001 ( .A(\U_0/U_2/U_2/cache_1 [5]), .Y(n10841) );
  INVX2 U11002 ( .A(\U_0/U_2/U_2/current_crc[13] ), .Y(n10842) );
  INVX2 U11003 ( .A(\U_0/U_2/U_2/current_crc[6] ), .Y(n10843) );
  INVX2 U11004 ( .A(\U_0/U_2/U_2/cache_1 [6]), .Y(n10844) );
  INVX2 U11005 ( .A(\U_0/U_2/U_2/current_crc[14] ), .Y(n10845) );
  INVX2 U11006 ( .A(\U_0/U_2/U_2/cache_1 [14]), .Y(n10846) );
  INVX2 U11007 ( .A(\U_0/U_2/U_2/current_crc[7] ), .Y(n10847) );
  INVX2 U11008 ( .A(\U_0/U_2/U_2/cache_1 [7]), .Y(n10848) );
  INVX2 U11009 ( .A(\U_0/U_2/U_2/cache_1 [13]), .Y(n10849) );
  INVX2 U11010 ( .A(\U_0/U_2/U_2/cache_1 [11]), .Y(n10850) );
  INVX2 U11011 ( .A(\U_0/U_2/U_2/current_crc[1] ), .Y(n10851) );
  INVX2 U11012 ( .A(\U_0/U_2/U_2/cache_1 [1]), .Y(n10852) );
  INVX2 U11013 ( .A(\U_0/U_2/U_2/current_crc[9] ), .Y(n10853) );
  INVX2 U11014 ( .A(\U_0/U_2/U_2/cache_1 [9]), .Y(n10854) );
  INVX2 U11015 ( .A(\U_0/U_2/U_2/cache_1 [10]), .Y(n10855) );
  INVX2 U11016 ( .A(\U_0/U_2/U_2/cache_1 [8]), .Y(n10856) );
  INVX2 U11017 ( .A(\U_0/U_2/U_2/cache_1 [15]), .Y(n10857) );
  INVX2 U11018 ( .A(\U_0/U_2/rx_CHECK_CRC [0]), .Y(n10858) );
  INVX2 U11019 ( .A(\U_0/U_2/rx_CHECK_CRC [2]), .Y(n10859) );
  INVX2 U11020 ( .A(\U_0/U_2/rx_CHECK_CRC [3]), .Y(n10860) );
  INVX2 U11021 ( .A(\U_0/U_2/rx_CHECK_CRC [4]), .Y(n10861) );
  INVX2 U11022 ( .A(\U_0/U_2/rx_CHECK_CRC [5]), .Y(n10862) );
  INVX2 U11023 ( .A(\U_0/U_2/rx_CHECK_CRC [6]), .Y(n10863) );
  INVX2 U11024 ( .A(\U_0/U_2/U_7/count[0] ), .Y(n10864) );
  INVX2 U11025 ( .A(\U_0/U_2/U_7/count[1] ), .Y(n10865) );
  INVX2 U11026 ( .A(\U_0/U_2/U_5/curR_ERROR ), .Y(n10866) );
  INVX2 U11027 ( .A(\U_0/U_2/U_5/curCRC_ERROR ), .Y(n10867) );
  INVX2 U11028 ( .A(n3303), .Y(n10868) );
  INVX2 U11029 ( .A(n6441), .Y(n10869) );
  INVX2 U11030 ( .A(n6445), .Y(n10870) );
  INVX2 U11031 ( .A(\U_0/U_3/U_0/N59 ), .Y(n10871) );
  INVX2 U11032 ( .A(n9243), .Y(n10872) );
  INVX2 U11033 ( .A(n3334), .Y(n10873) );
  INVX2 U11034 ( .A(n3308), .Y(n10874) );
  INVX2 U11035 ( .A(\U_0/U_3/U_0/state[3] ), .Y(n10875) );
  INVX2 U11036 ( .A(n6413), .Y(n10876) );
  INVX2 U11037 ( .A(n6420), .Y(n10877) );
  INVX2 U11038 ( .A(n6424), .Y(n10878) );
  INVX2 U11039 ( .A(\U_0/U_3/U_0/DE_holdout ), .Y(n10879) );
  INVX2 U11040 ( .A(\U_0/U_3/U_0/DE_holdout_last ), .Y(n10880) );
  INVX2 U11041 ( .A(n3307), .Y(n10881) );
  INVX2 U11042 ( .A(n6432), .Y(n10882) );
  INVX2 U11043 ( .A(n6418), .Y(n10883) );
  INVX2 U11044 ( .A(n6446), .Y(n10884) );
  INVX2 U11045 ( .A(\U_0/U_3/U_0/state[2] ), .Y(n10885) );
  INVX2 U11046 ( .A(\U_0/U_3/U_0/state[0] ), .Y(n10886) );
  INVX2 U11047 ( .A(\U_0/U_3/U_0/state[1] ), .Y(n10887) );
  INVX2 U11048 ( .A(host_is_sending), .Y(n10888) );
  INVX2 U11049 ( .A(n3312), .Y(n10889) );
  INVX2 U11050 ( .A(n6379), .Y(n10890) );
  INVX2 U11051 ( .A(n6460), .Y(n10891) );
  INVX2 U11052 ( .A(n6380), .Y(n10892) );
  INVX2 U11053 ( .A(n3384), .Y(n10893) );
  INVX2 U11054 ( .A(n4501), .Y(n10894) );
  INVX2 U11055 ( .A(n6389), .Y(n10895) );
  INVX2 U11056 ( .A(n3387), .Y(n10896) );
  INVX2 U11057 ( .A(n518), .Y(n10897) );
  INVX2 U11058 ( .A(n3400), .Y(n10898) );
  INVX2 U11059 ( .A(n6582), .Y(n10899) );
  INVX2 U11060 ( .A(n3398), .Y(n10900) );
  INVX2 U11061 ( .A(\U_0/U_3/U_3/state[1] ), .Y(n10901) );
  INVX2 U11062 ( .A(n6385), .Y(n10902) );
  INVX2 U11063 ( .A(\U_0/U_3/U_3/state[2] ), .Y(n10903) );
  INVX2 U11064 ( .A(\U_0/U_3/U_3/state[0] ), .Y(n10904) );
  INVX2 U11065 ( .A(\U_0/U_1/U_0/state[2] ), .Y(n10905) );
  INVX2 U11066 ( .A(n6591), .Y(n10906) );
  INVX2 U11067 ( .A(n6596), .Y(n10907) );
  INVX2 U11068 ( .A(\U_0/U_1/R_ENABLE ), .Y(n10908) );
  INVX2 U11069 ( .A(n4116), .Y(n10909) );
  INVX2 U11070 ( .A(n4131), .Y(n10910) );
  INVX2 U11071 ( .A(n4147), .Y(n10911) );
  INVX2 U11072 ( .A(n4160), .Y(n10912) );
  INVX2 U11073 ( .A(n4115), .Y(n10913) );
  INVX2 U11074 ( .A(n4129), .Y(n10914) );
  INVX2 U11075 ( .A(n4145), .Y(n10915) );
  INVX2 U11076 ( .A(n4161), .Y(n10916) );
  INVX2 U11077 ( .A(\U_0/U_1/U_1/writeptr[0] ), .Y(n10917) );
  INVX2 U11078 ( .A(\U_0/U_1/U_1/opcode[4][0] ), .Y(n10918) );
  INVX2 U11079 ( .A(\U_0/U_1/U_1/opcode[4][1] ), .Y(n10919) );
  INVX2 U11080 ( .A(\U_0/U_1/U_1/memory[4][0] ), .Y(n10920) );
  INVX2 U11081 ( .A(\U_0/U_1/U_1/memory[4][1] ), .Y(n10921) );
  INVX2 U11082 ( .A(\U_0/U_1/U_1/memory[4][2] ), .Y(n10922) );
  INVX2 U11083 ( .A(\U_0/U_1/U_1/memory[4][3] ), .Y(n10923) );
  INVX2 U11084 ( .A(\U_0/U_1/U_1/memory[4][4] ), .Y(n10924) );
  INVX2 U11085 ( .A(\U_0/U_1/U_1/memory[4][5] ), .Y(n10925) );
  INVX2 U11086 ( .A(\U_0/U_1/U_1/memory[4][6] ), .Y(n10926) );
  INVX2 U11087 ( .A(\U_0/U_1/U_1/memory[4][7] ), .Y(n10927) );
  INVX2 U11088 ( .A(\U_0/U_1/U_1/opcode[5][0] ), .Y(n10928) );
  INVX2 U11089 ( .A(\U_0/U_1/U_1/opcode[5][1] ), .Y(n10929) );
  INVX2 U11090 ( .A(\U_0/U_1/U_1/memory[5][0] ), .Y(n10930) );
  INVX2 U11091 ( .A(\U_0/U_1/U_1/memory[5][1] ), .Y(n10931) );
  INVX2 U11092 ( .A(\U_0/U_1/U_1/memory[5][2] ), .Y(n10932) );
  INVX2 U11093 ( .A(\U_0/U_1/U_1/memory[5][3] ), .Y(n10933) );
  INVX2 U11094 ( .A(\U_0/U_1/U_1/memory[5][4] ), .Y(n10934) );
  INVX2 U11095 ( .A(\U_0/U_1/U_1/memory[5][5] ), .Y(n10935) );
  INVX2 U11096 ( .A(\U_0/U_1/U_1/memory[5][6] ), .Y(n10936) );
  INVX2 U11097 ( .A(\U_0/U_1/U_1/memory[5][7] ), .Y(n10937) );
  INVX2 U11098 ( .A(\U_0/U_1/U_1/memory[6][0] ), .Y(n10938) );
  INVX2 U11099 ( .A(\U_0/U_1/U_1/memory[6][1] ), .Y(n10939) );
  INVX2 U11100 ( .A(\U_0/U_1/U_1/memory[6][2] ), .Y(n10940) );
  INVX2 U11101 ( .A(\U_0/U_1/U_1/memory[6][3] ), .Y(n10941) );
  INVX2 U11102 ( .A(\U_0/U_1/U_1/memory[6][4] ), .Y(n10942) );
  INVX2 U11103 ( .A(\U_0/U_1/U_1/memory[6][5] ), .Y(n10943) );
  INVX2 U11104 ( .A(\U_0/U_1/U_1/memory[6][6] ), .Y(n10944) );
  INVX2 U11105 ( .A(\U_0/U_1/U_1/memory[6][7] ), .Y(n10945) );
  INVX2 U11106 ( .A(\U_0/U_1/U_1/memory[7][6] ), .Y(n10946) );
  INVX2 U11107 ( .A(\U_0/U_1/U_1/memory[7][7] ), .Y(n10947) );
  INVX2 U11108 ( .A(\U_0/U_1/U_1/memory[7][0] ), .Y(n10948) );
  INVX2 U11109 ( .A(\U_0/U_1/U_1/memory[7][1] ), .Y(n10949) );
  INVX2 U11110 ( .A(\U_0/U_1/U_1/memory[7][2] ), .Y(n10950) );
  INVX2 U11111 ( .A(\U_0/U_1/U_1/memory[7][3] ), .Y(n10951) );
  INVX2 U11112 ( .A(\U_0/U_1/U_1/memory[7][4] ), .Y(n10952) );
  INVX2 U11113 ( .A(\U_0/U_1/U_1/memory[7][5] ), .Y(n10953) );
  INVX2 U11114 ( .A(\U_0/U_1/U_1/opcode[11][1] ), .Y(n10954) );
  INVX2 U11115 ( .A(\U_0/U_1/U_1/opcode[11][0] ), .Y(n10955) );
  INVX2 U11116 ( .A(\U_0/U_1/U_1/opcode[6][0] ), .Y(n10956) );
  INVX2 U11117 ( .A(\U_0/U_1/U_1/opcode[6][1] ), .Y(n10957) );
  INVX2 U11118 ( .A(\U_0/U_1/U_1/opcode[7][0] ), .Y(n10958) );
  INVX2 U11119 ( .A(\U_0/U_1/U_1/opcode[7][1] ), .Y(n10959) );
  INVX2 U11120 ( .A(\U_0/U_1/U_1/memory[11][0] ), .Y(n10960) );
  INVX2 U11121 ( .A(\U_0/U_1/U_1/memory[11][1] ), .Y(n10961) );
  INVX2 U11122 ( .A(\U_0/U_1/U_1/memory[11][2] ), .Y(n10962) );
  INVX2 U11123 ( .A(\U_0/U_1/U_1/memory[11][3] ), .Y(n10963) );
  INVX2 U11124 ( .A(\U_0/U_1/U_1/memory[11][4] ), .Y(n10964) );
  INVX2 U11125 ( .A(\U_0/U_1/U_1/memory[11][5] ), .Y(n10965) );
  INVX2 U11126 ( .A(\U_0/U_1/U_1/memory[11][6] ), .Y(n10966) );
  INVX2 U11127 ( .A(\U_0/U_1/U_1/memory[11][7] ), .Y(n10967) );
  INVX2 U11128 ( .A(\U_0/U_1/U_1/opcode[8][0] ), .Y(n10968) );
  INVX2 U11129 ( .A(\U_0/U_1/U_1/opcode[8][1] ), .Y(n10969) );
  INVX2 U11130 ( .A(\U_0/U_1/U_1/memory[8][0] ), .Y(n10970) );
  INVX2 U11131 ( .A(\U_0/U_1/U_1/memory[8][1] ), .Y(n10971) );
  INVX2 U11132 ( .A(\U_0/U_1/U_1/memory[8][2] ), .Y(n10972) );
  INVX2 U11133 ( .A(\U_0/U_1/U_1/memory[8][3] ), .Y(n10973) );
  INVX2 U11134 ( .A(\U_0/U_1/U_1/memory[8][4] ), .Y(n10974) );
  INVX2 U11135 ( .A(\U_0/U_1/U_1/memory[8][5] ), .Y(n10975) );
  INVX2 U11136 ( .A(\U_0/U_1/U_1/memory[8][6] ), .Y(n10976) );
  INVX2 U11137 ( .A(\U_0/U_1/U_1/memory[8][7] ), .Y(n10977) );
  INVX2 U11138 ( .A(\U_0/U_1/U_1/opcode[9][0] ), .Y(n10978) );
  INVX2 U11139 ( .A(\U_0/U_1/U_1/opcode[9][1] ), .Y(n10979) );
  INVX2 U11140 ( .A(\U_0/U_1/U_1/memory[9][0] ), .Y(n10980) );
  INVX2 U11141 ( .A(\U_0/U_1/U_1/memory[9][1] ), .Y(n10981) );
  INVX2 U11142 ( .A(\U_0/U_1/U_1/memory[9][2] ), .Y(n10982) );
  INVX2 U11143 ( .A(\U_0/U_1/U_1/memory[9][3] ), .Y(n10983) );
  INVX2 U11144 ( .A(\U_0/U_1/U_1/memory[9][4] ), .Y(n10984) );
  INVX2 U11145 ( .A(\U_0/U_1/U_1/memory[9][5] ), .Y(n10985) );
  INVX2 U11146 ( .A(\U_0/U_1/U_1/memory[9][6] ), .Y(n10986) );
  INVX2 U11147 ( .A(\U_0/U_1/U_1/memory[9][7] ), .Y(n10987) );
  INVX2 U11148 ( .A(\U_0/U_1/U_1/opcode[10][0] ), .Y(n10988) );
  INVX2 U11149 ( .A(\U_0/U_1/U_1/opcode[10][1] ), .Y(n10989) );
  INVX2 U11150 ( .A(\U_0/U_1/U_1/memory[10][0] ), .Y(n10990) );
  INVX2 U11151 ( .A(\U_0/U_1/U_1/memory[10][1] ), .Y(n10991) );
  INVX2 U11152 ( .A(\U_0/U_1/U_1/memory[10][2] ), .Y(n10992) );
  INVX2 U11153 ( .A(\U_0/U_1/U_1/memory[10][3] ), .Y(n10993) );
  INVX2 U11154 ( .A(\U_0/U_1/U_1/memory[10][4] ), .Y(n10994) );
  INVX2 U11155 ( .A(\U_0/U_1/U_1/memory[10][5] ), .Y(n10995) );
  INVX2 U11156 ( .A(\U_0/U_1/U_1/memory[10][6] ), .Y(n10996) );
  INVX2 U11157 ( .A(\U_0/U_1/U_1/memory[10][7] ), .Y(n10997) );
  INVX2 U11158 ( .A(\U_0/U_1/U_1/opcode[28][0] ), .Y(n10998) );
  INVX2 U11159 ( .A(\U_0/U_1/U_1/opcode[28][1] ), .Y(n10999) );
  INVX2 U11160 ( .A(\U_0/U_1/U_1/memory[28][0] ), .Y(n11000) );
  INVX2 U11161 ( .A(\U_0/U_1/U_1/memory[28][1] ), .Y(n11001) );
  INVX2 U11162 ( .A(\U_0/U_1/U_1/memory[28][2] ), .Y(n11002) );
  INVX2 U11163 ( .A(\U_0/U_1/U_1/memory[28][3] ), .Y(n11003) );
  INVX2 U11164 ( .A(\U_0/U_1/U_1/memory[28][4] ), .Y(n11004) );
  INVX2 U11165 ( .A(\U_0/U_1/U_1/memory[28][5] ), .Y(n11005) );
  INVX2 U11166 ( .A(\U_0/U_1/U_1/memory[28][6] ), .Y(n11006) );
  INVX2 U11167 ( .A(\U_0/U_1/U_1/memory[28][7] ), .Y(n11007) );
  INVX2 U11168 ( .A(\U_0/U_1/U_1/opcode[29][0] ), .Y(n11008) );
  INVX2 U11169 ( .A(\U_0/U_1/U_1/opcode[29][1] ), .Y(n11009) );
  INVX2 U11170 ( .A(\U_0/U_1/U_1/memory[29][0] ), .Y(n11010) );
  INVX2 U11171 ( .A(\U_0/U_1/U_1/memory[29][1] ), .Y(n11011) );
  INVX2 U11172 ( .A(\U_0/U_1/U_1/memory[29][2] ), .Y(n11012) );
  INVX2 U11173 ( .A(\U_0/U_1/U_1/memory[29][3] ), .Y(n11013) );
  INVX2 U11174 ( .A(\U_0/U_1/U_1/memory[29][4] ), .Y(n11014) );
  INVX2 U11175 ( .A(\U_0/U_1/U_1/memory[29][5] ), .Y(n11015) );
  INVX2 U11176 ( .A(\U_0/U_1/U_1/memory[29][6] ), .Y(n11016) );
  INVX2 U11177 ( .A(\U_0/U_1/U_1/memory[29][7] ), .Y(n11017) );
  INVX2 U11178 ( .A(\U_0/U_1/U_1/opcode[30][0] ), .Y(n11018) );
  INVX2 U11179 ( .A(\U_0/U_1/U_1/opcode[30][1] ), .Y(n11019) );
  INVX2 U11180 ( .A(\U_0/U_1/U_1/memory[30][0] ), .Y(n11020) );
  INVX2 U11181 ( .A(\U_0/U_1/U_1/memory[30][1] ), .Y(n11021) );
  INVX2 U11182 ( .A(\U_0/U_1/U_1/memory[30][2] ), .Y(n11022) );
  INVX2 U11183 ( .A(\U_0/U_1/U_1/memory[30][3] ), .Y(n11023) );
  INVX2 U11184 ( .A(\U_0/U_1/U_1/memory[30][4] ), .Y(n11024) );
  INVX2 U11185 ( .A(\U_0/U_1/U_1/memory[30][5] ), .Y(n11025) );
  INVX2 U11186 ( .A(\U_0/U_1/U_1/memory[30][6] ), .Y(n11026) );
  INVX2 U11187 ( .A(\U_0/U_1/U_1/memory[30][7] ), .Y(n11027) );
  INVX2 U11188 ( .A(\U_0/U_1/U_1/opcode[31][0] ), .Y(n11028) );
  INVX2 U11189 ( .A(\U_0/U_1/U_1/opcode[31][1] ), .Y(n11029) );
  INVX2 U11190 ( .A(\U_0/U_1/U_1/memory[31][0] ), .Y(n11030) );
  INVX2 U11191 ( .A(\U_0/U_1/U_1/memory[31][1] ), .Y(n11031) );
  INVX2 U11192 ( .A(\U_0/U_1/U_1/memory[31][2] ), .Y(n11032) );
  INVX2 U11193 ( .A(\U_0/U_1/U_1/memory[31][3] ), .Y(n11033) );
  INVX2 U11194 ( .A(\U_0/U_1/U_1/memory[31][4] ), .Y(n11034) );
  INVX2 U11195 ( .A(\U_0/U_1/U_1/memory[31][5] ), .Y(n11035) );
  INVX2 U11196 ( .A(\U_0/U_1/U_1/memory[31][6] ), .Y(n11036) );
  INVX2 U11197 ( .A(\U_0/U_1/U_1/memory[31][7] ), .Y(n11037) );
  INVX2 U11198 ( .A(\U_0/U_1/U_1/opcode[16][0] ), .Y(n11038) );
  INVX2 U11199 ( .A(\U_0/U_1/U_1/opcode[16][1] ), .Y(n11039) );
  INVX2 U11200 ( .A(\U_0/U_1/U_1/memory[16][0] ), .Y(n11040) );
  INVX2 U11201 ( .A(\U_0/U_1/U_1/memory[16][1] ), .Y(n11041) );
  INVX2 U11202 ( .A(\U_0/U_1/U_1/memory[16][2] ), .Y(n11042) );
  INVX2 U11203 ( .A(\U_0/U_1/U_1/memory[16][3] ), .Y(n11043) );
  INVX2 U11204 ( .A(\U_0/U_1/U_1/memory[16][4] ), .Y(n11044) );
  INVX2 U11205 ( .A(\U_0/U_1/U_1/memory[16][5] ), .Y(n11045) );
  INVX2 U11206 ( .A(\U_0/U_1/U_1/memory[16][6] ), .Y(n11046) );
  INVX2 U11207 ( .A(\U_0/U_1/U_1/memory[16][7] ), .Y(n11047) );
  INVX2 U11208 ( .A(\U_0/U_1/U_1/opcode[17][0] ), .Y(n11048) );
  INVX2 U11209 ( .A(\U_0/U_1/U_1/opcode[17][1] ), .Y(n11049) );
  INVX2 U11210 ( .A(\U_0/U_1/U_1/memory[17][0] ), .Y(n11050) );
  INVX2 U11211 ( .A(\U_0/U_1/U_1/memory[17][1] ), .Y(n11051) );
  INVX2 U11212 ( .A(\U_0/U_1/U_1/memory[17][2] ), .Y(n11052) );
  INVX2 U11213 ( .A(\U_0/U_1/U_1/memory[17][3] ), .Y(n11053) );
  INVX2 U11214 ( .A(\U_0/U_1/U_1/memory[17][4] ), .Y(n11054) );
  INVX2 U11215 ( .A(\U_0/U_1/U_1/memory[17][5] ), .Y(n11055) );
  INVX2 U11216 ( .A(\U_0/U_1/U_1/memory[17][6] ), .Y(n11056) );
  INVX2 U11217 ( .A(\U_0/U_1/U_1/memory[17][7] ), .Y(n11057) );
  INVX2 U11218 ( .A(\U_0/U_1/U_1/opcode[18][0] ), .Y(n11058) );
  INVX2 U11219 ( .A(\U_0/U_1/U_1/opcode[18][1] ), .Y(n11059) );
  INVX2 U11220 ( .A(\U_0/U_1/U_1/memory[18][0] ), .Y(n11060) );
  INVX2 U11221 ( .A(\U_0/U_1/U_1/memory[18][1] ), .Y(n11061) );
  INVX2 U11222 ( .A(\U_0/U_1/U_1/memory[18][2] ), .Y(n11062) );
  INVX2 U11223 ( .A(\U_0/U_1/U_1/memory[18][3] ), .Y(n11063) );
  INVX2 U11224 ( .A(\U_0/U_1/U_1/memory[18][4] ), .Y(n11064) );
  INVX2 U11225 ( .A(\U_0/U_1/U_1/memory[18][5] ), .Y(n11065) );
  INVX2 U11226 ( .A(\U_0/U_1/U_1/memory[18][6] ), .Y(n11066) );
  INVX2 U11227 ( .A(\U_0/U_1/U_1/memory[18][7] ), .Y(n11067) );
  INVX2 U11228 ( .A(\U_0/U_1/U_1/opcode[19][0] ), .Y(n11068) );
  INVX2 U11229 ( .A(\U_0/U_1/U_1/opcode[19][1] ), .Y(n11069) );
  INVX2 U11230 ( .A(\U_0/U_1/U_1/memory[19][3] ), .Y(n11070) );
  INVX2 U11231 ( .A(\U_0/U_1/U_1/memory[19][4] ), .Y(n11071) );
  INVX2 U11232 ( .A(\U_0/U_1/U_1/memory[19][5] ), .Y(n11072) );
  INVX2 U11233 ( .A(\U_0/U_1/U_1/memory[19][6] ), .Y(n11073) );
  INVX2 U11234 ( .A(\U_0/U_1/U_1/memory[19][7] ), .Y(n11074) );
  INVX2 U11235 ( .A(\U_0/U_1/U_1/memory[19][0] ), .Y(n11075) );
  INVX2 U11236 ( .A(\U_0/U_1/U_1/memory[19][1] ), .Y(n11076) );
  INVX2 U11237 ( .A(\U_0/U_1/U_1/memory[19][2] ), .Y(n11077) );
  INVX2 U11238 ( .A(n6592), .Y(n11078) );
  INVX2 U11239 ( .A(\U_0/U_1/DATA [0]), .Y(n11079) );
  INVX2 U11240 ( .A(\U_0/U_1/DATA [1]), .Y(n11080) );
  INVX2 U11241 ( .A(\U_0/U_1/DATA [2]), .Y(n11081) );
  INVX2 U11242 ( .A(\U_0/U_1/DATA [3]), .Y(n11082) );
  INVX2 U11243 ( .A(\U_0/U_1/DATA [4]), .Y(n11083) );
  INVX2 U11244 ( .A(\U_0/U_1/DATA [5]), .Y(n11084) );
  INVX2 U11245 ( .A(\U_0/U_1/DATA [6]), .Y(n11085) );
  INVX2 U11246 ( .A(\U_0/U_1/DATA [7]), .Y(n11086) );
  INVX2 U11247 ( .A(\U_0/U_1/OUT_OPCODE [0]), .Y(n11087) );
  INVX2 U11248 ( .A(\U_0/U_1/OUT_OPCODE [1]), .Y(n11088) );
  INVX2 U11249 ( .A(n6585), .Y(n11089) );
  INVX2 U11250 ( .A(\U_0/U_1/U_0/state[0] ), .Y(n11090) );
  INVX2 U11251 ( .A(\U_0/U_1/U_0/state[1] ), .Y(n11091) );
  INVX2 U11252 ( .A(\U_0/B_READY ), .Y(n11092) );
  INVX2 U11253 ( .A(n6383), .Y(n11093) );
  INVX2 U11254 ( .A(n6775), .Y(n11094) );
  INVX2 U11255 ( .A(\U_0/PRGA_OPCODE[0] ), .Y(n11095) );
  INVX2 U11256 ( .A(\U_0/U_1/U_0/tempOpcode [0]), .Y(n11096) );
  INVX2 U11257 ( .A(\U_0/U_1/U_0/tempData [7]), .Y(n11097) );
  INVX2 U11258 ( .A(\U_0/PRGA_IN [7]), .Y(n11098) );
  INVX2 U11259 ( .A(\U_0/U_1/U_0/tempData [6]), .Y(n11099) );
  INVX2 U11260 ( .A(\U_0/PRGA_IN [6]), .Y(n11100) );
  INVX2 U11261 ( .A(\U_0/U_1/U_0/tempData [5]), .Y(n11101) );
  INVX2 U11262 ( .A(\U_0/PRGA_IN [5]), .Y(n11102) );
  INVX2 U11263 ( .A(\U_0/U_1/U_0/tempData [4]), .Y(n11103) );
  INVX2 U11264 ( .A(\U_0/PRGA_IN [4]), .Y(n11104) );
  INVX2 U11265 ( .A(\U_0/U_1/U_0/tempData [3]), .Y(n11105) );
  INVX2 U11266 ( .A(\U_0/PRGA_IN [3]), .Y(n11106) );
  INVX2 U11267 ( .A(\U_0/U_1/U_0/tempData [2]), .Y(n11107) );
  INVX2 U11268 ( .A(\U_0/PRGA_IN [2]), .Y(n11108) );
  INVX2 U11269 ( .A(\U_0/U_1/U_0/tempData [1]), .Y(n11109) );
  INVX2 U11270 ( .A(\U_0/PRGA_IN [1]), .Y(n11110) );
  INVX2 U11271 ( .A(\U_0/U_1/U_0/tempData [0]), .Y(n11111) );
  INVX2 U11272 ( .A(\U_0/PRGA_IN [0]), .Y(n11112) );
  INVX2 U11273 ( .A(\U_0/PRGA_OPCODE[1] ), .Y(n11113) );
  INVX2 U11274 ( .A(\U_0/U_3/U_3/count[0] ), .Y(n11114) );
  INVX2 U11275 ( .A(\U_0/U_3/U_3/count[5] ), .Y(n11115) );
  INVX2 U11276 ( .A(n6402), .Y(n11116) );
  INVX2 U11277 ( .A(\U_0/U_3/U_3/count[1] ), .Y(n11117) );
  INVX2 U11278 ( .A(\U_0/U_3/U_3/count[2] ), .Y(n11118) );
  INVX2 U11279 ( .A(\U_0/U_3/U_3/count[3] ), .Y(n11119) );
  INVX2 U11280 ( .A(\U_0/U_3/U_3/count[4] ), .Y(n11120) );
  INVX2 U11281 ( .A(\U_0/U_0/U_0/nfaddr[0] ), .Y(n11121) );
  INVX2 U11282 ( .A(\U_0/U_0/U_0/nfaddr[1] ), .Y(n11122) );
  INVX2 U11283 ( .A(\U_0/U_0/U_0/nfaddr[2] ), .Y(n11123) );
  INVX2 U11284 ( .A(\U_0/U_0/U_0/nfaddr[3] ), .Y(n11124) );
  INVX2 U11285 ( .A(\U_0/U_0/U_0/nfaddr[4] ), .Y(n11125) );
  INVX2 U11286 ( .A(\U_0/U_0/U_0/nfaddr[5] ), .Y(n11126) );
  INVX2 U11287 ( .A(\U_0/U_0/U_0/nfaddr[6] ), .Y(n11127) );
  INVX2 U11288 ( .A(\U_0/U_0/U_0/nfaddr[7] ), .Y(n11128) );
  INVX2 U11289 ( .A(n6654), .Y(n11129) );
  INVX2 U11290 ( .A(n6658), .Y(n11130) );
  INVX2 U11291 ( .A(n3481), .Y(n11131) );
  INVX2 U11292 ( .A(n6763), .Y(n11132) );
  INVX2 U11293 ( .A(n3496), .Y(n11133) );
  INVX2 U11294 ( .A(n557), .Y(n11135) );
  INVX2 U11295 ( .A(n6676), .Y(n11136) );
  INVX2 U11296 ( .A(n3569), .Y(n11137) );
  INVX2 U11297 ( .A(n3502), .Y(n11138) );
  INVX2 U11298 ( .A(n3566), .Y(n11139) );
  INVX2 U11299 ( .A(n602), .Y(n11140) );
  INVX2 U11300 ( .A(n3563), .Y(n11141) );
  INVX2 U11301 ( .A(n3585), .Y(n11142) );
  INVX2 U11302 ( .A(n3501), .Y(n11143) );
  INVX2 U11303 ( .A(n6625), .Y(n11145) );
  INVX2 U11304 ( .A(n3674), .Y(n11146) );
  INVX2 U11305 ( .A(n3672), .Y(n11147) );
  INVX2 U11306 ( .A(n3438), .Y(n11148) );
  INVX2 U11307 ( .A(n6717), .Y(n11149) );
  INVX2 U11308 ( .A(n6753), .Y(n11150) );
  INVX2 U11309 ( .A(n3571), .Y(n11151) );
  INVX2 U11310 ( .A(n6742), .Y(n11152) );
  INVX2 U11311 ( .A(n3673), .Y(n11153) );
  INVX2 U11312 ( .A(n6837), .Y(n11154) );
  INVX2 U11313 ( .A(\U_0/U_0/U_0/state[0] ), .Y(n11156) );
  INVX2 U11314 ( .A(n6762), .Y(n11157) );
  INVX2 U11315 ( .A(n3655), .Y(n11158) );
  INVX2 U11316 ( .A(n6671), .Y(n11159) );
  INVX2 U11317 ( .A(n9188), .Y(n11160) );
  INVX2 U11318 ( .A(n6842), .Y(n11161) );
  INVX2 U11319 ( .A(n3669), .Y(n11162) );
  INVX2 U11320 ( .A(n567), .Y(n11163) );
  INVX2 U11321 ( .A(n6751), .Y(n11164) );
  INVX2 U11322 ( .A(n6833), .Y(n11165) );
  INVX2 U11323 ( .A(n6661), .Y(n11166) );
  INVX2 U11324 ( .A(\U_0/U_0/U_0/state[3] ), .Y(n11167) );
  INVX2 U11325 ( .A(n6664), .Y(n11168) );
  INVX2 U11326 ( .A(n3670), .Y(n11169) );
  INVX2 U11327 ( .A(n6764), .Y(n11170) );
  INVX2 U11328 ( .A(n9320), .Y(n11171) );
  INVX2 U11329 ( .A(\U_0/U_0/U_0/prefillCounter[7] ), .Y(n11172) );
  INVX2 U11330 ( .A(\U_0/U_0/U_0/state[1] ), .Y(n11173) );
  INVX2 U11331 ( .A(\U_0/U_0/U_0/prefillCounter[0] ), .Y(n11174) );
  INVX2 U11332 ( .A(\U_0/U_0/U_0/prefillCounter[1] ), .Y(n11175) );
  INVX2 U11333 ( .A(\U_0/U_0/U_0/prefillCounter[2] ), .Y(n11176) );
  INVX2 U11334 ( .A(\U_0/U_0/U_0/prefillCounter[3] ), .Y(n11177) );
  INVX2 U11335 ( .A(\U_0/U_0/U_0/prefillCounter[4] ), .Y(n11178) );
  INVX2 U11336 ( .A(\U_0/U_0/U_0/prefillCounter[5] ), .Y(n11179) );
  INVX2 U11337 ( .A(\U_0/U_0/U_0/prefillCounter[6] ), .Y(n11180) );
  INVX2 U11338 ( .A(\U_0/PDATA_READY ), .Y(n11181) );
  INVX2 U11339 ( .A(\U_0/U_0/U_0/intj[7] ), .Y(n11182) );
  INVX2 U11340 ( .A(\U_0/U_0/U_0/intj[0] ), .Y(n11183) );
  INVX2 U11341 ( .A(\U_0/U_0/U_0/intj[1] ), .Y(n11184) );
  INVX2 U11342 ( .A(\U_0/U_0/U_0/intj[2] ), .Y(n11185) );
  INVX2 U11343 ( .A(\U_0/U_0/U_0/intj[3] ), .Y(n11186) );
  INVX2 U11344 ( .A(\U_0/U_0/U_0/intj[4] ), .Y(n11187) );
  INVX2 U11345 ( .A(\U_0/U_0/U_0/intj[5] ), .Y(n11188) );
  INVX2 U11346 ( .A(\U_0/U_0/U_0/intj[6] ), .Y(n11189) );
  INVX2 U11347 ( .A(\U_0/U_0/U_0/sj[7] ), .Y(n11190) );
  INVX2 U11348 ( .A(\U_0/U_0/U_0/sj[6] ), .Y(n11191) );
  INVX2 U11349 ( .A(\U_0/U_0/U_0/sj[5] ), .Y(n11192) );
  INVX2 U11350 ( .A(\U_0/U_0/U_0/sj[4] ), .Y(n11193) );
  INVX2 U11351 ( .A(\U_0/U_0/U_0/sj[3] ), .Y(n11194) );
  INVX2 U11352 ( .A(\U_0/U_0/U_0/sj[2] ), .Y(n11195) );
  INVX2 U11353 ( .A(\U_0/U_0/U_0/sj[1] ), .Y(n11196) );
  INVX2 U11354 ( .A(\U_0/U_0/U_0/sj[0] ), .Y(n11197) );
  INVX2 U11355 ( .A(\U_0/U_0/U_0/temp[6] ), .Y(n11198) );
  INVX2 U11356 ( .A(\U_0/U_0/U_0/temp[0] ), .Y(n11199) );
  INVX2 U11357 ( .A(\U_0/U_0/U_0/temp[1] ), .Y(n11200) );
  INVX2 U11358 ( .A(\U_0/U_0/U_0/temp[2] ), .Y(n11201) );
  INVX2 U11359 ( .A(\U_0/U_0/U_0/temp[3] ), .Y(n11202) );
  INVX2 U11360 ( .A(\U_0/U_0/U_0/temp[4] ), .Y(n11203) );
  INVX2 U11361 ( .A(\U_0/U_0/U_0/temp[5] ), .Y(n11204) );
  INVX2 U11362 ( .A(\U_0/U_0/U_0/temp[7] ), .Y(n11205) );
  INVX2 U11363 ( .A(\U_0/U_0/U_0/currentProcessedData [7]), .Y(n11206) );
  INVX2 U11364 ( .A(\U_0/PROCESSED_DATA [7]), .Y(n11207) );
  INVX2 U11365 ( .A(\U_0/U_0/U_0/currentProcessedData [6]), .Y(n11208) );
  INVX2 U11366 ( .A(n3361), .Y(n11209) );
  INVX2 U11367 ( .A(\U_0/PROCESSED_DATA [6]), .Y(n11210) );
  INVX2 U11368 ( .A(\U_0/U_0/U_0/currentProcessedData [5]), .Y(n11211) );
  INVX2 U11369 ( .A(\U_0/U_0/U_0/currentProcessedData [4]), .Y(n11212) );
  INVX2 U11370 ( .A(\U_0/PROCESSED_DATA [4]), .Y(n11213) );
  INVX2 U11371 ( .A(\U_0/U_0/U_0/currentProcessedData [3]), .Y(n11214) );
  INVX2 U11372 ( .A(\U_0/U_0/U_0/currentProcessedData [2]), .Y(n11215) );
  INVX2 U11373 ( .A(\U_0/U_0/U_0/currentProcessedData [1]), .Y(n11216) );
  INVX2 U11374 ( .A(\U_0/U_0/U_0/currentProcessedData [0]), .Y(n11217) );
  INVX2 U11375 ( .A(\U_0/U_3/TX_CRC [15]), .Y(n11218) );
  INVX2 U11376 ( .A(\U_0/U_3/TX_CRC [1]), .Y(n11219) );
  INVX2 U11377 ( .A(\U_0/U_3/TX_CRC [9]), .Y(n11220) );
  INVX2 U11378 ( .A(\U_0/U_3/TX_CRC [2]), .Y(n11221) );
  INVX2 U11379 ( .A(\U_0/U_3/TX_CRC [10]), .Y(n11222) );
  INVX2 U11380 ( .A(\U_0/U_3/TX_CRC [3]), .Y(n11223) );
  INVX2 U11381 ( .A(\U_0/U_3/TX_CRC [11]), .Y(n11224) );
  INVX2 U11382 ( .A(\U_0/U_3/TX_CRC [4]), .Y(n11225) );
  INVX2 U11383 ( .A(\U_0/U_3/TX_CRC [12]), .Y(n11226) );
  INVX2 U11384 ( .A(\U_0/U_3/TX_CRC [5]), .Y(n11227) );
  INVX2 U11385 ( .A(\U_0/U_3/TX_CRC [13]), .Y(n11228) );
  INVX2 U11386 ( .A(\U_0/U_3/TX_CRC [6]), .Y(n11229) );
  INVX2 U11387 ( .A(\U_0/U_3/TX_CRC [14]), .Y(n11230) );
  INVX2 U11388 ( .A(\U_0/U_3/TX_CRC [7]), .Y(n11231) );
  INVX2 U11389 ( .A(\U_0/U_3/TX_CRC [0]), .Y(n11232) );
  INVX2 U11390 ( .A(\U_0/U_3/TX_CRC [8]), .Y(n11233) );
  INVX2 U11391 ( .A(\U_0/U_0/U_0/fdata [6]), .Y(n11234) );
  INVX2 U11392 ( .A(\U_0/U_0/U_0/fdata [5]), .Y(n11235) );
  INVX2 U11393 ( .A(\U_0/U_0/U_0/fdata [4]), .Y(n11236) );
  INVX2 U11394 ( .A(\U_0/U_0/U_0/fdata [3]), .Y(n11237) );
  INVX2 U11395 ( .A(\U_0/U_0/U_0/fdata [2]), .Y(n11238) );
  INVX2 U11396 ( .A(\U_0/U_0/U_0/fdata [1]), .Y(n11239) );
  INVX2 U11397 ( .A(\U_0/U_0/U_0/fdata [0]), .Y(n11240) );
  INVX2 U11398 ( .A(\U_0/U_0/U_0/si[7] ), .Y(n11241) );
  INVX2 U11399 ( .A(\U_0/U_0/U_0/si[0] ), .Y(n11242) );
  INVX2 U11400 ( .A(n6920), .Y(n11243) );
  INVX2 U11401 ( .A(n6921), .Y(n11244) );
  INVX2 U11402 ( .A(\U_0/U_0/U_0/keyi[1] ), .Y(n11245) );
  INVX2 U11403 ( .A(n6922), .Y(n11246) );
  INVX2 U11404 ( .A(n6923), .Y(n11247) );
  INVX2 U11405 ( .A(\U_0/U_0/U_0/si[2] ), .Y(n11248) );
  INVX2 U11406 ( .A(\U_0/U_0/U_0/keyi[2] ), .Y(n11249) );
  INVX2 U11407 ( .A(\U_0/U_0/U_0/si[4] ), .Y(n11250) );
  INVX2 U11408 ( .A(\U_0/U_0/U_0/si[5] ), .Y(n11251) );
  INVX2 U11409 ( .A(\U_0/U_0/U_0/si[6] ), .Y(n11252) );
  INVX2 U11410 ( .A(\U_0/U_0/U_0/keyi[0] ), .Y(n11253) );
  INVX2 U11411 ( .A(\U_0/U_0/U_0/fdata [7]), .Y(n11254) );
  INVX2 U11412 ( .A(\U_0/U_0/U_0/keyTable[0][6] ), .Y(n11255) );
  INVX2 U11413 ( .A(\U_0/U_0/U_0/keyTable[0][5] ), .Y(n11256) );
  INVX2 U11414 ( .A(\U_0/U_0/U_0/keyTable[0][4] ), .Y(n11257) );
  INVX2 U11415 ( .A(\U_0/U_0/U_0/keyTable[0][3] ), .Y(n11258) );
  INVX2 U11416 ( .A(\U_0/U_0/U_0/keyTable[0][2] ), .Y(n11259) );
  INVX2 U11417 ( .A(\U_0/U_0/U_0/keyTable[0][1] ), .Y(n11260) );
  INVX2 U11418 ( .A(\U_0/U_0/U_0/keyTable[0][0] ), .Y(n11261) );
  INVX2 U11419 ( .A(\U_0/U_0/U_0/keyTable[1][7] ), .Y(n11262) );
  INVX2 U11420 ( .A(\U_0/U_0/U_0/keyTable[0][7] ), .Y(n11263) );
  INVX2 U11421 ( .A(\U_0/U_0/U_0/keyTable[3][0] ), .Y(n11264) );
  INVX2 U11422 ( .A(\U_0/U_0/U_0/keyTable[3][1] ), .Y(n11265) );
  INVX2 U11423 ( .A(\U_0/U_0/U_0/keyTable[3][2] ), .Y(n11266) );
  INVX2 U11424 ( .A(\U_0/U_0/U_0/keyTable[3][3] ), .Y(n11267) );
  INVX2 U11425 ( .A(\U_0/U_0/U_0/keyTable[3][4] ), .Y(n11268) );
  INVX2 U11426 ( .A(\U_0/U_0/U_0/keyTable[3][5] ), .Y(n11269) );
  INVX2 U11427 ( .A(\U_0/U_0/U_0/keyTable[3][6] ), .Y(n11270) );
  INVX2 U11428 ( .A(\U_0/U_0/U_0/keyTable[3][7] ), .Y(n11271) );
  INVX2 U11429 ( .A(\U_0/U_0/U_0/keyTable[2][0] ), .Y(n11272) );
  INVX2 U11430 ( .A(\U_0/U_0/U_0/keyTable[2][1] ), .Y(n11273) );
  INVX2 U11431 ( .A(\U_0/U_0/U_0/keyTable[2][2] ), .Y(n11274) );
  INVX2 U11432 ( .A(\U_0/U_0/U_0/keyTable[2][3] ), .Y(n11275) );
  INVX2 U11433 ( .A(\U_0/U_0/U_0/keyTable[2][4] ), .Y(n11276) );
  INVX2 U11434 ( .A(\U_0/U_0/U_0/keyTable[2][5] ), .Y(n11277) );
  INVX2 U11435 ( .A(\U_0/U_0/U_0/keyTable[2][6] ), .Y(n11278) );
  INVX2 U11436 ( .A(\U_0/U_0/U_0/keyTable[2][7] ), .Y(n11279) );
  INVX2 U11437 ( .A(\U_0/U_0/U_0/keyTable[1][0] ), .Y(n11280) );
  INVX2 U11438 ( .A(\U_0/U_0/U_0/keyTable[1][1] ), .Y(n11281) );
  INVX2 U11439 ( .A(\U_0/U_0/U_0/keyTable[1][2] ), .Y(n11282) );
  INVX2 U11440 ( .A(\U_0/U_0/U_0/keyTable[1][3] ), .Y(n11283) );
  INVX2 U11441 ( .A(\U_0/U_0/U_0/keyTable[1][4] ), .Y(n11284) );
  INVX2 U11442 ( .A(\U_0/U_0/U_0/keyTable[1][5] ), .Y(n11285) );
  INVX2 U11443 ( .A(\U_0/U_0/U_0/keyTable[1][6] ), .Y(n11286) );
  INVX2 U11444 ( .A(\U_0/U_1/U_0/tempOpcode [1]), .Y(n11287) );
  INVX2 U11445 ( .A(\U_0/U_3/U_3/flop_data [7]), .Y(n11288) );
  INVX2 U11446 ( .A(\U_0/U_3/U_3/current_send_data [6]), .Y(n11289) );
  INVX2 U11447 ( .A(\U_0/U_3/send_data [6]), .Y(n11290) );
  INVX2 U11448 ( .A(\U_0/U_3/U_3/current_send_data [5]), .Y(n11291) );
  INVX2 U11449 ( .A(\U_0/U_3/send_data [5]), .Y(n11292) );
  INVX2 U11450 ( .A(\U_0/U_3/U_3/current_send_data [4]), .Y(n11293) );
  INVX2 U11451 ( .A(\U_0/U_3/send_data [4]), .Y(n11294) );
  INVX2 U11452 ( .A(\U_0/U_3/U_3/current_send_data [3]), .Y(n11295) );
  INVX2 U11453 ( .A(\U_0/U_3/send_data [3]), .Y(n11296) );
  INVX2 U11454 ( .A(\U_0/U_3/U_3/current_send_data [2]), .Y(n11297) );
  INVX2 U11455 ( .A(\U_0/U_3/send_data [2]), .Y(n11298) );
  INVX2 U11456 ( .A(\U_0/U_3/U_3/current_send_data [1]), .Y(n11299) );
  INVX2 U11457 ( .A(\U_0/U_3/send_data [1]), .Y(n11300) );
  INVX2 U11458 ( .A(\U_0/U_3/U_3/current_send_data [0]), .Y(n11301) );
  INVX2 U11459 ( .A(\U_0/U_3/send_data [0]), .Y(n11302) );
  INVX2 U11460 ( .A(\U_0/U_3/U_3/current_send_data [7]), .Y(n11303) );
  INVX2 U11461 ( .A(\U_0/U_3/U_4/count[0] ), .Y(n11304) );
  INVX2 U11462 ( .A(\U_0/U_3/U_4/count[2] ), .Y(n11305) );
  INVX2 U11463 ( .A(\U_0/U_3/U_4/count[1] ), .Y(n11306) );
  INVX2 U11464 ( .A(\U_0/U_3/U_2/count[1] ), .Y(n11307) );
  INVX2 U11465 ( .A(\U_0/U_3/U_2/count[2] ), .Y(n11308) );
  INVX2 U11466 ( .A(\U_0/U_3/U_2/count[0] ), .Y(n11309) );
  INVX2 U11467 ( .A(\U_0/U_3/d_encode ), .Y(n11310) );
  INVX2 U11468 ( .A(\U_0/U_3/U_0/DE_holdout_BS ), .Y(n11311) );
  INVX2 U11469 ( .A(\U_1/U_0/U_1/U_2/nextState[0] ), .Y(n11312) );
  INVX2 U11470 ( .A(\U_1/U_0/U_1/U_7/nextState[7] ), .Y(n11313) );
  INVX2 U11471 ( .A(\U_1/U_0/U_1/U_7/nextState[6] ), .Y(n11314) );
  INVX2 U11472 ( .A(n3266), .Y(n11315) );
  INVX2 U11473 ( .A(\U_1/U_0/U_1/U_7/nextState[5] ), .Y(n11316) );
  INVX2 U11474 ( .A(\U_1/U_0/U_1/U_7/state[5] ), .Y(n11317) );
  INVX2 U11475 ( .A(\U_1/U_0/U_1/STOP_DATA [1]), .Y(n11318) );
  INVX2 U11476 ( .A(\U_1/U_0/U_1/STOP_DATA [0]), .Y(n11319) );
  INVX2 U11477 ( .A(\U_1/U_0/U_1/U_2/nextState[2] ), .Y(n11320) );
  INVX2 U11478 ( .A(n6055), .Y(n11321) );
  INVX2 U11479 ( .A(\U_1/U_0/U_1/U_2/nextState[1] ), .Y(n11322) );
  INVX2 U11480 ( .A(\U_1/U_0/U_1/U_2/timerRunning ), .Y(n11323) );
  INVX2 U11481 ( .A(\U_1/U_0/U_1/U_2/N99 ), .Y(n11324) );
  INVX2 U11482 ( .A(\U_1/U_0/U_1/U_2/state[1] ), .Y(n11325) );
  INVX2 U11483 ( .A(\U_1/U_0/U_1/U_2/state[2] ), .Y(n11326) );
  INVX2 U11484 ( .A(n460), .Y(n11327) );
  INVX2 U11485 ( .A(\U_1/U_0/U_1/CHK_ERROR ), .Y(n11328) );
  INVX2 U11486 ( .A(\U_1/U_0/U_1/SBC_CLR ), .Y(n11329) );
  INVX2 U11487 ( .A(\U_1/U_0/U_1/TIMER_TRIG ), .Y(n11330) );
  INVX2 U11488 ( .A(\U_1/U_0/U_1/U_7/nextState[0] ), .Y(n11331) );
  INVX2 U11489 ( .A(\U_1/U_0/U_1/U_7/nextState[1] ), .Y(n11332) );
  INVX2 U11490 ( .A(\U_1/U_0/U_1/U_7/state[1] ), .Y(n11333) );
  INVX2 U11491 ( .A(\U_1/U_0/U_1/U_7/nextState[2] ), .Y(n11334) );
  INVX2 U11492 ( .A(\U_1/U_0/U_1/U_7/state[2] ), .Y(n11335) );
  INVX2 U11493 ( .A(\U_1/U_0/U_1/U_7/nextState[3] ), .Y(n11336) );
  INVX2 U11494 ( .A(\U_1/U_0/U_1/U_7/nextState[4] ), .Y(n11337) );
  INVX2 U11495 ( .A(\U_1/U_0/U_1/U_7/state[4] ), .Y(n11338) );
  INVX2 U11496 ( .A(\U_1/U_0/U_1/SBC_EN ), .Y(n11339) );
  INVX2 U11497 ( .A(n3203), .Y(n11340) );
  INVX2 U11498 ( .A(\U_1/U_0/U_1/SBE ), .Y(n11341) );
  INVX2 U11499 ( .A(n3132), .Y(n11342) );
  INVX2 U11500 ( .A(n6219), .Y(n11343) );
  INVX2 U11501 ( .A(n6218), .Y(n11344) );
  INVX2 U11502 ( .A(n6232), .Y(n11345) );
  INVX2 U11503 ( .A(n3162), .Y(n11346) );
  INVX2 U11504 ( .A(n3227), .Y(n11347) );
  INVX2 U11505 ( .A(n3200), .Y(n11348) );
  INVX2 U11506 ( .A(\U_1/U_0/U_1/U_8/state[0] ), .Y(n11349) );
  INVX2 U11507 ( .A(n3183), .Y(n11350) );
  INVX2 U11508 ( .A(n3231), .Y(n11351) );
  INVX2 U11509 ( .A(n3223), .Y(n11352) );
  INVX2 U11510 ( .A(n3184), .Y(n11353) );
  INVX2 U11511 ( .A(n3222), .Y(n11354) );
  INVX2 U11512 ( .A(\U_1/U_0/U_1/U_8/keyCount[1] ), .Y(n11355) );
  INVX2 U11513 ( .A(\U_1/U_0/U_1/U_8/keyCount[2] ), .Y(n11356) );
  INVX2 U11514 ( .A(\U_1/U_0/U_1/U_8/state[2] ), .Y(n11357) );
  INVX2 U11515 ( .A(\U_1/U_0/U_1/U_8/keyCount[0] ), .Y(n11358) );
  INVX2 U11516 ( .A(\U_1/U_0/U_1/U_8/state[3] ), .Y(n11359) );
  INVX2 U11517 ( .A(\U_1/U_0/U_1/U_8/state[1] ), .Y(n11360) );
  INVX2 U11518 ( .A(\U_1/RBUF_FULL ), .Y(n11361) );
  INVX2 U11519 ( .A(\U_1/U_0/U_1/OE ), .Y(n11362) );
  INVX2 U11520 ( .A(n2327), .Y(n11363) );
  INVX2 U11521 ( .A(n2411), .Y(n11364) );
  INVX2 U11522 ( .A(n2530), .Y(n11365) );
  INVX2 U11523 ( .A(n2566), .Y(n11366) );
  INVX2 U11524 ( .A(n2645), .Y(n11367) );
  INVX2 U11525 ( .A(n2760), .Y(n11368) );
  INVX2 U11526 ( .A(n2796), .Y(n11369) );
  INVX2 U11527 ( .A(n2875), .Y(n11370) );
  INVX2 U11528 ( .A(n2990), .Y(n11371) );
  INVX2 U11529 ( .A(n3026), .Y(n11372) );
  INVX2 U11530 ( .A(n3109), .Y(n11373) );
  INVX2 U11531 ( .A(n3112), .Y(n11375) );
  INVX2 U11532 ( .A(n2911), .Y(n11376) );
  INVX2 U11533 ( .A(n2681), .Y(n11377) );
  INVX2 U11534 ( .A(n2451), .Y(n11378) );
  INVX2 U11535 ( .A(n2176), .Y(n11379) );
  INVX2 U11536 ( .A(n2216), .Y(n11380) );
  INVX2 U11537 ( .A(n2284), .Y(n11381) );
  INVX2 U11538 ( .A(n2358), .Y(n11382) );
  INVX2 U11539 ( .A(n2443), .Y(n11383) );
  INVX2 U11540 ( .A(n2558), .Y(n11384) );
  INVX2 U11541 ( .A(n2595), .Y(n11385) );
  INVX2 U11542 ( .A(n2673), .Y(n11386) );
  INVX2 U11543 ( .A(n2788), .Y(n11387) );
  INVX2 U11544 ( .A(n2825), .Y(n11388) );
  INVX2 U11545 ( .A(n2903), .Y(n11389) );
  INVX2 U11546 ( .A(n3018), .Y(n11390) );
  INVX2 U11547 ( .A(n3056), .Y(n11391) );
  INVX2 U11548 ( .A(n3140), .Y(n11392) );
  INVX2 U11549 ( .A(n2940), .Y(n11394) );
  INVX2 U11550 ( .A(n2710), .Y(n11395) );
  INVX2 U11551 ( .A(n2480), .Y(n11396) );
  INVX2 U11552 ( .A(n2169), .Y(n11397) );
  INVX2 U11553 ( .A(n2299), .Y(n11398) );
  INVX2 U11554 ( .A(n2256), .Y(n11399) );
  INVX2 U11555 ( .A(n2351), .Y(n11400) );
  INVX2 U11556 ( .A(n2474), .Y(n11401) );
  INVX2 U11557 ( .A(n2508), .Y(n11402) );
  INVX2 U11558 ( .A(n2589), .Y(n11403) );
  INVX2 U11559 ( .A(n2704), .Y(n11404) );
  INVX2 U11560 ( .A(n2738), .Y(n11405) );
  INVX2 U11561 ( .A(n2819), .Y(n11406) );
  INVX2 U11562 ( .A(n2934), .Y(n11407) );
  INVX2 U11563 ( .A(n2968), .Y(n11408) );
  INVX2 U11564 ( .A(n3049), .Y(n11409) );
  INVX2 U11565 ( .A(n3095), .Y(n11411) );
  INVX2 U11566 ( .A(n2853), .Y(n11412) );
  INVX2 U11567 ( .A(n2623), .Y(n11413) );
  INVX2 U11568 ( .A(n2388), .Y(n11414) );
  INVX2 U11569 ( .A(n2191), .Y(n11415) );
  INVX2 U11570 ( .A(n2293), .Y(n11416) );
  INVX2 U11571 ( .A(n2381), .Y(n11417) );
  INVX2 U11572 ( .A(n2502), .Y(n11418) );
  INVX2 U11573 ( .A(n2536), .Y(n11419) );
  INVX2 U11574 ( .A(n2617), .Y(n11420) );
  INVX2 U11575 ( .A(n2732), .Y(n11421) );
  INVX2 U11576 ( .A(n2766), .Y(n11422) );
  INVX2 U11577 ( .A(n2847), .Y(n11423) );
  INVX2 U11578 ( .A(n2962), .Y(n11424) );
  INVX2 U11579 ( .A(n2996), .Y(n11425) );
  INVX2 U11580 ( .A(n3078), .Y(n11426) );
  INVX2 U11581 ( .A(n3081), .Y(n11428) );
  INVX2 U11582 ( .A(n2881), .Y(n11429) );
  INVX2 U11583 ( .A(n2651), .Y(n11430) );
  INVX2 U11584 ( .A(n2418), .Y(n11431) );
  INVX2 U11585 ( .A(n2183), .Y(n11432) );
  INVX2 U11586 ( .A(\U_1/U_0/U_1/U_8/address[0] ), .Y(n11433) );
  INVX2 U11587 ( .A(n2343), .Y(n11434) );
  INVX2 U11588 ( .A(n2426), .Y(n11435) );
  INVX2 U11589 ( .A(n2544), .Y(n11436) );
  INVX2 U11590 ( .A(n2581), .Y(n11437) );
  INVX2 U11591 ( .A(n2659), .Y(n11438) );
  INVX2 U11592 ( .A(n2774), .Y(n11439) );
  INVX2 U11593 ( .A(n2811), .Y(n11440) );
  INVX2 U11594 ( .A(n2889), .Y(n11441) );
  INVX2 U11595 ( .A(n3004), .Y(n11442) );
  INVX2 U11596 ( .A(n3041), .Y(n11443) );
  INVX2 U11597 ( .A(n3122), .Y(n11444) );
  INVX2 U11598 ( .A(n3125), .Y(n11446) );
  INVX2 U11599 ( .A(n2926), .Y(n11447) );
  INVX2 U11600 ( .A(n2696), .Y(n11448) );
  INVX2 U11601 ( .A(n2466), .Y(n11449) );
  INVX2 U11602 ( .A(n2217), .Y(n11450) );
  INVX2 U11603 ( .A(n2335), .Y(n11451) );
  INVX2 U11604 ( .A(n2459), .Y(n11452) );
  INVX2 U11605 ( .A(n2494), .Y(n11453) );
  INVX2 U11606 ( .A(n2574), .Y(n11454) );
  INVX2 U11607 ( .A(n2689), .Y(n11455) );
  INVX2 U11608 ( .A(n2724), .Y(n11456) );
  INVX2 U11609 ( .A(n2804), .Y(n11457) );
  INVX2 U11610 ( .A(n2919), .Y(n11458) );
  INVX2 U11611 ( .A(n2954), .Y(n11459) );
  INVX2 U11612 ( .A(n3034), .Y(n11460) );
  INVX2 U11613 ( .A(n3070), .Y(n11462) );
  INVX2 U11614 ( .A(n2839), .Y(n11463) );
  INVX2 U11615 ( .A(n2609), .Y(n11464) );
  INVX2 U11616 ( .A(n2373), .Y(n11465) );
  INVX2 U11617 ( .A(n2194), .Y(n11466) );
  INVX2 U11618 ( .A(n2366), .Y(n11468) );
  INVX2 U11619 ( .A(n2488), .Y(n11469) );
  INVX2 U11620 ( .A(n2522), .Y(n11470) );
  INVX2 U11621 ( .A(n2603), .Y(n11471) );
  INVX2 U11622 ( .A(n2718), .Y(n11472) );
  INVX2 U11623 ( .A(n2752), .Y(n11473) );
  INVX2 U11624 ( .A(n2833), .Y(n11474) );
  INVX2 U11625 ( .A(n2948), .Y(n11475) );
  INVX2 U11626 ( .A(n2982), .Y(n11476) );
  INVX2 U11627 ( .A(n3064), .Y(n11477) );
  INVX2 U11628 ( .A(n3083), .Y(n11479) );
  INVX2 U11629 ( .A(n2867), .Y(n11480) );
  INVX2 U11630 ( .A(n2637), .Y(n11481) );
  INVX2 U11631 ( .A(n2403), .Y(n11482) );
  INVX2 U11632 ( .A(n2187), .Y(n11483) );
  INVX2 U11633 ( .A(n2230), .Y(n11484) );
  INVX2 U11634 ( .A(n2309), .Y(n11485) );
  INVX2 U11635 ( .A(n2396), .Y(n11486) );
  INVX2 U11636 ( .A(n2516), .Y(n11487) );
  INVX2 U11637 ( .A(n2550), .Y(n11488) );
  INVX2 U11638 ( .A(n2631), .Y(n11489) );
  INVX2 U11639 ( .A(n2746), .Y(n11490) );
  INVX2 U11640 ( .A(n2780), .Y(n11491) );
  INVX2 U11641 ( .A(n2861), .Y(n11492) );
  INVX2 U11642 ( .A(n2976), .Y(n11493) );
  INVX2 U11643 ( .A(n3010), .Y(n11494) );
  INVX2 U11644 ( .A(n3094), .Y(n11495) );
  INVX2 U11645 ( .A(n3098), .Y(n11497) );
  INVX2 U11646 ( .A(n2895), .Y(n11498) );
  INVX2 U11647 ( .A(n2665), .Y(n11499) );
  INVX2 U11648 ( .A(n2435), .Y(n11500) );
  INVX2 U11649 ( .A(n2181), .Y(n11501) );
  INVX2 U11650 ( .A(n2264), .Y(n11502) );
  INVX2 U11651 ( .A(\U_1/U_0/U_1/U_8/address[1] ), .Y(n11503) );
  INVX2 U11652 ( .A(\U_1/U_0/U_1/U_8/address[2] ), .Y(n11504) );
  INVX2 U11653 ( .A(\U_1/U_0/U_1/U_8/address[6] ), .Y(n11505) );
  INVX2 U11654 ( .A(n3141), .Y(n11506) );
  INVX2 U11655 ( .A(\U_1/U_0/U_1/U_8/address[7] ), .Y(n11507) );
  INVX2 U11656 ( .A(n2196), .Y(n11509) );
  INVX2 U11657 ( .A(\U_1/U_0/U_1/U_8/address[5] ), .Y(n11510) );
  INVX2 U11658 ( .A(\U_1/U_0/U_1/U_8/address[4] ), .Y(n11511) );
  INVX2 U11659 ( .A(\U_1/U_0/U_1/LOAD_DATA [7]), .Y(n11512) );
  INVX2 U11660 ( .A(\U_1/U_0/U_1/RCV_DATA [7]), .Y(n11513) );
  INVX2 U11661 ( .A(\U_1/U_0/U_1/LOAD_DATA [6]), .Y(n11514) );
  INVX2 U11662 ( .A(\U_1/U_0/U_1/LOAD_DATA [5]), .Y(n11515) );
  INVX2 U11663 ( .A(\U_1/U_0/U_1/RCV_DATA [5]), .Y(n11516) );
  INVX2 U11664 ( .A(\U_1/U_0/U_1/LOAD_DATA [4]), .Y(n11517) );
  INVX2 U11665 ( .A(\U_1/U_0/U_1/RCV_DATA [4]), .Y(n11518) );
  INVX2 U11666 ( .A(\U_1/U_0/U_1/LOAD_DATA [3]), .Y(n11519) );
  INVX2 U11667 ( .A(\U_1/U_0/U_1/RCV_DATA [3]), .Y(n11520) );
  INVX2 U11668 ( .A(\U_1/U_0/U_1/LOAD_DATA [2]), .Y(n11521) );
  INVX2 U11669 ( .A(\U_1/U_0/U_1/LOAD_DATA [1]), .Y(n11522) );
  INVX2 U11670 ( .A(\U_1/U_0/U_1/RCV_DATA [1]), .Y(n11523) );
  INVX2 U11671 ( .A(\U_1/U_0/U_1/LOAD_DATA [0]), .Y(n11524) );
  INVX2 U11672 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[0] ), .Y(n11525) );
  INVX2 U11673 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[1] ), .Y(n11526) );
  INVX2 U11674 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[2] ), .Y(n11527) );
  INVX2 U11675 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[3] ), .Y(n11528) );
  INVX2 U11676 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[4] ), .Y(n11529) );
  INVX2 U11677 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[5] ), .Y(n11530) );
  INVX2 U11678 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[6] ), .Y(n11531) );
  INVX2 U11679 ( .A(\U_1/U_0/U_1/U_8/parityAccumulator[7] ), .Y(n11532) );
  INVX2 U11680 ( .A(\U_1/U_0/U_1/U_8/parityError ), .Y(n11533) );
  INVX2 U11681 ( .A(\U_1/U_0/U_1/U_8/currentPlainKey[0] ), .Y(n11534) );
  INVX2 U11682 ( .A(\U_1/U_0/PLAINKEY [0]), .Y(n11535) );
  INVX2 U11683 ( .A(\U_1/U_0/U_1/U_8/currentPlainKey[1] ), .Y(n11536) );
  INVX2 U11684 ( .A(\U_1/U_0/PLAINKEY [1]), .Y(n11537) );
  INVX2 U11685 ( .A(\U_1/U_0/U_1/U_8/currentPlainKey[2] ), .Y(n11538) );
  INVX2 U11686 ( .A(\U_1/U_0/PLAINKEY [2]), .Y(n11539) );
  INVX2 U11687 ( .A(\U_1/U_0/U_1/U_8/currentPlainKey[3] ), .Y(n11540) );
  INVX2 U11688 ( .A(\U_1/U_0/PLAINKEY [3]), .Y(n11541) );
  INVX2 U11689 ( .A(\U_1/U_0/U_1/U_8/currentPlainKey[63] ), .Y(n11542) );
  INVX2 U11690 ( .A(\U_1/U_0/PLAINKEY [63]), .Y(n11543) );
  INVX2 U11691 ( .A(n5932), .Y(n11544) );
  INVX2 U11692 ( .A(n1914), .Y(n11545) );
  INVX2 U11693 ( .A(n5913), .Y(n11546) );
  INVX2 U11694 ( .A(n6008), .Y(n11547) );
  INVX2 U11695 ( .A(n2128), .Y(n11548) );
  INVX2 U11696 ( .A(n5948), .Y(n11549) );
  INVX2 U11697 ( .A(n6007), .Y(n11550) );
  INVX2 U11698 ( .A(n5947), .Y(n11551) );
  INVX2 U11699 ( .A(\U_1/U_2/U_5/state[0] ), .Y(n11552) );
  INVX2 U11700 ( .A(n6006), .Y(n11553) );
  INVX2 U11701 ( .A(n5951), .Y(n11554) );
  INVX2 U11702 ( .A(n2115), .Y(n11555) );
  INVX2 U11703 ( .A(n2110), .Y(n11556) );
  INVX2 U11704 ( .A(\U_1/U_2/U_5/state[3] ), .Y(n11558) );
  INVX2 U11705 ( .A(n5907), .Y(n11559) );
  INVX2 U11706 ( .A(\U_1/U_2/U_7/count[2] ), .Y(n11560) );
  INVX2 U11707 ( .A(n5929), .Y(BSE_S) );
  INVX2 U11708 ( .A(n774), .Y(n11562) );
  INVX2 U11709 ( .A(n2162), .Y(n11563) );
  INVX2 U11710 ( .A(\U_1/U_2/U_1/state[0] ), .Y(n11564) );
  INVX2 U11711 ( .A(n2155), .Y(n11565) );
  INVX2 U11712 ( .A(\U_1/U_2/U_1/DP_hold2 ), .Y(n11566) );
  INVX2 U11713 ( .A(\U_1/U_2/U_1/state[3] ), .Y(n11567) );
  INVX2 U11714 ( .A(\U_1/U_2/U_1/state[1] ), .Y(n11568) );
  INVX2 U11715 ( .A(n5953), .Y(n11569) );
  INVX2 U11716 ( .A(\U_1/U_2/U_5/N170 ), .Y(n11570) );
  INVX2 U11717 ( .A(\U_1/U_2/rx_CHECK_CRC [7]), .Y(n11571) );
  INVX2 U11718 ( .A(n2142), .Y(n11572) );
  INVX2 U11719 ( .A(\U_1/U_2/U_5/count[0] ), .Y(n11573) );
  INVX2 U11720 ( .A(\U_1/U_2/U_5/count[1] ), .Y(n11574) );
  INVX2 U11721 ( .A(\U_1/U_2/U_5/count[2] ), .Y(n11575) );
  INVX2 U11722 ( .A(\U_1/U_2/U_5/count[3] ), .Y(n11576) );
  INVX2 U11723 ( .A(\U_1/U_2/U_2/current_crc[15] ), .Y(n11578) );
  INVX2 U11724 ( .A(\U_1/U_2/U_2/current_crc[0] ), .Y(n11579) );
  INVX2 U11725 ( .A(\U_1/U_2/U_2/cache_1 [0]), .Y(n11580) );
  INVX2 U11726 ( .A(\U_1/U_2/U_2/current_crc[8] ), .Y(n11581) );
  INVX2 U11727 ( .A(\U_1/U_2/U_2/current_crc[2] ), .Y(n11582) );
  INVX2 U11728 ( .A(\U_1/U_2/U_2/cache_1 [2]), .Y(n11583) );
  INVX2 U11729 ( .A(\U_1/U_2/U_2/current_crc[10] ), .Y(n11584) );
  INVX2 U11730 ( .A(\U_1/U_2/U_2/current_crc[3] ), .Y(n11585) );
  INVX2 U11731 ( .A(\U_1/U_2/U_2/cache_1 [3]), .Y(n11586) );
  INVX2 U11732 ( .A(\U_1/U_2/U_2/current_crc[11] ), .Y(n11587) );
  INVX2 U11733 ( .A(\U_1/U_2/U_2/current_crc[4] ), .Y(n11588) );
  INVX2 U11734 ( .A(\U_1/U_2/U_2/cache_1 [4]), .Y(n11589) );
  INVX2 U11735 ( .A(\U_1/U_2/U_2/current_crc[12] ), .Y(n11590) );
  INVX2 U11736 ( .A(\U_1/U_2/U_2/cache_1 [12]), .Y(n11591) );
  INVX2 U11737 ( .A(\U_1/U_2/U_2/current_crc[5] ), .Y(n11592) );
  INVX2 U11738 ( .A(\U_1/U_2/U_2/cache_1 [5]), .Y(n11593) );
  INVX2 U11739 ( .A(\U_1/U_2/U_2/current_crc[13] ), .Y(n11594) );
  INVX2 U11740 ( .A(\U_1/U_2/U_2/current_crc[6] ), .Y(n11595) );
  INVX2 U11741 ( .A(\U_1/U_2/U_2/cache_1 [6]), .Y(n11596) );
  INVX2 U11742 ( .A(\U_1/U_2/U_2/current_crc[14] ), .Y(n11597) );
  INVX2 U11743 ( .A(\U_1/U_2/U_2/cache_1 [14]), .Y(n11598) );
  INVX2 U11744 ( .A(\U_1/U_2/U_2/current_crc[7] ), .Y(n11599) );
  INVX2 U11745 ( .A(\U_1/U_2/U_2/cache_1 [7]), .Y(n11600) );
  INVX2 U11746 ( .A(\U_1/U_2/U_2/cache_1 [13]), .Y(n11601) );
  INVX2 U11747 ( .A(\U_1/U_2/U_2/cache_1 [11]), .Y(n11602) );
  INVX2 U11748 ( .A(\U_1/U_2/U_2/current_crc[1] ), .Y(n11603) );
  INVX2 U11749 ( .A(\U_1/U_2/U_2/cache_1 [1]), .Y(n11604) );
  INVX2 U11750 ( .A(\U_1/U_2/U_2/current_crc[9] ), .Y(n11605) );
  INVX2 U11751 ( .A(\U_1/U_2/U_2/cache_1 [9]), .Y(n11606) );
  INVX2 U11752 ( .A(\U_1/U_2/U_2/cache_1 [10]), .Y(n11607) );
  INVX2 U11753 ( .A(\U_1/U_2/U_2/cache_1 [8]), .Y(n11608) );
  INVX2 U11754 ( .A(\U_1/U_2/U_2/cache_1 [15]), .Y(n11609) );
  INVX2 U11755 ( .A(\U_1/U_2/rx_CHECK_CRC [0]), .Y(n11610) );
  INVX2 U11756 ( .A(\U_1/U_2/rx_CHECK_CRC [2]), .Y(n11611) );
  INVX2 U11757 ( .A(\U_1/U_2/rx_CHECK_CRC [3]), .Y(n11612) );
  INVX2 U11758 ( .A(\U_1/U_2/rx_CHECK_CRC [4]), .Y(n11613) );
  INVX2 U11759 ( .A(\U_1/U_2/rx_CHECK_CRC [5]), .Y(n11614) );
  INVX2 U11760 ( .A(\U_1/U_2/rx_CHECK_CRC [6]), .Y(n11615) );
  INVX2 U11761 ( .A(\U_1/U_2/U_7/count[0] ), .Y(n11616) );
  INVX2 U11762 ( .A(\U_1/U_2/U_7/count[1] ), .Y(n11617) );
  INVX2 U11763 ( .A(\U_1/U_2/U_5/curR_ERROR ), .Y(n11618) );
  INVX2 U11764 ( .A(\U_1/U_2/U_5/curCRC_ERROR ), .Y(n11619) );
  INVX2 U11765 ( .A(n781), .Y(n11620) );
  INVX2 U11766 ( .A(n5877), .Y(n11621) );
  INVX2 U11767 ( .A(n5881), .Y(n11622) );
  INVX2 U11768 ( .A(\U_1/U_3/U_0/N59 ), .Y(n11623) );
  INVX2 U11769 ( .A(n9285), .Y(n11624) );
  INVX2 U11770 ( .A(n812), .Y(n11625) );
  INVX2 U11771 ( .A(n786), .Y(n11626) );
  INVX2 U11772 ( .A(\U_1/U_3/U_0/state[3] ), .Y(n11627) );
  INVX2 U11773 ( .A(n5849), .Y(n11628) );
  INVX2 U11774 ( .A(n5856), .Y(n11629) );
  INVX2 U11775 ( .A(n5860), .Y(n11630) );
  INVX2 U11776 ( .A(\U_1/U_3/U_0/DE_holdout ), .Y(n11631) );
  INVX2 U11777 ( .A(\U_1/U_3/U_0/DE_holdout_last ), .Y(n11632) );
  INVX2 U11778 ( .A(n785), .Y(n11633) );
  INVX2 U11779 ( .A(n5868), .Y(n11634) );
  INVX2 U11780 ( .A(n5854), .Y(n11635) );
  INVX2 U11781 ( .A(n5882), .Y(n11636) );
  INVX2 U11782 ( .A(\U_1/U_3/U_0/state[2] ), .Y(n11637) );
  INVX2 U11783 ( .A(\U_1/U_3/U_0/state[0] ), .Y(n11638) );
  INVX2 U11784 ( .A(\U_1/U_3/U_0/state[1] ), .Y(n11639) );
  INVX2 U11785 ( .A(slave_is_sending), .Y(n11640) );
  INVX2 U11786 ( .A(n790), .Y(n11641) );
  INVX2 U11787 ( .A(n5896), .Y(n11642) );
  INVX2 U11788 ( .A(n5816), .Y(n11643) );
  INVX2 U11789 ( .A(\U_1/U_3/U_3/N188 ), .Y(n11644) );
  INVX2 U11790 ( .A(n862), .Y(n11645) );
  INVX2 U11791 ( .A(n2004), .Y(n11646) );
  INVX2 U11792 ( .A(n5825), .Y(n11647) );
  INVX2 U11793 ( .A(n865), .Y(n11648) );
  INVX2 U11794 ( .A(n6018), .Y(n11649) );
  INVX2 U11795 ( .A(n6034), .Y(n11650) );
  INVX2 U11796 ( .A(\U_1/U_3/U_3/state[1] ), .Y(n11651) );
  INVX2 U11797 ( .A(n5815), .Y(n11652) );
  INVX2 U11798 ( .A(n877), .Y(n11653) );
  INVX2 U11799 ( .A(n5821), .Y(n11654) );
  INVX2 U11800 ( .A(\U_1/U_3/U_3/state[2] ), .Y(n11655) );
  INVX2 U11801 ( .A(\U_1/U_3/U_3/state[0] ), .Y(n11656) );
  INVX2 U11802 ( .A(\U_1/U_1/U_0/state[2] ), .Y(n11657) );
  INVX2 U11803 ( .A(n6027), .Y(n11658) );
  INVX2 U11804 ( .A(n6032), .Y(n11659) );
  INVX2 U11805 ( .A(\U_1/U_1/R_ENABLE ), .Y(n11660) );
  INVX2 U11806 ( .A(n1613), .Y(n11661) );
  INVX2 U11807 ( .A(n1628), .Y(n11662) );
  INVX2 U11808 ( .A(n1644), .Y(n11663) );
  INVX2 U11809 ( .A(n1657), .Y(n11664) );
  INVX2 U11810 ( .A(n1612), .Y(n11665) );
  INVX2 U11811 ( .A(n1626), .Y(n11666) );
  INVX2 U11812 ( .A(n1642), .Y(n11667) );
  INVX2 U11813 ( .A(n1658), .Y(n11668) );
  INVX2 U11814 ( .A(\U_1/U_1/U_1/writeptr[0] ), .Y(n11669) );
  INVX2 U11815 ( .A(\U_1/U_1/U_1/opcode[4][0] ), .Y(n11670) );
  INVX2 U11816 ( .A(\U_1/U_1/U_1/opcode[4][1] ), .Y(n11671) );
  INVX2 U11817 ( .A(\U_1/U_1/U_1/memory[4][0] ), .Y(n11672) );
  INVX2 U11818 ( .A(\U_1/U_1/U_1/memory[4][1] ), .Y(n11673) );
  INVX2 U11819 ( .A(\U_1/U_1/U_1/memory[4][2] ), .Y(n11674) );
  INVX2 U11820 ( .A(\U_1/U_1/U_1/memory[4][3] ), .Y(n11675) );
  INVX2 U11821 ( .A(\U_1/U_1/U_1/memory[4][4] ), .Y(n11676) );
  INVX2 U11822 ( .A(\U_1/U_1/U_1/memory[4][5] ), .Y(n11677) );
  INVX2 U11823 ( .A(\U_1/U_1/U_1/memory[4][6] ), .Y(n11678) );
  INVX2 U11824 ( .A(\U_1/U_1/U_1/memory[4][7] ), .Y(n11679) );
  INVX2 U11825 ( .A(\U_1/U_1/U_1/opcode[5][0] ), .Y(n11680) );
  INVX2 U11826 ( .A(\U_1/U_1/U_1/opcode[5][1] ), .Y(n11681) );
  INVX2 U11827 ( .A(\U_1/U_1/U_1/memory[5][0] ), .Y(n11682) );
  INVX2 U11828 ( .A(\U_1/U_1/U_1/memory[5][1] ), .Y(n11683) );
  INVX2 U11829 ( .A(\U_1/U_1/U_1/memory[5][2] ), .Y(n11684) );
  INVX2 U11830 ( .A(\U_1/U_1/U_1/memory[5][3] ), .Y(n11685) );
  INVX2 U11831 ( .A(\U_1/U_1/U_1/memory[5][4] ), .Y(n11686) );
  INVX2 U11832 ( .A(\U_1/U_1/U_1/memory[5][5] ), .Y(n11687) );
  INVX2 U11833 ( .A(\U_1/U_1/U_1/memory[5][6] ), .Y(n11688) );
  INVX2 U11834 ( .A(\U_1/U_1/U_1/memory[5][7] ), .Y(n11689) );
  INVX2 U11835 ( .A(\U_1/U_1/U_1/memory[6][0] ), .Y(n11690) );
  INVX2 U11836 ( .A(\U_1/U_1/U_1/memory[6][1] ), .Y(n11691) );
  INVX2 U11837 ( .A(\U_1/U_1/U_1/memory[6][2] ), .Y(n11692) );
  INVX2 U11838 ( .A(\U_1/U_1/U_1/memory[6][3] ), .Y(n11693) );
  INVX2 U11839 ( .A(\U_1/U_1/U_1/memory[6][4] ), .Y(n11694) );
  INVX2 U11840 ( .A(\U_1/U_1/U_1/memory[6][5] ), .Y(n11695) );
  INVX2 U11841 ( .A(\U_1/U_1/U_1/memory[6][6] ), .Y(n11696) );
  INVX2 U11842 ( .A(\U_1/U_1/U_1/memory[6][7] ), .Y(n11697) );
  INVX2 U11843 ( .A(\U_1/U_1/U_1/memory[7][6] ), .Y(n11698) );
  INVX2 U11844 ( .A(\U_1/U_1/U_1/memory[7][7] ), .Y(n11699) );
  INVX2 U11845 ( .A(\U_1/U_1/U_1/memory[7][0] ), .Y(n11700) );
  INVX2 U11846 ( .A(\U_1/U_1/U_1/memory[7][1] ), .Y(n11701) );
  INVX2 U11847 ( .A(\U_1/U_1/U_1/memory[7][2] ), .Y(n11702) );
  INVX2 U11848 ( .A(\U_1/U_1/U_1/memory[7][3] ), .Y(n11703) );
  INVX2 U11849 ( .A(\U_1/U_1/U_1/memory[7][4] ), .Y(n11704) );
  INVX2 U11850 ( .A(\U_1/U_1/U_1/memory[7][5] ), .Y(n11705) );
  INVX2 U11851 ( .A(\U_1/U_1/U_1/opcode[11][1] ), .Y(n11706) );
  INVX2 U11852 ( .A(\U_1/U_1/U_1/opcode[11][0] ), .Y(n11707) );
  INVX2 U11853 ( .A(\U_1/U_1/U_1/opcode[6][0] ), .Y(n11708) );
  INVX2 U11854 ( .A(\U_1/U_1/U_1/opcode[6][1] ), .Y(n11709) );
  INVX2 U11855 ( .A(\U_1/U_1/U_1/opcode[7][0] ), .Y(n11710) );
  INVX2 U11856 ( .A(\U_1/U_1/U_1/opcode[7][1] ), .Y(n11711) );
  INVX2 U11857 ( .A(\U_1/U_1/U_1/memory[11][0] ), .Y(n11712) );
  INVX2 U11858 ( .A(\U_1/U_1/U_1/memory[11][1] ), .Y(n11713) );
  INVX2 U11859 ( .A(\U_1/U_1/U_1/memory[11][2] ), .Y(n11714) );
  INVX2 U11860 ( .A(\U_1/U_1/U_1/memory[11][3] ), .Y(n11715) );
  INVX2 U11861 ( .A(\U_1/U_1/U_1/memory[11][4] ), .Y(n11716) );
  INVX2 U11862 ( .A(\U_1/U_1/U_1/memory[11][5] ), .Y(n11717) );
  INVX2 U11863 ( .A(\U_1/U_1/U_1/memory[11][6] ), .Y(n11718) );
  INVX2 U11864 ( .A(\U_1/U_1/U_1/memory[11][7] ), .Y(n11719) );
  INVX2 U11865 ( .A(\U_1/U_1/U_1/opcode[8][0] ), .Y(n11720) );
  INVX2 U11866 ( .A(\U_1/U_1/U_1/opcode[8][1] ), .Y(n11721) );
  INVX2 U11867 ( .A(\U_1/U_1/U_1/memory[8][0] ), .Y(n11722) );
  INVX2 U11868 ( .A(\U_1/U_1/U_1/memory[8][1] ), .Y(n11723) );
  INVX2 U11869 ( .A(\U_1/U_1/U_1/memory[8][2] ), .Y(n11724) );
  INVX2 U11870 ( .A(\U_1/U_1/U_1/memory[8][3] ), .Y(n11725) );
  INVX2 U11871 ( .A(\U_1/U_1/U_1/memory[8][4] ), .Y(n11726) );
  INVX2 U11872 ( .A(\U_1/U_1/U_1/memory[8][5] ), .Y(n11727) );
  INVX2 U11873 ( .A(\U_1/U_1/U_1/memory[8][6] ), .Y(n11728) );
  INVX2 U11874 ( .A(\U_1/U_1/U_1/memory[8][7] ), .Y(n11729) );
  INVX2 U11875 ( .A(\U_1/U_1/U_1/opcode[9][0] ), .Y(n11730) );
  INVX2 U11876 ( .A(\U_1/U_1/U_1/opcode[9][1] ), .Y(n11731) );
  INVX2 U11877 ( .A(\U_1/U_1/U_1/memory[9][0] ), .Y(n11732) );
  INVX2 U11878 ( .A(\U_1/U_1/U_1/memory[9][1] ), .Y(n11733) );
  INVX2 U11879 ( .A(\U_1/U_1/U_1/memory[9][2] ), .Y(n11734) );
  INVX2 U11880 ( .A(\U_1/U_1/U_1/memory[9][3] ), .Y(n11735) );
  INVX2 U11881 ( .A(\U_1/U_1/U_1/memory[9][4] ), .Y(n11736) );
  INVX2 U11882 ( .A(\U_1/U_1/U_1/memory[9][5] ), .Y(n11737) );
  INVX2 U11883 ( .A(\U_1/U_1/U_1/memory[9][6] ), .Y(n11738) );
  INVX2 U11884 ( .A(\U_1/U_1/U_1/memory[9][7] ), .Y(n11739) );
  INVX2 U11885 ( .A(\U_1/U_1/U_1/opcode[10][0] ), .Y(n11740) );
  INVX2 U11886 ( .A(\U_1/U_1/U_1/opcode[10][1] ), .Y(n11741) );
  INVX2 U11887 ( .A(\U_1/U_1/U_1/memory[10][0] ), .Y(n11742) );
  INVX2 U11888 ( .A(\U_1/U_1/U_1/memory[10][1] ), .Y(n11743) );
  INVX2 U11889 ( .A(\U_1/U_1/U_1/memory[10][2] ), .Y(n11744) );
  INVX2 U11890 ( .A(\U_1/U_1/U_1/memory[10][3] ), .Y(n11745) );
  INVX2 U11891 ( .A(\U_1/U_1/U_1/memory[10][4] ), .Y(n11746) );
  INVX2 U11892 ( .A(\U_1/U_1/U_1/memory[10][5] ), .Y(n11747) );
  INVX2 U11893 ( .A(\U_1/U_1/U_1/memory[10][6] ), .Y(n11748) );
  INVX2 U11894 ( .A(\U_1/U_1/U_1/memory[10][7] ), .Y(n11749) );
  INVX2 U11895 ( .A(\U_1/U_1/U_1/opcode[28][0] ), .Y(n11750) );
  INVX2 U11896 ( .A(\U_1/U_1/U_1/opcode[28][1] ), .Y(n11751) );
  INVX2 U11897 ( .A(\U_1/U_1/U_1/memory[28][0] ), .Y(n11752) );
  INVX2 U11898 ( .A(\U_1/U_1/U_1/memory[28][1] ), .Y(n11753) );
  INVX2 U11899 ( .A(\U_1/U_1/U_1/memory[28][2] ), .Y(n11754) );
  INVX2 U11900 ( .A(\U_1/U_1/U_1/memory[28][3] ), .Y(n11755) );
  INVX2 U11901 ( .A(\U_1/U_1/U_1/memory[28][4] ), .Y(n11756) );
  INVX2 U11902 ( .A(\U_1/U_1/U_1/memory[28][5] ), .Y(n11757) );
  INVX2 U11903 ( .A(\U_1/U_1/U_1/memory[28][6] ), .Y(n11758) );
  INVX2 U11904 ( .A(\U_1/U_1/U_1/memory[28][7] ), .Y(n11759) );
  INVX2 U11905 ( .A(\U_1/U_1/U_1/opcode[29][0] ), .Y(n11760) );
  INVX2 U11906 ( .A(\U_1/U_1/U_1/opcode[29][1] ), .Y(n11761) );
  INVX2 U11907 ( .A(\U_1/U_1/U_1/memory[29][0] ), .Y(n11762) );
  INVX2 U11908 ( .A(\U_1/U_1/U_1/memory[29][1] ), .Y(n11763) );
  INVX2 U11909 ( .A(\U_1/U_1/U_1/memory[29][2] ), .Y(n11764) );
  INVX2 U11910 ( .A(\U_1/U_1/U_1/memory[29][3] ), .Y(n11765) );
  INVX2 U11911 ( .A(\U_1/U_1/U_1/memory[29][4] ), .Y(n11766) );
  INVX2 U11912 ( .A(\U_1/U_1/U_1/memory[29][5] ), .Y(n11767) );
  INVX2 U11913 ( .A(\U_1/U_1/U_1/memory[29][6] ), .Y(n11768) );
  INVX2 U11914 ( .A(\U_1/U_1/U_1/memory[29][7] ), .Y(n11769) );
  INVX2 U11915 ( .A(\U_1/U_1/U_1/opcode[30][0] ), .Y(n11770) );
  INVX2 U11916 ( .A(\U_1/U_1/U_1/opcode[30][1] ), .Y(n11771) );
  INVX2 U11917 ( .A(\U_1/U_1/U_1/memory[30][0] ), .Y(n11772) );
  INVX2 U11918 ( .A(\U_1/U_1/U_1/memory[30][1] ), .Y(n11773) );
  INVX2 U11919 ( .A(\U_1/U_1/U_1/memory[30][2] ), .Y(n11774) );
  INVX2 U11920 ( .A(\U_1/U_1/U_1/memory[30][3] ), .Y(n11775) );
  INVX2 U11921 ( .A(\U_1/U_1/U_1/memory[30][4] ), .Y(n11776) );
  INVX2 U11922 ( .A(\U_1/U_1/U_1/memory[30][5] ), .Y(n11777) );
  INVX2 U11923 ( .A(\U_1/U_1/U_1/memory[30][6] ), .Y(n11778) );
  INVX2 U11924 ( .A(\U_1/U_1/U_1/memory[30][7] ), .Y(n11779) );
  INVX2 U11925 ( .A(\U_1/U_1/U_1/opcode[31][0] ), .Y(n11780) );
  INVX2 U11926 ( .A(\U_1/U_1/U_1/opcode[31][1] ), .Y(n11781) );
  INVX2 U11927 ( .A(\U_1/U_1/U_1/memory[31][0] ), .Y(n11782) );
  INVX2 U11928 ( .A(\U_1/U_1/U_1/memory[31][1] ), .Y(n11783) );
  INVX2 U11929 ( .A(\U_1/U_1/U_1/memory[31][2] ), .Y(n11784) );
  INVX2 U11930 ( .A(\U_1/U_1/U_1/memory[31][3] ), .Y(n11785) );
  INVX2 U11931 ( .A(\U_1/U_1/U_1/memory[31][4] ), .Y(n11786) );
  INVX2 U11932 ( .A(\U_1/U_1/U_1/memory[31][5] ), .Y(n11787) );
  INVX2 U11933 ( .A(\U_1/U_1/U_1/memory[31][6] ), .Y(n11788) );
  INVX2 U11934 ( .A(\U_1/U_1/U_1/memory[31][7] ), .Y(n11789) );
  INVX2 U11935 ( .A(\U_1/U_1/U_1/opcode[16][0] ), .Y(n11790) );
  INVX2 U11936 ( .A(\U_1/U_1/U_1/opcode[16][1] ), .Y(n11791) );
  INVX2 U11937 ( .A(\U_1/U_1/U_1/memory[16][0] ), .Y(n11792) );
  INVX2 U11938 ( .A(\U_1/U_1/U_1/memory[16][1] ), .Y(n11793) );
  INVX2 U11939 ( .A(\U_1/U_1/U_1/memory[16][2] ), .Y(n11794) );
  INVX2 U11940 ( .A(\U_1/U_1/U_1/memory[16][3] ), .Y(n11795) );
  INVX2 U11941 ( .A(\U_1/U_1/U_1/memory[16][4] ), .Y(n11796) );
  INVX2 U11942 ( .A(\U_1/U_1/U_1/memory[16][5] ), .Y(n11797) );
  INVX2 U11943 ( .A(\U_1/U_1/U_1/memory[16][6] ), .Y(n11798) );
  INVX2 U11944 ( .A(\U_1/U_1/U_1/memory[16][7] ), .Y(n11799) );
  INVX2 U11945 ( .A(\U_1/U_1/U_1/opcode[17][0] ), .Y(n11800) );
  INVX2 U11946 ( .A(\U_1/U_1/U_1/opcode[17][1] ), .Y(n11801) );
  INVX2 U11947 ( .A(\U_1/U_1/U_1/memory[17][0] ), .Y(n11802) );
  INVX2 U11948 ( .A(\U_1/U_1/U_1/memory[17][1] ), .Y(n11803) );
  INVX2 U11949 ( .A(\U_1/U_1/U_1/memory[17][2] ), .Y(n11804) );
  INVX2 U11950 ( .A(\U_1/U_1/U_1/memory[17][3] ), .Y(n11805) );
  INVX2 U11951 ( .A(\U_1/U_1/U_1/memory[17][4] ), .Y(n11806) );
  INVX2 U11952 ( .A(\U_1/U_1/U_1/memory[17][5] ), .Y(n11807) );
  INVX2 U11953 ( .A(\U_1/U_1/U_1/memory[17][6] ), .Y(n11808) );
  INVX2 U11954 ( .A(\U_1/U_1/U_1/memory[17][7] ), .Y(n11809) );
  INVX2 U11955 ( .A(\U_1/U_1/U_1/opcode[18][0] ), .Y(n11810) );
  INVX2 U11956 ( .A(\U_1/U_1/U_1/opcode[18][1] ), .Y(n11811) );
  INVX2 U11957 ( .A(\U_1/U_1/U_1/memory[18][0] ), .Y(n11812) );
  INVX2 U11958 ( .A(\U_1/U_1/U_1/memory[18][1] ), .Y(n11813) );
  INVX2 U11959 ( .A(\U_1/U_1/U_1/memory[18][2] ), .Y(n11814) );
  INVX2 U11960 ( .A(\U_1/U_1/U_1/memory[18][3] ), .Y(n11815) );
  INVX2 U11961 ( .A(\U_1/U_1/U_1/memory[18][4] ), .Y(n11816) );
  INVX2 U11962 ( .A(\U_1/U_1/U_1/memory[18][5] ), .Y(n11817) );
  INVX2 U11963 ( .A(\U_1/U_1/U_1/memory[18][6] ), .Y(n11818) );
  INVX2 U11964 ( .A(\U_1/U_1/U_1/memory[18][7] ), .Y(n11819) );
  INVX2 U11965 ( .A(\U_1/U_1/U_1/opcode[19][0] ), .Y(n11820) );
  INVX2 U11966 ( .A(\U_1/U_1/U_1/opcode[19][1] ), .Y(n11821) );
  INVX2 U11967 ( .A(\U_1/U_1/U_1/memory[19][3] ), .Y(n11822) );
  INVX2 U11968 ( .A(\U_1/U_1/U_1/memory[19][4] ), .Y(n11823) );
  INVX2 U11969 ( .A(\U_1/U_1/U_1/memory[19][5] ), .Y(n11824) );
  INVX2 U11970 ( .A(\U_1/U_1/U_1/memory[19][6] ), .Y(n11825) );
  INVX2 U11971 ( .A(\U_1/U_1/U_1/memory[19][7] ), .Y(n11826) );
  INVX2 U11972 ( .A(\U_1/U_1/U_1/memory[19][0] ), .Y(n11827) );
  INVX2 U11973 ( .A(\U_1/U_1/U_1/memory[19][1] ), .Y(n11828) );
  INVX2 U11974 ( .A(\U_1/U_1/U_1/memory[19][2] ), .Y(n11829) );
  INVX2 U11975 ( .A(n6028), .Y(n11830) );
  INVX2 U11976 ( .A(\U_1/U_1/DATA [0]), .Y(n11831) );
  INVX2 U11977 ( .A(\U_1/U_1/DATA [1]), .Y(n11832) );
  INVX2 U11978 ( .A(\U_1/U_1/DATA [2]), .Y(n11833) );
  INVX2 U11979 ( .A(\U_1/U_1/DATA [3]), .Y(n11834) );
  INVX2 U11980 ( .A(\U_1/U_1/DATA [4]), .Y(n11835) );
  INVX2 U11981 ( .A(\U_1/U_1/DATA [5]), .Y(n11836) );
  INVX2 U11982 ( .A(\U_1/U_1/DATA [6]), .Y(n11837) );
  INVX2 U11983 ( .A(\U_1/U_1/DATA [7]), .Y(n11838) );
  INVX2 U11984 ( .A(\U_1/U_1/OUT_OPCODE [0]), .Y(n11839) );
  INVX2 U11985 ( .A(\U_1/U_1/OUT_OPCODE [1]), .Y(n11840) );
  INVX2 U11986 ( .A(n6021), .Y(n11841) );
  INVX2 U11987 ( .A(\U_1/U_1/U_0/state[0] ), .Y(n11842) );
  INVX2 U11988 ( .A(\U_1/U_1/U_0/state[1] ), .Y(n11843) );
  INVX2 U11989 ( .A(\U_1/B_READY ), .Y(n11844) );
  INVX2 U11990 ( .A(n5819), .Y(n11845) );
  INVX2 U11991 ( .A(n6216), .Y(n11846) );
  INVX2 U11992 ( .A(\U_1/PRGA_OPCODE[0] ), .Y(n11847) );
  INVX2 U11993 ( .A(\U_1/U_1/U_0/tempOpcode [0]), .Y(n11848) );
  INVX2 U11994 ( .A(\U_1/U_1/U_0/tempData [7]), .Y(n11849) );
  INVX2 U11995 ( .A(\U_1/PRGA_IN [7]), .Y(n11850) );
  INVX2 U11996 ( .A(\U_1/U_1/U_0/tempData [6]), .Y(n11851) );
  INVX2 U11997 ( .A(\U_1/PRGA_IN [6]), .Y(n11852) );
  INVX2 U11998 ( .A(\U_1/U_1/U_0/tempData [5]), .Y(n11853) );
  INVX2 U11999 ( .A(\U_1/PRGA_IN [5]), .Y(n11854) );
  INVX2 U12000 ( .A(\U_1/U_1/U_0/tempData [4]), .Y(n11855) );
  INVX2 U12001 ( .A(\U_1/PRGA_IN [4]), .Y(n11856) );
  INVX2 U12002 ( .A(\U_1/U_1/U_0/tempData [3]), .Y(n11857) );
  INVX2 U12003 ( .A(\U_1/PRGA_IN [3]), .Y(n11858) );
  INVX2 U12004 ( .A(\U_1/U_1/U_0/tempData [2]), .Y(n11859) );
  INVX2 U12005 ( .A(\U_1/PRGA_IN [2]), .Y(n11860) );
  INVX2 U12006 ( .A(\U_1/U_1/U_0/tempData [1]), .Y(n11861) );
  INVX2 U12007 ( .A(\U_1/PRGA_IN [1]), .Y(n11862) );
  INVX2 U12008 ( .A(\U_1/U_1/U_0/tempData [0]), .Y(n11863) );
  INVX2 U12009 ( .A(\U_1/PRGA_IN [0]), .Y(n11864) );
  INVX2 U12010 ( .A(\U_1/PRGA_OPCODE[1] ), .Y(n11865) );
  INVX2 U12011 ( .A(\U_1/U_3/U_3/count[0] ), .Y(n11866) );
  INVX2 U12012 ( .A(\U_1/U_3/U_3/count[5] ), .Y(n11867) );
  INVX2 U12013 ( .A(n5838), .Y(n11868) );
  INVX2 U12014 ( .A(\U_1/U_3/U_3/count[1] ), .Y(n11869) );
  INVX2 U12015 ( .A(\U_1/U_3/U_3/count[2] ), .Y(n11870) );
  INVX2 U12016 ( .A(\U_1/U_3/U_3/count[3] ), .Y(n11871) );
  INVX2 U12017 ( .A(\U_1/U_3/U_3/count[4] ), .Y(n11872) );
  INVX2 U12018 ( .A(\U_1/U_0/U_0/nfaddr[0] ), .Y(n11873) );
  INVX2 U12019 ( .A(\U_1/U_0/U_0/nfaddr[1] ), .Y(n11874) );
  INVX2 U12020 ( .A(\U_1/U_0/U_0/nfaddr[2] ), .Y(n11875) );
  INVX2 U12021 ( .A(\U_1/U_0/U_0/nfaddr[3] ), .Y(n11876) );
  INVX2 U12022 ( .A(\U_1/U_0/U_0/nfaddr[4] ), .Y(n11877) );
  INVX2 U12023 ( .A(\U_1/U_0/U_0/nfaddr[5] ), .Y(n11878) );
  INVX2 U12024 ( .A(\U_1/U_0/U_0/nfaddr[6] ), .Y(n11879) );
  INVX2 U12025 ( .A(\U_1/U_0/U_0/nfaddr[7] ), .Y(n11880) );
  INVX2 U12026 ( .A(n300), .Y(n11881) );
  INVX2 U12027 ( .A(n1097), .Y(n11882) );
  INVX2 U12028 ( .A(n975), .Y(n11884) );
  INVX2 U12029 ( .A(n1090), .Y(n11885) );
  INVX2 U12030 ( .A(n6227), .Y(n11887) );
  INVX2 U12031 ( .A(n6156), .Y(n11888) );
  INVX2 U12032 ( .A(n1054), .Y(n11889) );
  INVX2 U12033 ( .A(n6272), .Y(n11890) );
  INVX2 U12034 ( .A(n981), .Y(n11891) );
  INVX2 U12035 ( .A(n301), .Y(n11893) );
  INVX2 U12036 ( .A(n6189), .Y(n11894) );
  INVX2 U12037 ( .A(n980), .Y(n11895) );
  INVX2 U12038 ( .A(n312), .Y(n11897) );
  INVX2 U12039 ( .A(n6152), .Y(n11898) );
  INVX2 U12040 ( .A(n1089), .Y(n11900) );
  INVX2 U12041 ( .A(n6165), .Y(n11901) );
  INVX2 U12042 ( .A(n6093), .Y(n11902) );
  INVX2 U12043 ( .A(n6089), .Y(n11903) );
  INVX2 U12044 ( .A(n6085), .Y(n11904) );
  INVX2 U12045 ( .A(n6081), .Y(n11905) );
  INVX2 U12046 ( .A(n6077), .Y(n11906) );
  INVX2 U12047 ( .A(n6073), .Y(n11907) );
  INVX2 U12048 ( .A(n6069), .Y(n11908) );
  INVX2 U12049 ( .A(n6063), .Y(n11909) );
  INVX2 U12050 ( .A(n921), .Y(n11910) );
  INVX2 U12051 ( .A(n1096), .Y(n11911) );
  INVX2 U12052 ( .A(n6100), .Y(n11912) );
  INVX2 U12053 ( .A(n912), .Y(n11915) );
  INVX2 U12054 ( .A(n6183), .Y(n11916) );
  INVX2 U12055 ( .A(\U_1/U_0/U_0/state[0] ), .Y(n11917) );
  INVX2 U12056 ( .A(n6221), .Y(n11919) );
  INVX2 U12057 ( .A(n6240), .Y(n11920) );
  INVX2 U12058 ( .A(n307), .Y(n11921) );
  INVX2 U12059 ( .A(n6177), .Y(n11922) );
  INVX2 U12060 ( .A(\U_1/U_0/U_0/si[0] ), .Y(n11923) );
  INVX2 U12061 ( .A(\U_1/U_0/U_0/permuteComplete ), .Y(n11924) );
  INVX2 U12062 ( .A(n6155), .Y(n11925) );
  INVX2 U12063 ( .A(\U_1/U_0/U_0/state[3] ), .Y(n11926) );
  INVX2 U12064 ( .A(n6278), .Y(n11927) );
  INVX2 U12065 ( .A(n6193), .Y(n11928) );
  INVX2 U12066 ( .A(n9196), .Y(n11929) );
  INVX2 U12067 ( .A(n9286), .Y(n11930) );
  INVX2 U12068 ( .A(\U_1/U_0/U_0/state[1] ), .Y(n11931) );
  INVX2 U12069 ( .A(\U_1/PDATA_READY ), .Y(n11932) );
  INVX2 U12070 ( .A(\U_1/U_0/U_0/state[2] ), .Y(n11933) );
  INVX2 U12071 ( .A(\U_1/U_0/U_0/prefillCounter[0] ), .Y(n11934) );
  INVX2 U12072 ( .A(\U_1/U_0/U_0/prefillCounter[1] ), .Y(n11935) );
  INVX2 U12073 ( .A(\U_1/U_0/U_0/prefillCounter[2] ), .Y(n11936) );
  INVX2 U12074 ( .A(\U_1/U_0/U_0/prefillCounter[3] ), .Y(n11937) );
  INVX2 U12075 ( .A(\U_1/U_0/U_0/prefillCounter[4] ), .Y(n11938) );
  INVX2 U12076 ( .A(\U_1/U_0/U_0/prefillCounter[5] ), .Y(n11939) );
  INVX2 U12077 ( .A(\U_1/U_0/U_0/prefillCounter[6] ), .Y(n11940) );
  INVX2 U12078 ( .A(\U_1/U_0/U_0/prefillCounter[7] ), .Y(n11941) );
  INVX2 U12079 ( .A(\U_1/U_0/U_0/keyTable[0][6] ), .Y(n11942) );
  INVX2 U12080 ( .A(\U_1/U_0/U_0/keyTable[0][5] ), .Y(n11943) );
  INVX2 U12081 ( .A(\U_1/U_0/U_0/keyTable[0][4] ), .Y(n11944) );
  INVX2 U12082 ( .A(\U_1/U_0/U_0/keyTable[0][3] ), .Y(n11945) );
  INVX2 U12083 ( .A(\U_1/U_0/U_0/keyTable[0][2] ), .Y(n11946) );
  INVX2 U12084 ( .A(\U_1/U_0/U_0/keyTable[0][1] ), .Y(n11947) );
  INVX2 U12085 ( .A(\U_1/U_0/U_0/keyTable[0][0] ), .Y(n11948) );
  INVX2 U12086 ( .A(\U_1/U_0/U_0/keyTable[1][7] ), .Y(n11949) );
  INVX2 U12087 ( .A(\U_1/U_0/U_0/keyTable[0][7] ), .Y(n11950) );
  INVX2 U12088 ( .A(\U_1/U_0/U_0/keyTable[3][0] ), .Y(n11951) );
  INVX2 U12089 ( .A(\U_1/U_0/U_0/keyTable[3][1] ), .Y(n11952) );
  INVX2 U12090 ( .A(\U_1/U_0/U_0/keyTable[3][2] ), .Y(n11953) );
  INVX2 U12091 ( .A(\U_1/U_0/U_0/keyTable[3][3] ), .Y(n11954) );
  INVX2 U12092 ( .A(\U_1/U_0/U_0/keyTable[3][4] ), .Y(n11955) );
  INVX2 U12093 ( .A(\U_1/U_0/U_0/keyTable[3][5] ), .Y(n11956) );
  INVX2 U12094 ( .A(\U_1/U_0/U_0/keyTable[3][6] ), .Y(n11957) );
  INVX2 U12095 ( .A(\U_1/U_0/U_0/keyTable[3][7] ), .Y(n11958) );
  INVX2 U12096 ( .A(\U_1/U_0/U_0/keyTable[2][0] ), .Y(n11959) );
  INVX2 U12097 ( .A(\U_1/U_0/U_0/keyTable[2][1] ), .Y(n11960) );
  INVX2 U12098 ( .A(\U_1/U_0/U_0/keyTable[2][2] ), .Y(n11961) );
  INVX2 U12099 ( .A(\U_1/U_0/U_0/keyTable[2][3] ), .Y(n11962) );
  INVX2 U12100 ( .A(\U_1/U_0/U_0/keyTable[2][4] ), .Y(n11963) );
  INVX2 U12101 ( .A(\U_1/U_0/U_0/keyTable[2][5] ), .Y(n11964) );
  INVX2 U12102 ( .A(\U_1/U_0/U_0/keyTable[2][6] ), .Y(n11965) );
  INVX2 U12103 ( .A(\U_1/U_0/U_0/keyTable[2][7] ), .Y(n11966) );
  INVX2 U12104 ( .A(\U_1/U_0/U_0/keyTable[1][0] ), .Y(n11967) );
  INVX2 U12105 ( .A(\U_1/U_0/U_0/keyTable[1][1] ), .Y(n11968) );
  INVX2 U12106 ( .A(\U_1/U_0/U_0/keyTable[1][2] ), .Y(n11969) );
  INVX2 U12107 ( .A(\U_1/U_0/U_0/keyTable[1][3] ), .Y(n11970) );
  INVX2 U12108 ( .A(\U_1/U_0/U_0/keyTable[1][4] ), .Y(n11971) );
  INVX2 U12109 ( .A(\U_1/U_0/U_0/keyTable[1][5] ), .Y(n11972) );
  INVX2 U12110 ( .A(\U_1/U_0/U_0/keyTable[1][6] ), .Y(n11973) );
  INVX2 U12111 ( .A(\U_1/U_0/U_0/si[7] ), .Y(n11974) );
  INVX2 U12112 ( .A(\U_1/U_0/U_0/si[2] ), .Y(n11975) );
  INVX2 U12113 ( .A(\U_1/U_0/U_0/si[4] ), .Y(n11976) );
  INVX2 U12114 ( .A(\U_1/U_0/U_0/si[5] ), .Y(n11977) );
  INVX2 U12115 ( .A(\U_1/U_0/U_0/si[6] ), .Y(n11978) );
  INVX2 U12116 ( .A(\U_1/U_0/U_0/keyi[2] ), .Y(n11979) );
  INVX2 U12117 ( .A(n6363), .Y(n11980) );
  INVX2 U12118 ( .A(n6364), .Y(n11981) );
  INVX2 U12119 ( .A(n6365), .Y(n11982) );
  INVX2 U12120 ( .A(n6366), .Y(n11983) );
  INVX2 U12121 ( .A(\U_1/U_0/U_0/keyi[1] ), .Y(n11984) );
  INVX2 U12122 ( .A(\U_1/U_0/U_0/sj[7] ), .Y(n11985) );
  INVX2 U12123 ( .A(\U_1/U_0/U_0/sj[6] ), .Y(n11986) );
  INVX2 U12124 ( .A(\U_1/U_0/U_0/sj[5] ), .Y(n11987) );
  INVX2 U12125 ( .A(\U_1/U_0/U_0/sj[4] ), .Y(n11988) );
  INVX2 U12126 ( .A(\U_1/U_0/U_0/sj[3] ), .Y(n11989) );
  INVX2 U12127 ( .A(\U_1/U_0/U_0/sj[2] ), .Y(n11990) );
  INVX2 U12128 ( .A(\U_1/U_0/U_0/sj[1] ), .Y(n11991) );
  INVX2 U12129 ( .A(\U_1/U_0/U_0/sj[0] ), .Y(n11992) );
  INVX2 U12130 ( .A(\U_1/U_0/U_0/N503 ), .Y(n11993) );
  INVX2 U12131 ( .A(\U_1/U_0/U_0/inti[7] ), .Y(n11994) );
  INVX2 U12132 ( .A(\U_1/U_0/U_0/N502 ), .Y(n11995) );
  INVX2 U12133 ( .A(\U_1/U_0/U_0/N501 ), .Y(n11996) );
  INVX2 U12134 ( .A(\U_1/U_0/U_0/N500 ), .Y(n11997) );
  INVX2 U12135 ( .A(\U_1/U_0/U_0/N499 ), .Y(n11998) );
  INVX2 U12136 ( .A(\U_1/U_0/U_0/N498 ), .Y(n11999) );
  INVX2 U12137 ( .A(\U_1/U_0/U_0/N497 ), .Y(n12000) );
  INVX2 U12138 ( .A(\U_1/U_0/U_0/inti[0] ), .Y(n12001) );
  INVX2 U12139 ( .A(\U_1/U_0/U_0/inti[1] ), .Y(n12002) );
  INVX2 U12140 ( .A(\U_1/U_0/U_0/inti[2] ), .Y(n12003) );
  INVX2 U12141 ( .A(\U_1/U_0/U_0/inti[3] ), .Y(n12004) );
  INVX2 U12142 ( .A(\U_1/U_0/U_0/inti[4] ), .Y(n12005) );
  INVX2 U12143 ( .A(\U_1/U_0/U_0/inti[5] ), .Y(n12006) );
  INVX2 U12144 ( .A(\U_1/U_0/U_0/inti[6] ), .Y(n12007) );
  INVX2 U12145 ( .A(\U_1/U_0/U_0/intj[0] ), .Y(n12008) );
  INVX2 U12146 ( .A(\U_1/U_0/U_0/intj[1] ), .Y(n12009) );
  INVX2 U12147 ( .A(\U_1/U_0/U_0/intj[2] ), .Y(n12010) );
  INVX2 U12148 ( .A(\U_1/U_0/U_0/intj[3] ), .Y(n12011) );
  INVX2 U12149 ( .A(\U_1/U_0/U_0/intj[4] ), .Y(n12012) );
  INVX2 U12150 ( .A(\U_1/U_0/U_0/intj[5] ), .Y(n12013) );
  INVX2 U12151 ( .A(\U_1/U_0/U_0/intj[6] ), .Y(n12014) );
  INVX2 U12152 ( .A(\U_1/U_0/U_0/intj[7] ), .Y(n12015) );
  INVX2 U12153 ( .A(\U_1/U_0/U_0/temp[0] ), .Y(n12016) );
  INVX2 U12154 ( .A(\U_1/U_0/U_0/currentProcessedData [0]), .Y(n12017) );
  INVX2 U12155 ( .A(\U_1/U_0/U_0/temp[1] ), .Y(n12018) );
  INVX2 U12156 ( .A(\U_1/U_0/U_0/currentProcessedData [1]), .Y(n12019) );
  INVX2 U12157 ( .A(\U_1/U_0/U_0/temp[2] ), .Y(n12020) );
  INVX2 U12158 ( .A(\U_1/U_0/U_0/currentProcessedData [2]), .Y(n12021) );
  INVX2 U12159 ( .A(\U_1/U_0/U_0/temp[3] ), .Y(n12022) );
  INVX2 U12160 ( .A(\U_1/U_0/U_0/currentProcessedData [3]), .Y(n12023) );
  INVX2 U12161 ( .A(\U_1/U_0/U_0/temp[4] ), .Y(n12024) );
  INVX2 U12162 ( .A(\U_1/U_0/U_0/currentProcessedData [4]), .Y(n12025) );
  INVX2 U12163 ( .A(\U_1/PROCESSED_DATA [4]), .Y(n12026) );
  INVX2 U12164 ( .A(\U_1/U_0/U_0/temp[5] ), .Y(n12027) );
  INVX2 U12165 ( .A(\U_1/U_0/U_0/currentProcessedData [5]), .Y(n12028) );
  INVX2 U12166 ( .A(n839), .Y(n12029) );
  INVX2 U12167 ( .A(\U_1/U_0/U_0/temp[6] ), .Y(n12030) );
  INVX2 U12168 ( .A(\U_1/U_0/U_0/currentProcessedData [6]), .Y(n12031) );
  INVX2 U12169 ( .A(\U_1/PROCESSED_DATA [6]), .Y(n12032) );
  INVX2 U12170 ( .A(\U_1/U_0/U_0/temp[7] ), .Y(n12033) );
  INVX2 U12171 ( .A(\U_1/U_0/U_0/currentProcessedData [7]), .Y(n12034) );
  INVX2 U12172 ( .A(\U_1/PROCESSED_DATA [7]), .Y(n12035) );
  INVX2 U12173 ( .A(\U_1/U_3/TX_CRC [0]), .Y(n12036) );
  INVX2 U12174 ( .A(\U_1/U_3/TX_CRC [8]), .Y(n12037) );
  INVX2 U12175 ( .A(\U_1/U_3/TX_CRC [2]), .Y(n12038) );
  INVX2 U12176 ( .A(\U_1/U_3/TX_CRC [10]), .Y(n12039) );
  INVX2 U12177 ( .A(\U_1/U_3/TX_CRC [3]), .Y(n12040) );
  INVX2 U12178 ( .A(\U_1/U_3/TX_CRC [11]), .Y(n12041) );
  INVX2 U12179 ( .A(\U_1/U_3/TX_CRC [4]), .Y(n12042) );
  INVX2 U12180 ( .A(\U_1/U_3/TX_CRC [12]), .Y(n12043) );
  INVX2 U12181 ( .A(\U_1/U_3/TX_CRC [5]), .Y(n12044) );
  INVX2 U12182 ( .A(\U_1/U_3/TX_CRC [13]), .Y(n12045) );
  INVX2 U12183 ( .A(\U_1/U_3/TX_CRC [6]), .Y(n12046) );
  INVX2 U12184 ( .A(\U_1/U_3/TX_CRC [14]), .Y(n12047) );
  INVX2 U12185 ( .A(\U_1/U_3/TX_CRC [7]), .Y(n12048) );
  INVX2 U12186 ( .A(\U_1/U_3/TX_CRC [15]), .Y(n12049) );
  INVX2 U12187 ( .A(\U_1/U_3/TX_CRC [1]), .Y(n12050) );
  INVX2 U12188 ( .A(\U_1/U_3/TX_CRC [9]), .Y(n12051) );
  INVX2 U12189 ( .A(\U_1/U_0/U_0/keyi[0] ), .Y(n12052) );
  INVX2 U12190 ( .A(\U_1/U_1/U_0/tempOpcode [1]), .Y(n12053) );
  INVX2 U12191 ( .A(\U_1/U_3/U_3/flop_data [7]), .Y(n12054) );
  INVX2 U12192 ( .A(\U_1/U_3/U_3/current_send_data [6]), .Y(n12055) );
  INVX2 U12193 ( .A(\U_1/U_3/send_data [6]), .Y(n12056) );
  INVX2 U12194 ( .A(\U_1/U_3/U_3/current_send_data [5]), .Y(n12057) );
  INVX2 U12195 ( .A(\U_1/U_3/send_data [5]), .Y(n12058) );
  INVX2 U12196 ( .A(\U_1/U_3/U_3/current_send_data [4]), .Y(n12059) );
  INVX2 U12197 ( .A(\U_1/U_3/send_data [4]), .Y(n12060) );
  INVX2 U12198 ( .A(\U_1/U_3/U_3/current_send_data [3]), .Y(n12061) );
  INVX2 U12199 ( .A(\U_1/U_3/send_data [3]), .Y(n12062) );
  INVX2 U12200 ( .A(\U_1/U_3/U_3/current_send_data [2]), .Y(n12063) );
  INVX2 U12201 ( .A(\U_1/U_3/send_data [2]), .Y(n12064) );
  INVX2 U12202 ( .A(\U_1/U_3/U_3/current_send_data [1]), .Y(n12065) );
  INVX2 U12203 ( .A(\U_1/U_3/send_data [1]), .Y(n12066) );
  INVX2 U12204 ( .A(\U_1/U_3/U_3/current_send_data [0]), .Y(n12067) );
  INVX2 U12205 ( .A(\U_1/U_3/send_data [0]), .Y(n12068) );
  INVX2 U12206 ( .A(\U_1/U_3/U_3/current_send_data [7]), .Y(n12069) );
  INVX2 U12207 ( .A(\U_1/U_3/U_4/count[0] ), .Y(n12070) );
  INVX2 U12208 ( .A(\U_1/U_3/U_4/count[2] ), .Y(n12071) );
  INVX2 U12209 ( .A(\U_1/U_3/U_4/count[1] ), .Y(n12072) );
  INVX2 U12210 ( .A(\U_1/U_3/U_2/count[1] ), .Y(n12073) );
  INVX2 U12211 ( .A(\U_1/U_3/U_2/count[2] ), .Y(n12074) );
  INVX2 U12212 ( .A(\U_1/U_3/U_2/count[0] ), .Y(n12075) );
  INVX2 U12213 ( .A(\U_1/U_3/d_encode ), .Y(n12076) );
  INVX2 U12214 ( .A(\U_1/U_3/U_0/DE_holdout_BS ), .Y(n12077) );
endmodule

module  rmedt_square ( CLK, DPHS, DMHS, DPSS, DMSS, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN, BSE_H, BSE_S, CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, c_parity_error, c_prog_error, host_is_sending, slave_is_sending);

input   CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN;
output  BSE_H, BSE_S, CRCE_H, CRCE_S, EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, c_parity_error, c_prog_error, host_is_sending, slave_is_sending, DMTH, DMTS, DPTH, DPTS;
inout   DPHS, DMHS, DPSS, DMSS;
wire    nCLK, nDMRH, nDMRS, nDPRH, nDPRS, nRST, nSERIAL_IN, nBSE_H, nBSE_S, nCRCE_H, nCRCE_S, nDMTH, nDMTS, nDPTH, nDPTS, nEMPTY_H, nEMPTY_S, nFULL_H, nFULL_S, nRE_H, nRE_S, nc_key_error, nc_parity_error, nc_prog_error, nhost_is_sending, nslave_is_sending;

        rmedt_square_t I0 ( .CLK(nCLK), .DMRH(nDMRH), .DMRS(nDMRS), .DPRH(nDPRH),
    .DPRS(nDPRS), .RST(nRST), .SERIAL_IN(nSERIAL_IN), .BSE_H(nBSE_H), .BSE_S(nBSE_S),
    .CRCE_H(nCRCE_H), .CRCE_S(nCRCE_S), .DMTH(nDMTH), .DMTS(nDMTS),
    .DPTH(nDPTH), .DPTS(nDPTS), .EMPTY_H(nEMPTY_H), .EMPTY_S(nSERIAL_IN),
    .FULL_H(nFULL_H), .FULL_S(nFULL_S), .RE_H(nRE_H), .RE_S(nRE_S),
    .c_key_error(nc_key_error), .c_parity_error(nc_parity_error), .c_prog_error(nc_prog_error), .host_is_sending(nhost_is_sending),
    .slave_is_sending(nslave_is_sending));

PADVDD U1 (  );
PADGND U2 (  );
PADINC U3 ( .DI(nCLK), .YPAD(CLK) );
PADINC U8 ( .DI(nRST), .YPAD(RST) );
PADINC U9 ( .DI(nSERIAL_IN), .YPAD(SERIAL_IN) );
PADINOUT UIO1 ( .DI(nDPRH), .DO(nDPTH), .OEN(nslave_is_sending), .YPAD(DPHS));
PADINOUT UIO2 ( .DI(nDMRH), .DO(nDMTH), .OEN(nslave_is_sending), .YPAD(DMHS));
PADINOUT UIO3 ( .DI(nDPRS), .DO(nDPTS), .OEN(nhost_is_sending), .YPAD(DPSS));
PADINOUT UIO4 ( .DI(nDMRS), .DO(nDMTS), .OEN(nhost_is_sending), .YPAD(DMSS));
PADOUT UOUT1 ( .DO(BSE_H), .YPAD(nBSE_H) );
PADOUT UOUT2 ( .DO(BSE_S), .YPAD(nBSE_S) );
PADOUT UOUT3 ( .DO(CRCE_H), .YPAD(nCRCE_H) );
PADOUT UOUT4 ( .DO(CRCE_S), .YPAD(nCRCE_S) );
PADOUT UOUT5 ( .DO(EMPTY_H), .YPAD(nEMPTY_H) );
PADOUT UOUT6 ( .DO(EMPTY_S), .YPAD(nEMPTY_S) );
PADOUT UOUT7 ( .DO(FULL_H), .YPAD(nFULL_H) );
PADOUT UOUT8 ( .DO(FULL_S), .YPAD(nFULL_S) );
PADOUT UOUT9 ( .DO(RE_H), .YPAD(nRE_H) );
PADOUT UOUT10 ( .DO(RE_S), .YPAD(nRE_S) );
PADOUT UOUT11 ( .DO(c_key_error), .YPAD(nc_key_error) );
PADOUT UOUT12 ( .DO(c_parity_error), .YPAD(nc_parity_error) );
PADOUT UOUT13 ( .DO(c_prog_error), .YPAD(nc_prog_error) );

endmodule
