
module KSA_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module KSA_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module KSA_1_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_1_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_1_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_1_DW01_add_3 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [7:1] carry;

  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n6), .YC(carry[2]), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(B[3]), .B(A[3]), .Y(n1) );
  XOR2X1 U2 ( .A(carry[3]), .B(n1), .Y(SUM[3]) );
  NAND2X1 U3 ( .A(carry[3]), .B(B[3]), .Y(n2) );
  NAND2X1 U4 ( .A(carry[3]), .B(A[3]), .Y(n3) );
  NAND2X1 U5 ( .A(B[3]), .B(A[3]), .Y(n4) );
  NAND3X1 U6 ( .A(n3), .B(n2), .C(n4), .Y(carry[4]) );
  XOR2X1 U7 ( .A(B[7]), .B(A[7]), .Y(n5) );
  XOR2X1 U8 ( .A(carry[7]), .B(n5), .Y(SUM[7]) );
  AND2X2 U9 ( .A(B[0]), .B(A[0]), .Y(n6) );
  XOR2X1 U10 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module KSA_1_DW01_add_2 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(A[5]), .B(B[5]), .Y(n2) );
  XOR2X1 U3 ( .A(n2), .B(carry[5]), .Y(SUM[5]) );
  NAND2X1 U4 ( .A(A[5]), .B(B[5]), .Y(n3) );
  NAND2X1 U5 ( .A(A[5]), .B(carry[5]), .Y(n4) );
  NAND2X1 U6 ( .A(B[5]), .B(carry[5]), .Y(n5) );
  NAND3X1 U7 ( .A(n3), .B(n4), .C(n5), .Y(carry[6]) );
  XOR2X1 U8 ( .A(A[6]), .B(B[6]), .Y(n6) );
  XOR2X1 U9 ( .A(n6), .B(carry[6]), .Y(SUM[6]) );
  NAND2X1 U10 ( .A(A[6]), .B(B[6]), .Y(n7) );
  NAND2X1 U11 ( .A(A[6]), .B(carry[6]), .Y(n8) );
  NAND2X1 U12 ( .A(B[6]), .B(carry[6]), .Y(n9) );
  NAND3X1 U13 ( .A(n7), .B(n8), .C(n9), .Y(carry[7]) );
  XOR2X1 U14 ( .A(B[1]), .B(A[1]), .Y(n10) );
  XOR2X1 U15 ( .A(n1), .B(n10), .Y(SUM[1]) );
  NAND2X1 U16 ( .A(n1), .B(B[1]), .Y(n11) );
  NAND2X1 U17 ( .A(n1), .B(A[1]), .Y(n12) );
  NAND2X1 U18 ( .A(B[1]), .B(A[1]), .Y(n13) );
  NAND3X1 U19 ( .A(n12), .B(n11), .C(n13), .Y(carry[2]) );
  XOR2X1 U20 ( .A(A[2]), .B(B[2]), .Y(n14) );
  XOR2X1 U21 ( .A(n14), .B(carry[2]), .Y(SUM[2]) );
  NAND2X1 U22 ( .A(A[2]), .B(B[2]), .Y(n15) );
  NAND2X1 U23 ( .A(A[2]), .B(carry[2]), .Y(n16) );
  NAND2X1 U24 ( .A(B[2]), .B(carry[2]), .Y(n17) );
  NAND3X1 U25 ( .A(n15), .B(n16), .C(n17), .Y(carry[3]) );
  XOR2X1 U26 ( .A(A[3]), .B(B[3]), .Y(n18) );
  XOR2X1 U27 ( .A(n18), .B(carry[3]), .Y(SUM[3]) );
  NAND2X1 U28 ( .A(A[3]), .B(B[3]), .Y(n19) );
  NAND2X1 U29 ( .A(A[3]), .B(carry[3]), .Y(n20) );
  NAND2X1 U30 ( .A(B[3]), .B(carry[3]), .Y(n21) );
  NAND3X1 U31 ( .A(n19), .B(n20), .C(n21), .Y(carry[4]) );
  XOR2X1 U32 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module KSA_1 ( KEY, CLK, RST, KEY_ERROR, BYTE_READY, BYTE, OPCODE, DATA_IN, 
        PROCESSED_DATA, PDATA_READY, W_ENABLE, R_ENABLE, ADDR, DATA );
  input [63:0] KEY;
  input [7:0] BYTE;
  input [1:0] OPCODE;
  input [7:0] DATA_IN;
  output [7:0] PROCESSED_DATA;
  output [7:0] ADDR;
  output [7:0] DATA;
  input CLK, RST, KEY_ERROR, BYTE_READY;
  output PDATA_READY, W_ENABLE, R_ENABLE;
  wire   permuteComplete, \keyTable[0][7] , \keyTable[0][6] , \keyTable[0][5] ,
         \keyTable[0][4] , \keyTable[0][3] , \keyTable[0][2] ,
         \keyTable[0][1] , \keyTable[0][0] , \keyTable[1][7] ,
         \keyTable[1][6] , \keyTable[1][5] , \keyTable[1][4] ,
         \keyTable[1][3] , \keyTable[1][2] , \keyTable[1][1] ,
         \keyTable[1][0] , \keyTable[2][7] , \keyTable[2][6] ,
         \keyTable[2][5] , \keyTable[2][4] , \keyTable[2][3] ,
         \keyTable[2][2] , \keyTable[2][1] , \keyTable[2][0] ,
         \keyTable[3][7] , \keyTable[3][6] , \keyTable[3][5] ,
         \keyTable[3][4] , \keyTable[3][3] , \keyTable[3][2] ,
         \keyTable[3][1] , \keyTable[3][0] , \keyTable[4][7] ,
         \keyTable[4][6] , \keyTable[4][5] , \keyTable[4][4] ,
         \keyTable[4][3] , \keyTable[4][2] , \keyTable[4][1] ,
         \keyTable[4][0] , \keyTable[5][7] , \keyTable[5][6] ,
         \keyTable[5][5] , \keyTable[5][4] , \keyTable[5][3] ,
         \keyTable[5][2] , \keyTable[5][1] , \keyTable[5][0] ,
         \keyTable[6][7] , \keyTable[6][6] , \keyTable[6][5] ,
         \keyTable[6][4] , \keyTable[6][3] , \keyTable[6][2] ,
         \keyTable[6][1] , \keyTable[6][0] , \keyTable[7][7] ,
         \keyTable[7][6] , \keyTable[7][5] , \keyTable[7][4] ,
         \keyTable[7][3] , \keyTable[7][2] , \keyTable[7][1] ,
         \keyTable[7][0] , fw_enable, fr_enable, N407, N408, N409, N410, N411,
         N412, N413, N414, N424, N425, N426, N427, N428, N429, N430, N431,
         N442, N443, N444, N445, N446, N447, N448, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N496, N497, N498, N499, N500, N501, N502, N503, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, n11, n13, n18, n21, n23, n25, n26, n28, n30, n31,
         n33, n35, n36, n38, n40, n41, n43, n45, n46, n48, n50, n51, n53, n55,
         n56, n57, n58, n59, n60, n61, n63, n65, n66, n67, n68, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n123, n124, n125,
         n126, n127, n128, n130, n132, n133, n134, n137, n138, n139, n140,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n152, n153,
         n154, n155, n156, n157, n158, n159, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n173, n174, n176, n178, n179, n181,
         n182, n183, n184, n186, n189, n190, n191, n192, n193, n194, n195,
         n197, n198, n199, n200, n202, n204, n205, n207, n209, n211, n213,
         n215, n217, n219, n221, n222, n223, n224, n225, n226, n227, n229,
         n231, n232, n233, n234, n236, n242, n243, n245, n248, n251, n254,
         n257, n260, n263, n266, n269, n272, n273, n274, n276, n278, n279,
         n281, n283, n284, n286, n288, n289, n291, n293, n294, n296, n298,
         n299, n301, n303, n304, n306, n308, n309, n310, n312, n313, n314,
         n315, n316, n319, n320, n321, n322, n323, n324, n325, n328, n330,
         n332, n334, n336, n338, n340, n342, n344, n346, n348, n350, n352,
         n354, n356, n358, n360, n362, n364, n366, n368, n370, n372, n374,
         n376, n378, n380, n382, n384, n386, n388, n390, n392, n394, n396,
         n398, n400, n402, n404, n406, n408, n410, n412, n414, n416, n418,
         n420, n422, n424, n426, n428, n430, n432, n434, n436, n438, n440,
         n442, n444, n446, n448, n450, n452, n454, n456, n457, n460, n464,
         n466, n468, n470, n472, n474, n476, n477, n478, n479, n481, n483,
         n484, n485, n486, n487, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n499, n502, n508, n510, n511, n513, n515, n517, n519,
         n521, n523, n525, n526, n527, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n544, n546, n548, n550, n552, n554,
         n556, n558, n559, n560, n561, n563, n564, n565, n566, n567, n568,
         n570, n573, n574, n576, n578, n580, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n593, n595, n596, n597, n598, n599,
         n601, n602, n603, n607, n608, n609, n611, n613, n615, n617, n619,
         n620, n621, n622, n623, n625, n627, n628, n631, n633, n634, n635,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n693, n694, n695, n696, n697, n698,
         n699, n700, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n747, n749, n751, n753, n755, n757, n759, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, N456, N455, N454, N453,
         N452, N451, N450, N449, n3, n4, n5, n6, n7, n8, n9, n10, n12, n14,
         n15, n16, n161, n172, n175, n177, n180, n185, n187, n188, n196, n201,
         n203, n206, n208, n210, n212, n214, n216, n218, n220, n228, n230,
         n235, n237, n238, n239, n240, n241, n244, n246, n247, n249, n250,
         n252, n253, n255, n256, n258, n259, n261, n262, n264, n265, n267,
         n268, n270, n271, n275, n277, n280, n282, n285, n287, n290, n292,
         n295, n297, n300, n302, n305, n307, n311, n317, n318, n326, n327,
         n329, n331, n333, n335, n337, n339, n341, n343, n345, n347, n349,
         n351, n353, n355, n357, n359, n361, n363, n365, n367, n369, n371,
         n373, n375, n377, n379, n381, n383, n385, n387, n389, n391, n393,
         n395, n397, n399, n401, n403, n405, n407, n409, n411, n413, n415,
         n417, n419, n421, n423, n425, n427, n429, n431, n433, n435, n437,
         n439, n441, n443, n445, n447, n449, n451, n453, n455, n458, n459,
         n461, n462, n463, n465, n467, n469, n471, n473, n475, n480, n482,
         n488, n498, n500, n501, n503, n504, n505, n506, n507, n509, n512,
         n514, n516, n518, n520, n522, n524, n528, n540, n541, n542, n543,
         n545, n547, n549, n551, n553, n555, n557, n562, n569, n571, n572,
         n575, n577, n579, n581, n592, n594, n600, n604, n605, n606, n610,
         n612, n614, n616, n618, n624, n626, n629, n630, n632, n636, n637,
         n638, n648, n649, n650, n651, n692, n701, n746, n748, n750, n752,
         n754, n756, n758, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n864, n865, n866, n867, n868, n869, n870, n871, n883,
         n884, n885, n886, n887, n888, n889, n890, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975;
  wire   [4:0] state;
  wire   [7:0] si;
  wire   [7:0] sj;
  wire   [7:0] currentProcessedData;
  wire   [4:0] nextState;
  wire   [7:0] inti;
  wire   [7:0] intj;
  wire   [2:0] keyi;
  wire   [7:0] temp;
  wire   [7:0] extratemp;
  wire   [7:0] nextProcessedData;
  wire   [7:0] delaydata;
  wire   [7:0] prefillCounter;
  wire   [7:0] faddr;
  wire   [7:0] fdata;
  tri   [7:0] nfaddr;
  tri   [7:0] nfdata;

  DFFPOSX1 \prefillCounter_reg[0]  ( .D(n915), .CLK(CLK), .Q(prefillCounter[0]) );
  DFFPOSX1 permuteComplete_reg ( .D(n899), .CLK(CLK), .Q(permuteComplete) );
  DFFPOSX1 \extratemp_reg[7]  ( .D(n465), .CLK(CLK), .Q(extratemp[7]) );
  DFFPOSX1 \extratemp_reg[6]  ( .D(n463), .CLK(CLK), .Q(extratemp[6]) );
  DFFPOSX1 \extratemp_reg[5]  ( .D(n462), .CLK(CLK), .Q(extratemp[5]) );
  DFFPOSX1 \extratemp_reg[4]  ( .D(n461), .CLK(CLK), .Q(extratemp[4]) );
  DFFPOSX1 \extratemp_reg[3]  ( .D(n459), .CLK(CLK), .Q(extratemp[3]) );
  DFFPOSX1 \extratemp_reg[2]  ( .D(n458), .CLK(CLK), .Q(extratemp[2]) );
  DFFPOSX1 \extratemp_reg[1]  ( .D(n455), .CLK(CLK), .Q(extratemp[1]) );
  DFFPOSX1 \extratemp_reg[0]  ( .D(n453), .CLK(CLK), .Q(extratemp[0]) );
  DFFPOSX1 \keyTable_reg[7][0]  ( .D(n792), .CLK(CLK), .Q(\keyTable[7][0] ) );
  DFFPOSX1 \keyTable_reg[7][1]  ( .D(n793), .CLK(CLK), .Q(\keyTable[7][1] ) );
  DFFPOSX1 \keyTable_reg[7][2]  ( .D(n794), .CLK(CLK), .Q(\keyTable[7][2] ) );
  DFFPOSX1 \keyTable_reg[7][3]  ( .D(n795), .CLK(CLK), .Q(\keyTable[7][3] ) );
  DFFPOSX1 \keyTable_reg[7][4]  ( .D(n796), .CLK(CLK), .Q(\keyTable[7][4] ) );
  DFFPOSX1 \keyTable_reg[7][5]  ( .D(n797), .CLK(CLK), .Q(\keyTable[7][5] ) );
  DFFPOSX1 \keyTable_reg[7][6]  ( .D(n798), .CLK(CLK), .Q(\keyTable[7][6] ) );
  DFFPOSX1 \keyTable_reg[7][7]  ( .D(n799), .CLK(CLK), .Q(\keyTable[7][7] ) );
  DFFPOSX1 \keyTable_reg[6][0]  ( .D(n800), .CLK(CLK), .Q(\keyTable[6][0] ) );
  DFFPOSX1 \keyTable_reg[6][1]  ( .D(n801), .CLK(CLK), .Q(\keyTable[6][1] ) );
  DFFPOSX1 \keyTable_reg[6][2]  ( .D(n802), .CLK(CLK), .Q(\keyTable[6][2] ) );
  DFFPOSX1 \keyTable_reg[6][3]  ( .D(n803), .CLK(CLK), .Q(\keyTable[6][3] ) );
  DFFPOSX1 \keyTable_reg[6][4]  ( .D(n804), .CLK(CLK), .Q(\keyTable[6][4] ) );
  DFFPOSX1 \keyTable_reg[6][5]  ( .D(n805), .CLK(CLK), .Q(\keyTable[6][5] ) );
  DFFPOSX1 \keyTable_reg[6][6]  ( .D(n806), .CLK(CLK), .Q(\keyTable[6][6] ) );
  DFFPOSX1 \keyTable_reg[6][7]  ( .D(n807), .CLK(CLK), .Q(\keyTable[6][7] ) );
  DFFPOSX1 \keyTable_reg[5][0]  ( .D(n808), .CLK(CLK), .Q(\keyTable[5][0] ) );
  DFFPOSX1 \keyTable_reg[5][1]  ( .D(n809), .CLK(CLK), .Q(\keyTable[5][1] ) );
  DFFPOSX1 \keyTable_reg[5][2]  ( .D(n810), .CLK(CLK), .Q(\keyTable[5][2] ) );
  DFFPOSX1 \keyTable_reg[5][3]  ( .D(n811), .CLK(CLK), .Q(\keyTable[5][3] ) );
  DFFPOSX1 \keyTable_reg[5][4]  ( .D(n812), .CLK(CLK), .Q(\keyTable[5][4] ) );
  DFFPOSX1 \keyTable_reg[5][5]  ( .D(n813), .CLK(CLK), .Q(\keyTable[5][5] ) );
  DFFPOSX1 \keyTable_reg[5][6]  ( .D(n814), .CLK(CLK), .Q(\keyTable[5][6] ) );
  DFFPOSX1 \keyTable_reg[5][7]  ( .D(n815), .CLK(CLK), .Q(\keyTable[5][7] ) );
  DFFPOSX1 \keyTable_reg[4][0]  ( .D(n816), .CLK(CLK), .Q(\keyTable[4][0] ) );
  DFFPOSX1 \keyTable_reg[4][1]  ( .D(n817), .CLK(CLK), .Q(\keyTable[4][1] ) );
  DFFPOSX1 \keyTable_reg[4][2]  ( .D(n818), .CLK(CLK), .Q(\keyTable[4][2] ) );
  DFFPOSX1 \keyTable_reg[4][3]  ( .D(n819), .CLK(CLK), .Q(\keyTable[4][3] ) );
  DFFPOSX1 \keyTable_reg[4][4]  ( .D(n820), .CLK(CLK), .Q(\keyTable[4][4] ) );
  DFFPOSX1 \keyTable_reg[4][5]  ( .D(n821), .CLK(CLK), .Q(\keyTable[4][5] ) );
  DFFPOSX1 \keyTable_reg[4][6]  ( .D(n822), .CLK(CLK), .Q(\keyTable[4][6] ) );
  DFFPOSX1 \keyTable_reg[4][7]  ( .D(n823), .CLK(CLK), .Q(\keyTable[4][7] ) );
  DFFPOSX1 \keyTable_reg[3][0]  ( .D(n824), .CLK(CLK), .Q(\keyTable[3][0] ) );
  DFFPOSX1 \keyTable_reg[3][1]  ( .D(n825), .CLK(CLK), .Q(\keyTable[3][1] ) );
  DFFPOSX1 \keyTable_reg[3][2]  ( .D(n826), .CLK(CLK), .Q(\keyTable[3][2] ) );
  DFFPOSX1 \keyTable_reg[3][3]  ( .D(n827), .CLK(CLK), .Q(\keyTable[3][3] ) );
  DFFPOSX1 \keyTable_reg[3][4]  ( .D(n828), .CLK(CLK), .Q(\keyTable[3][4] ) );
  DFFPOSX1 \keyTable_reg[3][5]  ( .D(n829), .CLK(CLK), .Q(\keyTable[3][5] ) );
  DFFPOSX1 \keyTable_reg[3][6]  ( .D(n830), .CLK(CLK), .Q(\keyTable[3][6] ) );
  DFFPOSX1 \keyTable_reg[3][7]  ( .D(n831), .CLK(CLK), .Q(\keyTable[3][7] ) );
  DFFPOSX1 \keyTable_reg[2][0]  ( .D(n832), .CLK(CLK), .Q(\keyTable[2][0] ) );
  DFFPOSX1 \keyTable_reg[2][1]  ( .D(n833), .CLK(CLK), .Q(\keyTable[2][1] ) );
  DFFPOSX1 \keyTable_reg[2][2]  ( .D(n834), .CLK(CLK), .Q(\keyTable[2][2] ) );
  DFFPOSX1 \keyTable_reg[2][3]  ( .D(n835), .CLK(CLK), .Q(\keyTable[2][3] ) );
  DFFPOSX1 \keyTable_reg[2][4]  ( .D(n836), .CLK(CLK), .Q(\keyTable[2][4] ) );
  DFFPOSX1 \keyTable_reg[2][5]  ( .D(n837), .CLK(CLK), .Q(\keyTable[2][5] ) );
  DFFPOSX1 \keyTable_reg[2][6]  ( .D(n838), .CLK(CLK), .Q(\keyTable[2][6] ) );
  DFFPOSX1 \keyTable_reg[2][7]  ( .D(n839), .CLK(CLK), .Q(\keyTable[2][7] ) );
  DFFPOSX1 \keyTable_reg[1][0]  ( .D(n840), .CLK(CLK), .Q(\keyTable[1][0] ) );
  DFFPOSX1 \keyTable_reg[1][1]  ( .D(n841), .CLK(CLK), .Q(\keyTable[1][1] ) );
  DFFPOSX1 \keyTable_reg[1][2]  ( .D(n842), .CLK(CLK), .Q(\keyTable[1][2] ) );
  DFFPOSX1 \keyTable_reg[1][3]  ( .D(n843), .CLK(CLK), .Q(\keyTable[1][3] ) );
  DFFPOSX1 \keyTable_reg[1][4]  ( .D(n844), .CLK(CLK), .Q(\keyTable[1][4] ) );
  DFFPOSX1 \keyTable_reg[1][5]  ( .D(n845), .CLK(CLK), .Q(\keyTable[1][5] ) );
  DFFPOSX1 \keyTable_reg[1][6]  ( .D(n846), .CLK(CLK), .Q(\keyTable[1][6] ) );
  DFFPOSX1 \keyTable_reg[0][6]  ( .D(n847), .CLK(CLK), .Q(\keyTable[0][6] ) );
  DFFPOSX1 \keyTable_reg[0][5]  ( .D(n848), .CLK(CLK), .Q(\keyTable[0][5] ) );
  DFFPOSX1 \keyTable_reg[0][4]  ( .D(n849), .CLK(CLK), .Q(\keyTable[0][4] ) );
  DFFPOSX1 \keyTable_reg[0][3]  ( .D(n850), .CLK(CLK), .Q(\keyTable[0][3] ) );
  DFFPOSX1 \keyTable_reg[0][2]  ( .D(n851), .CLK(CLK), .Q(\keyTable[0][2] ) );
  DFFPOSX1 \keyTable_reg[0][1]  ( .D(n852), .CLK(CLK), .Q(\keyTable[0][1] ) );
  DFFPOSX1 \keyTable_reg[0][0]  ( .D(n853), .CLK(CLK), .Q(\keyTable[0][0] ) );
  DFFPOSX1 \keyTable_reg[1][7]  ( .D(n854), .CLK(CLK), .Q(\keyTable[1][7] ) );
  DFFPOSX1 \keyTable_reg[0][7]  ( .D(n855), .CLK(CLK), .Q(\keyTable[0][7] ) );
  DFFPOSX1 \prefillCounter_reg[7]  ( .D(n914), .CLK(CLK), .Q(prefillCounter[7]) );
  DFFPOSX1 \prefillCounter_reg[1]  ( .D(n913), .CLK(CLK), .Q(prefillCounter[1]) );
  DFFPOSX1 \prefillCounter_reg[2]  ( .D(n912), .CLK(CLK), .Q(prefillCounter[2]) );
  DFFPOSX1 \prefillCounter_reg[3]  ( .D(n911), .CLK(CLK), .Q(prefillCounter[3]) );
  DFFPOSX1 \prefillCounter_reg[4]  ( .D(n910), .CLK(CLK), .Q(prefillCounter[4]) );
  DFFPOSX1 \prefillCounter_reg[5]  ( .D(n909), .CLK(CLK), .Q(prefillCounter[5]) );
  DFFPOSX1 \prefillCounter_reg[6]  ( .D(n908), .CLK(CLK), .Q(prefillCounter[6]) );
  DFFPOSX1 \temp_reg[7]  ( .D(n856), .CLK(CLK), .Q(temp[7]) );
  DFFPOSX1 \temp_reg[0]  ( .D(n863), .CLK(CLK), .Q(temp[0]) );
  DFFPOSX1 \temp_reg[1]  ( .D(n862), .CLK(CLK), .Q(temp[1]) );
  DFFPOSX1 \temp_reg[2]  ( .D(n861), .CLK(CLK), .Q(temp[2]) );
  DFFPOSX1 \temp_reg[3]  ( .D(n860), .CLK(CLK), .Q(temp[3]) );
  DFFPOSX1 \temp_reg[4]  ( .D(n859), .CLK(CLK), .Q(temp[4]) );
  DFFPOSX1 \temp_reg[5]  ( .D(n858), .CLK(CLK), .Q(temp[5]) );
  DFFPOSX1 \temp_reg[6]  ( .D(n857), .CLK(CLK), .Q(temp[6]) );
  DFFPOSX1 \delaydata_reg[7]  ( .D(n371), .CLK(CLK), .Q(delaydata[7]) );
  DFFPOSX1 \delaydata_reg[0]  ( .D(n399), .CLK(CLK), .Q(delaydata[0]) );
  DFFPOSX1 \delaydata_reg[1]  ( .D(n395), .CLK(CLK), .Q(delaydata[1]) );
  DFFPOSX1 \delaydata_reg[2]  ( .D(n391), .CLK(CLK), .Q(delaydata[2]) );
  DFFPOSX1 \delaydata_reg[3]  ( .D(n387), .CLK(CLK), .Q(delaydata[3]) );
  DFFPOSX1 \delaydata_reg[4]  ( .D(n383), .CLK(CLK), .Q(delaydata[4]) );
  DFFPOSX1 \delaydata_reg[5]  ( .D(n379), .CLK(CLK), .Q(delaydata[5]) );
  DFFPOSX1 \delaydata_reg[6]  ( .D(n375), .CLK(CLK), .Q(delaydata[6]) );
  DFFPOSX1 \intj_reg[7]  ( .D(n875), .CLK(CLK), .Q(intj[7]) );
  DFFPOSX1 \intj_reg[0]  ( .D(n882), .CLK(CLK), .Q(intj[0]) );
  DFFPOSX1 \intj_reg[1]  ( .D(n881), .CLK(CLK), .Q(intj[1]) );
  DFFPOSX1 \intj_reg[2]  ( .D(n880), .CLK(CLK), .Q(intj[2]) );
  DFFPOSX1 \intj_reg[3]  ( .D(n879), .CLK(CLK), .Q(intj[3]) );
  DFFPOSX1 \intj_reg[4]  ( .D(n878), .CLK(CLK), .Q(intj[4]) );
  DFFPOSX1 \intj_reg[5]  ( .D(n877), .CLK(CLK), .Q(intj[5]) );
  DFFPOSX1 \intj_reg[6]  ( .D(n876), .CLK(CLK), .Q(intj[6]) );
  DFFPOSX1 \keyi_reg[2]  ( .D(n874), .CLK(CLK), .Q(keyi[2]) );
  DFFPOSX1 \keyi_reg[1]  ( .D(n873), .CLK(CLK), .Q(keyi[1]) );
  DFFPOSX1 \keyi_reg[0]  ( .D(n872), .CLK(CLK), .Q(keyi[0]) );
  DFFPOSX1 \inti_reg[7]  ( .D(n425), .CLK(CLK), .Q(inti[7]) );
  DFFPOSX1 \inti_reg[0]  ( .D(n411), .CLK(CLK), .Q(inti[0]) );
  DFFPOSX1 \inti_reg[1]  ( .D(n413), .CLK(CLK), .Q(inti[1]) );
  DFFPOSX1 \inti_reg[2]  ( .D(n415), .CLK(CLK), .Q(inti[2]) );
  DFFPOSX1 \inti_reg[3]  ( .D(n417), .CLK(CLK), .Q(inti[3]) );
  DFFPOSX1 \inti_reg[4]  ( .D(n419), .CLK(CLK), .Q(inti[4]) );
  DFFPOSX1 \inti_reg[5]  ( .D(n421), .CLK(CLK), .Q(inti[5]) );
  DFFPOSX1 \inti_reg[6]  ( .D(n423), .CLK(CLK), .Q(inti[6]) );
  DFFPOSX1 \PROCESSED_DATA_reg[0]  ( .D(n759), .CLK(CLK), .Q(PROCESSED_DATA[0]) );
  DFFPOSX1 \PROCESSED_DATA_reg[1]  ( .D(n757), .CLK(CLK), .Q(PROCESSED_DATA[1]) );
  DFFPOSX1 \PROCESSED_DATA_reg[2]  ( .D(n755), .CLK(CLK), .Q(PROCESSED_DATA[2]) );
  DFFPOSX1 \PROCESSED_DATA_reg[3]  ( .D(n753), .CLK(CLK), .Q(PROCESSED_DATA[3]) );
  DFFPOSX1 \PROCESSED_DATA_reg[4]  ( .D(n751), .CLK(CLK), .Q(PROCESSED_DATA[4]) );
  DFFPOSX1 \PROCESSED_DATA_reg[5]  ( .D(n749), .CLK(CLK), .Q(PROCESSED_DATA[5]) );
  DFFPOSX1 \PROCESSED_DATA_reg[6]  ( .D(n747), .CLK(CLK), .Q(PROCESSED_DATA[6]) );
  DFFPOSX1 \PROCESSED_DATA_reg[7]  ( .D(n745), .CLK(CLK), .Q(PROCESSED_DATA[7]) );
  DFFPOSX1 \faddr_reg[7]  ( .D(n744), .CLK(CLK), .Q(faddr[7]) );
  DFFPOSX1 \ADDR_reg[7]  ( .D(n743), .CLK(CLK), .Q(ADDR[7]) );
  DFFPOSX1 \faddr_reg[6]  ( .D(n742), .CLK(CLK), .Q(faddr[6]) );
  DFFPOSX1 \ADDR_reg[6]  ( .D(n741), .CLK(CLK), .Q(ADDR[6]) );
  DFFPOSX1 \faddr_reg[5]  ( .D(n740), .CLK(CLK), .Q(faddr[5]) );
  DFFPOSX1 \ADDR_reg[5]  ( .D(n739), .CLK(CLK), .Q(ADDR[5]) );
  DFFPOSX1 \faddr_reg[4]  ( .D(n738), .CLK(CLK), .Q(faddr[4]) );
  DFFPOSX1 \ADDR_reg[4]  ( .D(n737), .CLK(CLK), .Q(ADDR[4]) );
  DFFPOSX1 \faddr_reg[3]  ( .D(n736), .CLK(CLK), .Q(faddr[3]) );
  DFFPOSX1 \ADDR_reg[3]  ( .D(n735), .CLK(CLK), .Q(ADDR[3]) );
  DFFPOSX1 \faddr_reg[2]  ( .D(n734), .CLK(CLK), .Q(faddr[2]) );
  DFFPOSX1 \ADDR_reg[2]  ( .D(n733), .CLK(CLK), .Q(ADDR[2]) );
  DFFPOSX1 \faddr_reg[1]  ( .D(n732), .CLK(CLK), .Q(faddr[1]) );
  DFFPOSX1 \ADDR_reg[1]  ( .D(n731), .CLK(CLK), .Q(ADDR[1]) );
  DFFPOSX1 \faddr_reg[0]  ( .D(n730), .CLK(CLK), .Q(faddr[0]) );
  DFFPOSX1 \ADDR_reg[0]  ( .D(n729), .CLK(CLK), .Q(ADDR[0]) );
  DFFPOSX1 \fdata_reg[7]  ( .D(n728), .CLK(CLK), .Q(fdata[7]) );
  DFFPOSX1 \fdata_reg[6]  ( .D(n727), .CLK(CLK), .Q(fdata[6]) );
  DFFPOSX1 \fdata_reg[5]  ( .D(n726), .CLK(CLK), .Q(fdata[5]) );
  DFFPOSX1 \fdata_reg[4]  ( .D(n725), .CLK(CLK), .Q(fdata[4]) );
  DFFPOSX1 \fdata_reg[3]  ( .D(n724), .CLK(CLK), .Q(fdata[3]) );
  DFFPOSX1 \fdata_reg[2]  ( .D(n723), .CLK(CLK), .Q(fdata[2]) );
  DFFPOSX1 \fdata_reg[1]  ( .D(n722), .CLK(CLK), .Q(fdata[1]) );
  DFFPOSX1 \fdata_reg[0]  ( .D(n721), .CLK(CLK), .Q(fdata[0]) );
  DFFPOSX1 fw_enable_reg ( .D(n720), .CLK(CLK), .Q(fw_enable) );
  DFFPOSX1 fr_enable_reg ( .D(n719), .CLK(CLK), .Q(fr_enable) );
  DFFPOSX1 W_ENABLE_reg ( .D(n718), .CLK(CLK), .Q(W_ENABLE) );
  DFFPOSX1 R_ENABLE_reg ( .D(n717), .CLK(CLK), .Q(R_ENABLE) );
  DFFPOSX1 \DATA_reg[7]  ( .D(n716), .CLK(CLK), .Q(DATA[7]) );
  DFFPOSX1 \DATA_reg[6]  ( .D(n715), .CLK(CLK), .Q(DATA[6]) );
  DFFPOSX1 \DATA_reg[5]  ( .D(n714), .CLK(CLK), .Q(DATA[5]) );
  DFFPOSX1 \DATA_reg[4]  ( .D(n713), .CLK(CLK), .Q(DATA[4]) );
  DFFPOSX1 \DATA_reg[3]  ( .D(n712), .CLK(CLK), .Q(DATA[3]) );
  DFFPOSX1 \DATA_reg[2]  ( .D(n711), .CLK(CLK), .Q(DATA[2]) );
  DFFPOSX1 \DATA_reg[1]  ( .D(n710), .CLK(CLK), .Q(DATA[1]) );
  DFFPOSX1 \DATA_reg[0]  ( .D(n709), .CLK(CLK), .Q(DATA[0]) );
  NOR2X1 U3 ( .A(n11), .B(n553), .Y(n691) );
  AOI22X1 U7 ( .A(n246), .B(extratemp[7]), .C(n572), .D(temp[7]), .Y(n13) );
  OAI21X1 U8 ( .A(n451), .B(n968), .C(n18), .Y(n11) );
  AOI22X1 U9 ( .A(DATA_IN[7]), .B(n244), .C(prefillCounter[7]), .D(n247), .Y(
        n18) );
  NOR2X1 U10 ( .A(n21), .B(n551), .Y(n693) );
  AOI22X1 U12 ( .A(n246), .B(extratemp[6]), .C(n572), .D(temp[6]), .Y(n23) );
  OAI21X1 U13 ( .A(n451), .B(n969), .C(n25), .Y(n21) );
  AOI22X1 U14 ( .A(DATA_IN[6]), .B(n244), .C(prefillCounter[6]), .D(n247), .Y(
        n25) );
  NOR2X1 U15 ( .A(n26), .B(n549), .Y(n694) );
  AOI22X1 U17 ( .A(n246), .B(extratemp[5]), .C(n572), .D(temp[5]), .Y(n28) );
  OAI21X1 U18 ( .A(n451), .B(n970), .C(n30), .Y(n26) );
  AOI22X1 U19 ( .A(DATA_IN[5]), .B(n244), .C(prefillCounter[5]), .D(n247), .Y(
        n30) );
  NOR2X1 U20 ( .A(n31), .B(n547), .Y(n695) );
  AOI22X1 U22 ( .A(n246), .B(extratemp[4]), .C(n572), .D(temp[4]), .Y(n33) );
  OAI21X1 U23 ( .A(n451), .B(n971), .C(n35), .Y(n31) );
  AOI22X1 U24 ( .A(DATA_IN[4]), .B(n244), .C(prefillCounter[4]), .D(n247), .Y(
        n35) );
  NOR2X1 U25 ( .A(n36), .B(n545), .Y(n696) );
  AOI22X1 U27 ( .A(n246), .B(extratemp[3]), .C(n572), .D(temp[3]), .Y(n38) );
  OAI21X1 U28 ( .A(n451), .B(n972), .C(n40), .Y(n36) );
  AOI22X1 U29 ( .A(DATA_IN[3]), .B(n244), .C(prefillCounter[3]), .D(n247), .Y(
        n40) );
  NOR2X1 U30 ( .A(n41), .B(n543), .Y(n697) );
  AOI22X1 U32 ( .A(n246), .B(extratemp[2]), .C(n572), .D(temp[2]), .Y(n43) );
  OAI21X1 U33 ( .A(n451), .B(n973), .C(n45), .Y(n41) );
  AOI22X1 U34 ( .A(DATA_IN[2]), .B(n244), .C(prefillCounter[2]), .D(n247), .Y(
        n45) );
  NOR2X1 U35 ( .A(n46), .B(n542), .Y(n698) );
  AOI22X1 U37 ( .A(n246), .B(extratemp[1]), .C(n572), .D(temp[1]), .Y(n48) );
  OAI21X1 U38 ( .A(n451), .B(n974), .C(n50), .Y(n46) );
  AOI22X1 U39 ( .A(DATA_IN[1]), .B(n244), .C(prefillCounter[1]), .D(n247), .Y(
        n50) );
  NOR2X1 U40 ( .A(n51), .B(n541), .Y(n699) );
  AOI22X1 U42 ( .A(n246), .B(extratemp[0]), .C(n572), .D(temp[0]), .Y(n53) );
  OAI21X1 U43 ( .A(n451), .B(n975), .C(n55), .Y(n51) );
  AOI22X1 U44 ( .A(DATA_IN[0]), .B(n244), .C(prefillCounter[0]), .D(n247), .Y(
        n55) );
  NOR2X1 U46 ( .A(n57), .B(n58), .Y(n700) );
  NAND2X1 U47 ( .A(n59), .B(n60), .Y(n58) );
  AOI22X1 U48 ( .A(sj[7]), .B(n61), .C(N448), .D(n252), .Y(n60) );
  AOI22X1 U49 ( .A(intj[7]), .B(n250), .C(N503), .D(n241), .Y(n59) );
  NAND2X1 U50 ( .A(n65), .B(n66), .Y(n57) );
  AOI22X1 U51 ( .A(temp[7]), .B(n240), .C(inti[7]), .D(n68), .Y(n66) );
  AOI22X1 U52 ( .A(prefillCounter[7]), .B(n247), .C(faddr[7]), .D(n261), .Y(
        n65) );
  NOR2X1 U53 ( .A(n70), .B(n71), .Y(n702) );
  NAND2X1 U54 ( .A(n72), .B(n73), .Y(n71) );
  AOI22X1 U55 ( .A(sj[6]), .B(n61), .C(N447), .D(n252), .Y(n73) );
  AOI22X1 U56 ( .A(intj[6]), .B(n250), .C(N502), .D(n241), .Y(n72) );
  NAND2X1 U57 ( .A(n74), .B(n75), .Y(n70) );
  AOI22X1 U58 ( .A(temp[6]), .B(n240), .C(inti[6]), .D(n68), .Y(n75) );
  AOI22X1 U59 ( .A(prefillCounter[6]), .B(n247), .C(faddr[6]), .D(n261), .Y(
        n74) );
  NOR2X1 U60 ( .A(n76), .B(n77), .Y(n703) );
  NAND2X1 U61 ( .A(n78), .B(n79), .Y(n77) );
  AOI22X1 U62 ( .A(sj[5]), .B(n61), .C(N446), .D(n252), .Y(n79) );
  AOI22X1 U63 ( .A(intj[5]), .B(n250), .C(N501), .D(n241), .Y(n78) );
  NAND2X1 U64 ( .A(n80), .B(n81), .Y(n76) );
  AOI22X1 U65 ( .A(temp[5]), .B(n240), .C(inti[5]), .D(n68), .Y(n81) );
  AOI22X1 U66 ( .A(prefillCounter[5]), .B(n247), .C(faddr[5]), .D(n261), .Y(
        n80) );
  NOR2X1 U67 ( .A(n82), .B(n83), .Y(n704) );
  NAND2X1 U68 ( .A(n84), .B(n85), .Y(n83) );
  AOI22X1 U69 ( .A(sj[4]), .B(n61), .C(N445), .D(n252), .Y(n85) );
  AOI22X1 U70 ( .A(intj[4]), .B(n250), .C(N500), .D(n241), .Y(n84) );
  NAND2X1 U71 ( .A(n86), .B(n87), .Y(n82) );
  AOI22X1 U72 ( .A(temp[4]), .B(n240), .C(inti[4]), .D(n68), .Y(n87) );
  AOI22X1 U73 ( .A(prefillCounter[4]), .B(n247), .C(faddr[4]), .D(n261), .Y(
        n86) );
  NOR2X1 U74 ( .A(n88), .B(n89), .Y(n705) );
  NAND2X1 U75 ( .A(n90), .B(n91), .Y(n89) );
  AOI22X1 U76 ( .A(sj[3]), .B(n61), .C(N444), .D(n252), .Y(n91) );
  AOI22X1 U77 ( .A(intj[3]), .B(n250), .C(N499), .D(n241), .Y(n90) );
  NAND2X1 U78 ( .A(n92), .B(n93), .Y(n88) );
  AOI22X1 U79 ( .A(temp[3]), .B(n240), .C(inti[3]), .D(n68), .Y(n93) );
  AOI22X1 U80 ( .A(prefillCounter[3]), .B(n247), .C(faddr[3]), .D(n261), .Y(
        n92) );
  NOR2X1 U81 ( .A(n94), .B(n95), .Y(n706) );
  NAND2X1 U82 ( .A(n96), .B(n97), .Y(n95) );
  AOI22X1 U83 ( .A(sj[2]), .B(n61), .C(N443), .D(n252), .Y(n97) );
  AOI22X1 U84 ( .A(intj[2]), .B(n250), .C(N498), .D(n241), .Y(n96) );
  NAND2X1 U85 ( .A(n98), .B(n99), .Y(n94) );
  AOI22X1 U86 ( .A(temp[2]), .B(n240), .C(inti[2]), .D(n68), .Y(n99) );
  AOI22X1 U87 ( .A(prefillCounter[2]), .B(n247), .C(faddr[2]), .D(n261), .Y(
        n98) );
  NOR2X1 U88 ( .A(n100), .B(n101), .Y(n707) );
  NAND2X1 U89 ( .A(n102), .B(n103), .Y(n101) );
  AOI22X1 U90 ( .A(sj[1]), .B(n61), .C(N442), .D(n252), .Y(n103) );
  AOI22X1 U91 ( .A(intj[1]), .B(n250), .C(N497), .D(n241), .Y(n102) );
  NAND2X1 U92 ( .A(n104), .B(n105), .Y(n100) );
  AOI22X1 U93 ( .A(temp[1]), .B(n240), .C(inti[1]), .D(n68), .Y(n105) );
  AOI22X1 U94 ( .A(prefillCounter[1]), .B(n247), .C(faddr[1]), .D(n261), .Y(
        n104) );
  NOR2X1 U95 ( .A(n106), .B(n107), .Y(n708) );
  NAND2X1 U96 ( .A(n108), .B(n109), .Y(n107) );
  AOI22X1 U97 ( .A(sj[0]), .B(n61), .C(n924), .D(n252), .Y(n109) );
  OAI21X1 U98 ( .A(n110), .B(n111), .C(n112), .Y(n61) );
  AOI22X1 U99 ( .A(intj[0]), .B(n250), .C(N496), .D(n241), .Y(n108) );
  NAND2X1 U100 ( .A(n113), .B(n114), .Y(n106) );
  AOI22X1 U101 ( .A(temp[0]), .B(n240), .C(inti[0]), .D(n68), .Y(n114) );
  OAI21X1 U102 ( .A(n115), .B(n116), .C(n503), .Y(n68) );
  AOI22X1 U104 ( .A(prefillCounter[0]), .B(n247), .C(faddr[0]), .D(n261), .Y(
        n113) );
  OAI21X1 U106 ( .A(n218), .B(n188), .C(n249), .Y(n120) );
  OAI21X1 U108 ( .A(n123), .B(n124), .C(n125), .Y(n119) );
  AOI21X1 U109 ( .A(n126), .B(n127), .C(n540), .Y(n125) );
  NOR2X1 U110 ( .A(KEY_ERROR), .B(n128), .Y(n126) );
  OAI21X1 U111 ( .A(n361), .B(n130), .C(n359), .Y(n124) );
  NAND3X1 U112 ( .A(n132), .B(n133), .C(n134), .Y(nextState[3]) );
  AOI21X1 U113 ( .A(n571), .B(n606), .C(n137), .Y(n134) );
  NAND2X1 U114 ( .A(n138), .B(n139), .Y(n137) );
  AOI22X1 U115 ( .A(n140), .B(n359), .C(n522), .D(n142), .Y(n132) );
  NAND3X1 U116 ( .A(n143), .B(n144), .C(n145), .Y(nextState[2]) );
  NOR2X1 U117 ( .A(n146), .B(n147), .Y(n145) );
  OAI21X1 U118 ( .A(n148), .B(n110), .C(n133), .Y(n147) );
  AOI21X1 U119 ( .A(n149), .B(permuteComplete), .C(n150), .Y(n133) );
  NAND2X1 U120 ( .A(n507), .B(n152), .Y(n150) );
  OAI22X1 U121 ( .A(n116), .B(n153), .C(KEY_ERROR), .D(n154), .Y(n146) );
  AOI22X1 U122 ( .A(n155), .B(n156), .C(n157), .D(n158), .Y(n154) );
  NOR2X1 U123 ( .A(n159), .B(n361), .Y(n155) );
  NOR2X1 U124 ( .A(n246), .B(n600), .Y(n144) );
  NOR2X1 U125 ( .A(n594), .B(n162), .Y(n143) );
  NAND3X1 U126 ( .A(n163), .B(n164), .C(n165), .Y(nextState[1]) );
  NOR2X1 U127 ( .A(n166), .B(n167), .Y(n165) );
  OAI21X1 U128 ( .A(n168), .B(n169), .C(n170), .Y(n167) );
  NAND3X1 U129 ( .A(n171), .B(n401), .C(n173), .Y(n169) );
  NOR2X1 U130 ( .A(prefillCounter[2]), .B(prefillCounter[1]), .Y(n173) );
  NAND3X1 U131 ( .A(n174), .B(n889), .C(n176), .Y(n168) );
  NOR2X1 U132 ( .A(prefillCounter[4]), .B(prefillCounter[3]), .Y(n176) );
  NOR2X1 U133 ( .A(prefillCounter[7]), .B(prefillCounter[6]), .Y(n174) );
  AOI22X1 U135 ( .A(n178), .B(state[0]), .C(n179), .D(n359), .Y(n163) );
  OAI21X1 U137 ( .A(n518), .B(n158), .C(n181), .Y(n179) );
  NAND2X1 U138 ( .A(n142), .B(n182), .Y(n181) );
  OAI21X1 U139 ( .A(n183), .B(n158), .C(n184), .Y(n182) );
  OAI21X1 U140 ( .A(n159), .B(n361), .C(n569), .Y(n184) );
  NAND3X1 U143 ( .A(n367), .B(n365), .C(BYTE_READY), .Y(n158) );
  NOR2X1 U145 ( .A(state[1]), .B(n116), .Y(n178) );
  NAND3X1 U146 ( .A(n189), .B(n190), .C(n191), .Y(nextState[0]) );
  NOR2X1 U147 ( .A(n252), .B(n192), .Y(n191) );
  OAI21X1 U148 ( .A(KEY_ERROR), .B(n193), .C(n164), .Y(n192) );
  NOR2X1 U149 ( .A(n194), .B(n195), .Y(n164) );
  OAI21X1 U150 ( .A(permuteComplete), .B(n562), .C(n197), .Y(n195) );
  NAND3X1 U151 ( .A(n152), .B(n198), .C(n199), .Y(n194) );
  AOI21X1 U152 ( .A(n156), .B(n128), .C(n200), .Y(n193) );
  OAI21X1 U153 ( .A(n218), .B(n201), .C(n202), .Y(n200) );
  NAND3X1 U154 ( .A(BYTE_READY), .B(n157), .C(n363), .Y(n202) );
  NAND2X1 U156 ( .A(OPCODE[0]), .B(n365), .Y(n130) );
  NAND2X1 U158 ( .A(BYTE_READY), .B(n204), .Y(n128) );
  OAI21X1 U159 ( .A(OPCODE[0]), .B(OPCODE[1]), .C(n186), .Y(n204) );
  NAND2X1 U160 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n186) );
  NOR2X1 U161 ( .A(n540), .B(n246), .Y(n190) );
  NOR2X1 U162 ( .A(n171), .B(n205), .Y(n189) );
  OAI21X1 U163 ( .A(n300), .B(n403), .C(n207), .Y(n709) );
  NAND2X1 U164 ( .A(DATA[0]), .B(n290), .Y(n207) );
  OAI21X1 U165 ( .A(n302), .B(n449), .C(n209), .Y(n710) );
  NAND2X1 U166 ( .A(DATA[1]), .B(n305), .Y(n209) );
  OAI21X1 U167 ( .A(n302), .B(n447), .C(n211), .Y(n711) );
  NAND2X1 U168 ( .A(DATA[2]), .B(n305), .Y(n211) );
  OAI21X1 U169 ( .A(n302), .B(n445), .C(n213), .Y(n712) );
  NAND2X1 U170 ( .A(DATA[3]), .B(n305), .Y(n213) );
  OAI21X1 U171 ( .A(n302), .B(n443), .C(n215), .Y(n713) );
  NAND2X1 U172 ( .A(DATA[4]), .B(RST), .Y(n215) );
  OAI21X1 U173 ( .A(n302), .B(n441), .C(n217), .Y(n714) );
  NAND2X1 U174 ( .A(DATA[5]), .B(n305), .Y(n217) );
  OAI21X1 U175 ( .A(n302), .B(n439), .C(n219), .Y(n715) );
  NAND2X1 U176 ( .A(DATA[6]), .B(n305), .Y(n219) );
  OAI21X1 U177 ( .A(n302), .B(n437), .C(n221), .Y(n716) );
  NAND2X1 U178 ( .A(DATA[7]), .B(n305), .Y(n221) );
  OAI21X1 U179 ( .A(n302), .B(n222), .C(n223), .Y(n717) );
  NAND2X1 U180 ( .A(R_ENABLE), .B(n305), .Y(n223) );
  AOI21X1 U181 ( .A(fr_enable), .B(n224), .C(n225), .Y(n222) );
  OAI21X1 U182 ( .A(n300), .B(n226), .C(n227), .Y(n718) );
  NAND2X1 U183 ( .A(W_ENABLE), .B(n302), .Y(n227) );
  AOI21X1 U184 ( .A(fw_enable), .B(n185), .C(n229), .Y(n226) );
  OAI21X1 U185 ( .A(n300), .B(n504), .C(n231), .Y(n719) );
  OAI21X1 U186 ( .A(n300), .B(n224), .C(fr_enable), .Y(n231) );
  NAND3X1 U187 ( .A(n3), .B(n233), .C(n234), .Y(n224) );
  NOR2X1 U188 ( .A(n577), .B(n236), .Y(n234) );
  NAND2X1 U189 ( .A(n210), .B(n10), .Y(n236) );
  NAND2X1 U191 ( .A(n579), .B(n604), .Y(n112) );
  OAI21X1 U192 ( .A(n300), .B(n514), .C(n242), .Y(n720) );
  OAI21X1 U193 ( .A(n300), .B(n185), .C(fw_enable), .Y(n242) );
  NAND3X1 U195 ( .A(n210), .B(n10), .C(n243), .Y(n229) );
  NOR2X1 U196 ( .A(n244), .B(n572), .Y(n243) );
  OAI22X1 U197 ( .A(n331), .B(n975), .C(n297), .D(n403), .Y(n721) );
  OAI22X1 U200 ( .A(n331), .B(n974), .C(n295), .D(n449), .Y(n722) );
  OAI22X1 U203 ( .A(n331), .B(n973), .C(n297), .D(n447), .Y(n723) );
  OAI22X1 U206 ( .A(n331), .B(n972), .C(n295), .D(n445), .Y(n724) );
  OAI22X1 U209 ( .A(n333), .B(n971), .C(n297), .D(n443), .Y(n725) );
  OAI22X1 U212 ( .A(n329), .B(n970), .C(n295), .D(n441), .Y(n726) );
  OAI22X1 U215 ( .A(n329), .B(n969), .C(n297), .D(n439), .Y(n727) );
  OAI22X1 U218 ( .A(n329), .B(n968), .C(n295), .D(n437), .Y(n728) );
  OAI21X1 U221 ( .A(n300), .B(n405), .C(n245), .Y(n729) );
  NAND2X1 U222 ( .A(ADDR[0]), .B(n302), .Y(n245) );
  OAI22X1 U223 ( .A(n326), .B(n967), .C(n295), .D(n405), .Y(n730) );
  OAI21X1 U226 ( .A(n300), .B(n471), .C(n248), .Y(n731) );
  NAND2X1 U227 ( .A(ADDR[1]), .B(n305), .Y(n248) );
  OAI22X1 U228 ( .A(n335), .B(n966), .C(n295), .D(n471), .Y(n732) );
  OAI21X1 U231 ( .A(n300), .B(n473), .C(n251), .Y(n733) );
  NAND2X1 U232 ( .A(ADDR[2]), .B(n302), .Y(n251) );
  OAI22X1 U233 ( .A(n337), .B(n965), .C(n295), .D(n473), .Y(n734) );
  OAI21X1 U236 ( .A(n300), .B(n475), .C(n254), .Y(n735) );
  NAND2X1 U237 ( .A(ADDR[3]), .B(n305), .Y(n254) );
  OAI22X1 U238 ( .A(n327), .B(n964), .C(n295), .D(n475), .Y(n736) );
  OAI21X1 U241 ( .A(n300), .B(n480), .C(n257), .Y(n737) );
  NAND2X1 U242 ( .A(ADDR[4]), .B(n305), .Y(n257) );
  OAI22X1 U243 ( .A(n307), .B(n963), .C(n295), .D(n480), .Y(n738) );
  OAI21X1 U246 ( .A(n300), .B(n482), .C(n260), .Y(n739) );
  NAND2X1 U247 ( .A(ADDR[5]), .B(n305), .Y(n260) );
  OAI22X1 U248 ( .A(n318), .B(n962), .C(n295), .D(n482), .Y(n740) );
  OAI21X1 U251 ( .A(n297), .B(n488), .C(n263), .Y(n741) );
  NAND2X1 U252 ( .A(ADDR[6]), .B(n305), .Y(n263) );
  OAI22X1 U253 ( .A(n317), .B(n961), .C(n295), .D(n488), .Y(n742) );
  OAI21X1 U256 ( .A(n297), .B(n498), .C(n266), .Y(n743) );
  NAND2X1 U257 ( .A(ADDR[7]), .B(n305), .Y(n266) );
  OAI22X1 U258 ( .A(n311), .B(n960), .C(n295), .D(n498), .Y(n744) );
  OAI21X1 U261 ( .A(n297), .B(n369), .C(n269), .Y(n745) );
  NAND2X1 U262 ( .A(PROCESSED_DATA[7]), .B(n305), .Y(n269) );
  OAI21X1 U264 ( .A(n500), .B(n959), .C(n272), .Y(nextProcessedData[7]) );
  AOI22X1 U265 ( .A(n273), .B(n274), .C(BYTE[7]), .D(n575), .Y(n272) );
  XOR2X1 U266 ( .A(temp[7]), .B(delaydata[7]), .Y(n274) );
  OAI21X1 U268 ( .A(n297), .B(n373), .C(n276), .Y(n747) );
  NAND2X1 U269 ( .A(PROCESSED_DATA[6]), .B(n305), .Y(n276) );
  OAI21X1 U271 ( .A(n500), .B(n958), .C(n278), .Y(nextProcessedData[6]) );
  AOI22X1 U272 ( .A(n273), .B(n279), .C(BYTE[6]), .D(n575), .Y(n278) );
  XOR2X1 U273 ( .A(temp[6]), .B(delaydata[6]), .Y(n279) );
  OAI21X1 U275 ( .A(n297), .B(n377), .C(n281), .Y(n749) );
  NAND2X1 U276 ( .A(PROCESSED_DATA[5]), .B(n305), .Y(n281) );
  OAI21X1 U278 ( .A(n500), .B(n957), .C(n283), .Y(nextProcessedData[5]) );
  AOI22X1 U279 ( .A(n273), .B(n284), .C(BYTE[5]), .D(n575), .Y(n283) );
  XOR2X1 U280 ( .A(temp[5]), .B(delaydata[5]), .Y(n284) );
  OAI21X1 U282 ( .A(n297), .B(n381), .C(n286), .Y(n751) );
  NAND2X1 U283 ( .A(PROCESSED_DATA[4]), .B(n305), .Y(n286) );
  OAI21X1 U285 ( .A(n500), .B(n956), .C(n288), .Y(nextProcessedData[4]) );
  AOI22X1 U286 ( .A(n273), .B(n289), .C(BYTE[4]), .D(n575), .Y(n288) );
  XOR2X1 U287 ( .A(temp[4]), .B(delaydata[4]), .Y(n289) );
  OAI21X1 U289 ( .A(n300), .B(n385), .C(n291), .Y(n753) );
  NAND2X1 U290 ( .A(PROCESSED_DATA[3]), .B(n305), .Y(n291) );
  OAI21X1 U292 ( .A(n500), .B(n955), .C(n293), .Y(nextProcessedData[3]) );
  AOI22X1 U293 ( .A(n273), .B(n294), .C(BYTE[3]), .D(n575), .Y(n293) );
  XOR2X1 U294 ( .A(temp[3]), .B(delaydata[3]), .Y(n294) );
  OAI21X1 U296 ( .A(n297), .B(n389), .C(n296), .Y(n755) );
  NAND2X1 U297 ( .A(PROCESSED_DATA[2]), .B(n305), .Y(n296) );
  OAI21X1 U299 ( .A(n500), .B(n954), .C(n298), .Y(nextProcessedData[2]) );
  AOI22X1 U300 ( .A(n273), .B(n299), .C(BYTE[2]), .D(n575), .Y(n298) );
  XOR2X1 U301 ( .A(temp[2]), .B(delaydata[2]), .Y(n299) );
  OAI21X1 U303 ( .A(n297), .B(n393), .C(n301), .Y(n757) );
  NAND2X1 U304 ( .A(PROCESSED_DATA[1]), .B(RST), .Y(n301) );
  OAI21X1 U306 ( .A(n500), .B(n953), .C(n303), .Y(nextProcessedData[1]) );
  AOI22X1 U307 ( .A(n273), .B(n304), .C(BYTE[1]), .D(n575), .Y(n303) );
  XOR2X1 U308 ( .A(temp[1]), .B(delaydata[1]), .Y(n304) );
  OAI21X1 U310 ( .A(n297), .B(n397), .C(n306), .Y(n759) );
  NAND2X1 U311 ( .A(PROCESSED_DATA[0]), .B(RST), .Y(n306) );
  OAI21X1 U313 ( .A(n500), .B(n952), .C(n308), .Y(nextProcessedData[0]) );
  AOI22X1 U314 ( .A(n273), .B(n309), .C(BYTE[0]), .D(n575), .Y(n308) );
  XOR2X1 U315 ( .A(temp[0]), .B(delaydata[0]), .Y(n309) );
  NAND3X1 U318 ( .A(n253), .B(n505), .C(n312), .Y(n310) );
  NOR2X1 U319 ( .A(n313), .B(n314), .Y(n312) );
  AOI22X1 U322 ( .A(BYTE[7]), .B(n6), .C(n262), .D(delaydata[7]), .Y(n316) );
  AOI22X1 U324 ( .A(BYTE[0]), .B(n6), .C(n262), .D(delaydata[0]), .Y(n319) );
  AOI22X1 U326 ( .A(BYTE[1]), .B(n6), .C(n262), .D(delaydata[1]), .Y(n320) );
  AOI22X1 U328 ( .A(BYTE[2]), .B(n6), .C(n262), .D(delaydata[2]), .Y(n321) );
  AOI22X1 U330 ( .A(BYTE[3]), .B(n6), .C(n262), .D(delaydata[3]), .Y(n322) );
  AOI22X1 U332 ( .A(BYTE[4]), .B(n6), .C(n262), .D(delaydata[4]), .Y(n323) );
  AOI22X1 U334 ( .A(BYTE[5]), .B(n6), .C(n262), .D(delaydata[5]), .Y(n324) );
  AOI22X1 U336 ( .A(BYTE[6]), .B(n6), .C(n262), .D(delaydata[6]), .Y(n325) );
  OAI21X1 U339 ( .A(n271), .B(n616), .C(n330), .Y(n792) );
  NAND2X1 U340 ( .A(KEY[56]), .B(n287), .Y(n330) );
  OAI21X1 U342 ( .A(n268), .B(n618), .C(n332), .Y(n793) );
  NAND2X1 U343 ( .A(KEY[57]), .B(n287), .Y(n332) );
  OAI21X1 U345 ( .A(n268), .B(n624), .C(n334), .Y(n794) );
  NAND2X1 U346 ( .A(KEY[58]), .B(n287), .Y(n334) );
  OAI21X1 U348 ( .A(n268), .B(n626), .C(n336), .Y(n795) );
  NAND2X1 U349 ( .A(KEY[59]), .B(n287), .Y(n336) );
  OAI21X1 U351 ( .A(n268), .B(n629), .C(n338), .Y(n796) );
  NAND2X1 U352 ( .A(KEY[60]), .B(n287), .Y(n338) );
  OAI21X1 U354 ( .A(n268), .B(n630), .C(n340), .Y(n797) );
  NAND2X1 U355 ( .A(KEY[61]), .B(n285), .Y(n340) );
  OAI21X1 U357 ( .A(n268), .B(n632), .C(n342), .Y(n798) );
  NAND2X1 U358 ( .A(KEY[62]), .B(n285), .Y(n342) );
  OAI21X1 U360 ( .A(n268), .B(n636), .C(n344), .Y(n799) );
  NAND2X1 U361 ( .A(KEY[63]), .B(n285), .Y(n344) );
  OAI21X1 U363 ( .A(n268), .B(n637), .C(n346), .Y(n800) );
  NAND2X1 U364 ( .A(KEY[48]), .B(n285), .Y(n346) );
  OAI21X1 U366 ( .A(n268), .B(n638), .C(n348), .Y(n801) );
  NAND2X1 U367 ( .A(KEY[49]), .B(n285), .Y(n348) );
  OAI21X1 U369 ( .A(n268), .B(n648), .C(n350), .Y(n802) );
  NAND2X1 U370 ( .A(KEY[50]), .B(n285), .Y(n350) );
  OAI21X1 U372 ( .A(n268), .B(n649), .C(n352), .Y(n803) );
  NAND2X1 U373 ( .A(KEY[51]), .B(n285), .Y(n352) );
  OAI21X1 U375 ( .A(n268), .B(n650), .C(n354), .Y(n804) );
  NAND2X1 U376 ( .A(KEY[52]), .B(n285), .Y(n354) );
  OAI21X1 U378 ( .A(n268), .B(n651), .C(n356), .Y(n805) );
  NAND2X1 U379 ( .A(KEY[53]), .B(n285), .Y(n356) );
  OAI21X1 U381 ( .A(n270), .B(n692), .C(n358), .Y(n806) );
  NAND2X1 U382 ( .A(KEY[54]), .B(n285), .Y(n358) );
  OAI21X1 U384 ( .A(n270), .B(n701), .C(n360), .Y(n807) );
  NAND2X1 U385 ( .A(KEY[55]), .B(n282), .Y(n360) );
  OAI21X1 U387 ( .A(n270), .B(n746), .C(n362), .Y(n808) );
  NAND2X1 U388 ( .A(KEY[40]), .B(n285), .Y(n362) );
  OAI21X1 U390 ( .A(n270), .B(n748), .C(n364), .Y(n809) );
  NAND2X1 U391 ( .A(KEY[41]), .B(n285), .Y(n364) );
  OAI21X1 U393 ( .A(n270), .B(n750), .C(n366), .Y(n810) );
  NAND2X1 U394 ( .A(KEY[42]), .B(n282), .Y(n366) );
  OAI21X1 U396 ( .A(n270), .B(n752), .C(n368), .Y(n811) );
  NAND2X1 U397 ( .A(KEY[43]), .B(n285), .Y(n368) );
  OAI21X1 U399 ( .A(n270), .B(n754), .C(n370), .Y(n812) );
  NAND2X1 U400 ( .A(KEY[44]), .B(n282), .Y(n370) );
  OAI21X1 U402 ( .A(n270), .B(n756), .C(n372), .Y(n813) );
  NAND2X1 U403 ( .A(KEY[45]), .B(n282), .Y(n372) );
  OAI21X1 U405 ( .A(n270), .B(n758), .C(n374), .Y(n814) );
  NAND2X1 U406 ( .A(KEY[46]), .B(n282), .Y(n374) );
  OAI21X1 U408 ( .A(n270), .B(n760), .C(n376), .Y(n815) );
  NAND2X1 U409 ( .A(KEY[47]), .B(n282), .Y(n376) );
  OAI21X1 U411 ( .A(n270), .B(n761), .C(n378), .Y(n816) );
  NAND2X1 U412 ( .A(KEY[32]), .B(n282), .Y(n378) );
  OAI21X1 U414 ( .A(n270), .B(n762), .C(n380), .Y(n817) );
  NAND2X1 U415 ( .A(KEY[33]), .B(n282), .Y(n380) );
  OAI21X1 U417 ( .A(n270), .B(n763), .C(n382), .Y(n818) );
  NAND2X1 U418 ( .A(KEY[34]), .B(n280), .Y(n382) );
  OAI21X1 U420 ( .A(n271), .B(n764), .C(n384), .Y(n819) );
  NAND2X1 U421 ( .A(KEY[35]), .B(n280), .Y(n384) );
  OAI21X1 U423 ( .A(n271), .B(n765), .C(n386), .Y(n820) );
  NAND2X1 U424 ( .A(KEY[36]), .B(n282), .Y(n386) );
  OAI21X1 U426 ( .A(n271), .B(n766), .C(n388), .Y(n821) );
  NAND2X1 U427 ( .A(KEY[37]), .B(n280), .Y(n388) );
  OAI21X1 U429 ( .A(n271), .B(n767), .C(n390), .Y(n822) );
  NAND2X1 U430 ( .A(KEY[38]), .B(n280), .Y(n390) );
  OAI21X1 U432 ( .A(n271), .B(n768), .C(n392), .Y(n823) );
  NAND2X1 U433 ( .A(KEY[39]), .B(n282), .Y(n392) );
  OAI21X1 U435 ( .A(n275), .B(n769), .C(n394), .Y(n824) );
  NAND2X1 U436 ( .A(KEY[24]), .B(n280), .Y(n394) );
  OAI21X1 U437 ( .A(n271), .B(n770), .C(n396), .Y(n825) );
  NAND2X1 U438 ( .A(KEY[25]), .B(n280), .Y(n396) );
  OAI21X1 U439 ( .A(n271), .B(n771), .C(n398), .Y(n826) );
  NAND2X1 U440 ( .A(KEY[26]), .B(n280), .Y(n398) );
  OAI21X1 U441 ( .A(n271), .B(n772), .C(n400), .Y(n827) );
  NAND2X1 U442 ( .A(KEY[27]), .B(n280), .Y(n400) );
  OAI21X1 U443 ( .A(n271), .B(n773), .C(n402), .Y(n828) );
  NAND2X1 U444 ( .A(KEY[28]), .B(n280), .Y(n402) );
  OAI21X1 U445 ( .A(n271), .B(n774), .C(n404), .Y(n829) );
  NAND2X1 U446 ( .A(KEY[29]), .B(n280), .Y(n404) );
  OAI21X1 U447 ( .A(n271), .B(n775), .C(n406), .Y(n830) );
  NAND2X1 U448 ( .A(KEY[30]), .B(n280), .Y(n406) );
  OAI21X1 U449 ( .A(n271), .B(n776), .C(n408), .Y(n831) );
  NAND2X1 U450 ( .A(KEY[31]), .B(n280), .Y(n408) );
  OAI21X1 U451 ( .A(n275), .B(n777), .C(n410), .Y(n832) );
  NAND2X1 U452 ( .A(KEY[16]), .B(n280), .Y(n410) );
  OAI21X1 U453 ( .A(n275), .B(n778), .C(n412), .Y(n833) );
  NAND2X1 U454 ( .A(KEY[17]), .B(n277), .Y(n412) );
  OAI21X1 U455 ( .A(n275), .B(n779), .C(n414), .Y(n834) );
  NAND2X1 U456 ( .A(KEY[18]), .B(n280), .Y(n414) );
  OAI21X1 U457 ( .A(n275), .B(n780), .C(n416), .Y(n835) );
  NAND2X1 U458 ( .A(KEY[19]), .B(n280), .Y(n416) );
  OAI21X1 U459 ( .A(n275), .B(n781), .C(n418), .Y(n836) );
  NAND2X1 U460 ( .A(KEY[20]), .B(n282), .Y(n418) );
  OAI21X1 U461 ( .A(n275), .B(n782), .C(n420), .Y(n837) );
  NAND2X1 U462 ( .A(KEY[21]), .B(n280), .Y(n420) );
  OAI21X1 U463 ( .A(n275), .B(n783), .C(n422), .Y(n838) );
  NAND2X1 U464 ( .A(KEY[22]), .B(n282), .Y(n422) );
  OAI21X1 U465 ( .A(n275), .B(n784), .C(n424), .Y(n839) );
  NAND2X1 U466 ( .A(KEY[23]), .B(n280), .Y(n424) );
  OAI21X1 U467 ( .A(n277), .B(n785), .C(n426), .Y(n840) );
  NAND2X1 U468 ( .A(KEY[8]), .B(n282), .Y(n426) );
  OAI21X1 U469 ( .A(n277), .B(n786), .C(n428), .Y(n841) );
  NAND2X1 U470 ( .A(KEY[9]), .B(n282), .Y(n428) );
  OAI21X1 U471 ( .A(n275), .B(n787), .C(n430), .Y(n842) );
  NAND2X1 U472 ( .A(KEY[10]), .B(n280), .Y(n430) );
  OAI21X1 U473 ( .A(n277), .B(n788), .C(n432), .Y(n843) );
  NAND2X1 U474 ( .A(KEY[11]), .B(n282), .Y(n432) );
  OAI21X1 U475 ( .A(n277), .B(n789), .C(n434), .Y(n844) );
  NAND2X1 U476 ( .A(KEY[12]), .B(n282), .Y(n434) );
  OAI21X1 U477 ( .A(n275), .B(n790), .C(n436), .Y(n845) );
  NAND2X1 U478 ( .A(KEY[13]), .B(n282), .Y(n436) );
  OAI21X1 U479 ( .A(n275), .B(n791), .C(n438), .Y(n846) );
  NAND2X1 U480 ( .A(KEY[14]), .B(n285), .Y(n438) );
  OAI21X1 U481 ( .A(n277), .B(n864), .C(n440), .Y(n847) );
  NAND2X1 U482 ( .A(KEY[6]), .B(n282), .Y(n440) );
  OAI21X1 U483 ( .A(n275), .B(n865), .C(n442), .Y(n848) );
  NAND2X1 U484 ( .A(KEY[5]), .B(n285), .Y(n442) );
  OAI21X1 U485 ( .A(n277), .B(n866), .C(n444), .Y(n849) );
  NAND2X1 U486 ( .A(KEY[4]), .B(n285), .Y(n444) );
  OAI21X1 U487 ( .A(n277), .B(n867), .C(n446), .Y(n850) );
  NAND2X1 U488 ( .A(KEY[3]), .B(n285), .Y(n446) );
  OAI21X1 U489 ( .A(n277), .B(n868), .C(n448), .Y(n851) );
  NAND2X1 U490 ( .A(KEY[2]), .B(n285), .Y(n448) );
  OAI21X1 U491 ( .A(n277), .B(n869), .C(n450), .Y(n852) );
  NAND2X1 U492 ( .A(KEY[1]), .B(n287), .Y(n450) );
  OAI21X1 U493 ( .A(n277), .B(n870), .C(n452), .Y(n853) );
  NAND2X1 U494 ( .A(KEY[0]), .B(n287), .Y(n452) );
  OAI21X1 U495 ( .A(n277), .B(n871), .C(n454), .Y(n854) );
  NAND2X1 U496 ( .A(KEY[15]), .B(n287), .Y(n454) );
  OAI21X1 U497 ( .A(n277), .B(n883), .C(n456), .Y(n855) );
  NAND2X1 U498 ( .A(KEY[7]), .B(n287), .Y(n456) );
  NOR2X1 U499 ( .A(n457), .B(n313), .Y(n328) );
  OAI21X1 U500 ( .A(n469), .B(n916), .C(n460), .Y(n856) );
  AOI22X1 U501 ( .A(N527), .B(n14), .C(n180), .D(DATA_IN[7]), .Y(n460) );
  OAI21X1 U503 ( .A(n469), .B(n923), .C(n464), .Y(n857) );
  AOI22X1 U504 ( .A(N526), .B(n14), .C(n180), .D(DATA_IN[6]), .Y(n464) );
  OAI21X1 U506 ( .A(n469), .B(n922), .C(n466), .Y(n858) );
  AOI22X1 U507 ( .A(N525), .B(n14), .C(n180), .D(DATA_IN[5]), .Y(n466) );
  OAI21X1 U509 ( .A(n469), .B(n921), .C(n468), .Y(n859) );
  AOI22X1 U510 ( .A(N524), .B(n14), .C(n180), .D(DATA_IN[4]), .Y(n468) );
  OAI21X1 U512 ( .A(n469), .B(n920), .C(n470), .Y(n860) );
  AOI22X1 U513 ( .A(N523), .B(n14), .C(n180), .D(DATA_IN[3]), .Y(n470) );
  OAI21X1 U515 ( .A(n469), .B(n919), .C(n472), .Y(n861) );
  AOI22X1 U516 ( .A(N522), .B(n14), .C(n180), .D(DATA_IN[2]), .Y(n472) );
  OAI21X1 U518 ( .A(n469), .B(n918), .C(n474), .Y(n862) );
  AOI22X1 U519 ( .A(N521), .B(n14), .C(n180), .D(DATA_IN[1]), .Y(n474) );
  OAI21X1 U521 ( .A(n469), .B(n917), .C(n476), .Y(n863) );
  AOI22X1 U522 ( .A(N520), .B(n14), .C(n180), .D(DATA_IN[0]), .Y(n476) );
  NAND3X1 U527 ( .A(n479), .B(n509), .C(n481), .Y(n477) );
  NOR2X1 U528 ( .A(n315), .B(n261), .Y(n481) );
  NAND3X1 U530 ( .A(n483), .B(n210), .C(n484), .Y(n315) );
  NOR2X1 U532 ( .A(n302), .B(n171), .Y(n479) );
  AOI22X1 U534 ( .A(n259), .B(extratemp[0]), .C(DATA_IN[0]), .D(n258), .Y(n486) );
  AOI22X1 U536 ( .A(n259), .B(extratemp[1]), .C(DATA_IN[1]), .D(n258), .Y(n489) );
  AOI22X1 U538 ( .A(n259), .B(extratemp[2]), .C(DATA_IN[2]), .D(n258), .Y(n490) );
  AOI22X1 U540 ( .A(n259), .B(extratemp[3]), .C(DATA_IN[3]), .D(n258), .Y(n491) );
  AOI22X1 U542 ( .A(n259), .B(extratemp[4]), .C(DATA_IN[4]), .D(n258), .Y(n492) );
  AOI22X1 U544 ( .A(n259), .B(extratemp[5]), .C(DATA_IN[5]), .D(n258), .Y(n493) );
  AOI22X1 U546 ( .A(n259), .B(extratemp[6]), .C(DATA_IN[6]), .D(n258), .Y(n494) );
  AOI22X1 U548 ( .A(n259), .B(extratemp[7]), .C(DATA_IN[7]), .D(n258), .Y(n495) );
  NAND3X1 U550 ( .A(n138), .B(n210), .C(n496), .Y(n487) );
  NOR2X1 U551 ( .A(n497), .B(n56), .Y(n496) );
  NAND3X1 U552 ( .A(n5), .B(n520), .C(n3), .Y(n56) );
  NAND2X1 U553 ( .A(n579), .B(n142), .Y(n138) );
  OAI22X1 U555 ( .A(n429), .B(n924), .C(n502), .D(n951), .Y(n872) );
  OAI22X1 U556 ( .A(n429), .B(n357), .C(n502), .D(n228), .Y(n873) );
  OAI22X1 U557 ( .A(n429), .B(n925), .C(n502), .D(n945), .Y(n874) );
  NOR2X1 U559 ( .A(n508), .B(n313), .Y(n502) );
  OAI21X1 U560 ( .A(n409), .B(n930), .C(n510), .Y(n875) );
  NAND2X1 U561 ( .A(N519), .B(n511), .Y(n510) );
  OAI21X1 U563 ( .A(n409), .B(n937), .C(n513), .Y(n876) );
  NAND2X1 U564 ( .A(N518), .B(n511), .Y(n513) );
  OAI21X1 U566 ( .A(n409), .B(n936), .C(n515), .Y(n877) );
  NAND2X1 U567 ( .A(N517), .B(n511), .Y(n515) );
  OAI21X1 U569 ( .A(n409), .B(n935), .C(n517), .Y(n878) );
  NAND2X1 U570 ( .A(N516), .B(n511), .Y(n517) );
  OAI21X1 U572 ( .A(n409), .B(n934), .C(n519), .Y(n879) );
  NAND2X1 U573 ( .A(N515), .B(n511), .Y(n519) );
  OAI21X1 U575 ( .A(n409), .B(n933), .C(n521), .Y(n880) );
  NAND2X1 U576 ( .A(N514), .B(n511), .Y(n521) );
  OAI21X1 U578 ( .A(n409), .B(n932), .C(n523), .Y(n881) );
  NAND2X1 U579 ( .A(N513), .B(n511), .Y(n523) );
  OAI21X1 U581 ( .A(n409), .B(n931), .C(n525), .Y(n882) );
  NAND2X1 U582 ( .A(N512), .B(n511), .Y(n525) );
  NOR2X1 U583 ( .A(n152), .B(n526), .Y(n511) );
  NOR2X1 U587 ( .A(n302), .B(n594), .Y(n529) );
  AOI22X1 U589 ( .A(n256), .B(inti[7]), .C(N503), .D(n216), .Y(n530) );
  AOI22X1 U591 ( .A(n256), .B(inti[6]), .C(N502), .D(n216), .Y(n533) );
  AOI22X1 U593 ( .A(n256), .B(inti[5]), .C(N501), .D(n216), .Y(n534) );
  AOI22X1 U595 ( .A(n256), .B(inti[4]), .C(N500), .D(n216), .Y(n535) );
  AOI22X1 U597 ( .A(n256), .B(inti[3]), .C(N499), .D(n214), .Y(n536) );
  AOI22X1 U599 ( .A(n256), .B(inti[2]), .C(N498), .D(n214), .Y(n537) );
  AOI22X1 U601 ( .A(n256), .B(inti[1]), .C(N497), .D(n214), .Y(n538) );
  AOI22X1 U603 ( .A(n256), .B(inti[0]), .C(N496), .D(n214), .Y(n539) );
  NOR2X1 U604 ( .A(n256), .B(n507), .Y(n532) );
  NAND3X1 U605 ( .A(n557), .B(n520), .C(n431), .Y(n531) );
  OAI21X1 U606 ( .A(n407), .B(n220), .C(n544), .Y(n891) );
  NAND2X1 U607 ( .A(N480), .B(n594), .Y(n544) );
  OAI21X1 U609 ( .A(n407), .B(n944), .C(n546), .Y(n892) );
  NAND2X1 U610 ( .A(N481), .B(n594), .Y(n546) );
  OAI21X1 U612 ( .A(n407), .B(n943), .C(n548), .Y(n893) );
  NAND2X1 U613 ( .A(N482), .B(n594), .Y(n548) );
  OAI21X1 U615 ( .A(n407), .B(n942), .C(n550), .Y(n894) );
  NAND2X1 U616 ( .A(N483), .B(n594), .Y(n550) );
  OAI21X1 U618 ( .A(n407), .B(n941), .C(n552), .Y(n895) );
  NAND2X1 U619 ( .A(N484), .B(n594), .Y(n552) );
  OAI21X1 U621 ( .A(n407), .B(n940), .C(n554), .Y(n896) );
  NAND2X1 U622 ( .A(N485), .B(n594), .Y(n554) );
  OAI21X1 U624 ( .A(n407), .B(n939), .C(n556), .Y(n897) );
  NAND2X1 U625 ( .A(N486), .B(n594), .Y(n556) );
  NAND2X1 U628 ( .A(N487), .B(n594), .Y(n558) );
  NAND3X1 U631 ( .A(n528), .B(n152), .C(n527), .Y(n559) );
  NOR2X1 U632 ( .A(n560), .B(n561), .Y(n527) );
  NAND3X1 U633 ( .A(n3), .B(n557), .C(n435), .Y(n561) );
  NAND3X1 U634 ( .A(n581), .B(n520), .C(n563), .Y(n560) );
  OAI21X1 U637 ( .A(n557), .B(n565), .C(n566), .Y(n899) );
  OAI21X1 U638 ( .A(n567), .B(n508), .C(permuteComplete), .Y(n566) );
  NAND2X1 U639 ( .A(n568), .B(n427), .Y(n565) );
  NAND3X1 U641 ( .A(n172), .B(n507), .C(n431), .Y(n508) );
  NAND3X1 U643 ( .A(n253), .B(n329), .C(n435), .Y(n570) );
  OAI21X1 U646 ( .A(n433), .B(n929), .C(n573), .Y(n900) );
  NAND2X1 U647 ( .A(N431), .B(n574), .Y(n573) );
  OAI21X1 U649 ( .A(n433), .B(n928), .C(n576), .Y(n901) );
  NAND2X1 U650 ( .A(N430), .B(n574), .Y(n576) );
  OAI21X1 U652 ( .A(n433), .B(n927), .C(n578), .Y(n902) );
  NAND2X1 U653 ( .A(N429), .B(n574), .Y(n578) );
  OAI21X1 U654 ( .A(n433), .B(n926), .C(n580), .Y(n903) );
  NAND2X1 U655 ( .A(N428), .B(n574), .Y(n580) );
  OAI21X1 U656 ( .A(n433), .B(n355), .C(n582), .Y(n904) );
  NAND2X1 U657 ( .A(N427), .B(n574), .Y(n582) );
  OAI21X1 U659 ( .A(n433), .B(n925), .C(n583), .Y(n905) );
  NAND2X1 U660 ( .A(N426), .B(n574), .Y(n583) );
  OAI21X1 U662 ( .A(n433), .B(n357), .C(n584), .Y(n906) );
  NAND2X1 U663 ( .A(N425), .B(n574), .Y(n584) );
  OAI21X1 U664 ( .A(n433), .B(n924), .C(n585), .Y(n907) );
  NAND2X1 U665 ( .A(N424), .B(n574), .Y(n585) );
  NOR2X1 U666 ( .A(n557), .B(n568), .Y(n574) );
  NOR2X1 U667 ( .A(n586), .B(n587), .Y(n568) );
  NAND3X1 U668 ( .A(si[7]), .B(si[6]), .C(n588), .Y(n587) );
  NOR2X1 U669 ( .A(n926), .B(n927), .Y(n588) );
  NAND3X1 U672 ( .A(si[3]), .B(si[2]), .C(n589), .Y(n586) );
  NOR2X1 U673 ( .A(n924), .B(n357), .Y(n589) );
  NAND3X1 U677 ( .A(n435), .B(n253), .C(n591), .Y(n590) );
  NOR2X1 U678 ( .A(n241), .B(n313), .Y(n591) );
  NOR2X1 U679 ( .A(n203), .B(n116), .Y(n313) );
  OAI21X1 U681 ( .A(n218), .B(n499), .C(n524), .Y(n593) );
  NAND3X1 U684 ( .A(n123), .B(n484), .C(n597), .Y(n596) );
  NOR2X1 U685 ( .A(n598), .B(n599), .Y(n597) );
  OAI21X1 U686 ( .A(n218), .B(n170), .C(n139), .Y(n599) );
  OAI21X1 U690 ( .A(n111), .B(n602), .C(n10), .Y(n63) );
  OAI21X1 U693 ( .A(n467), .B(n890), .C(n607), .Y(n908) );
  NAND2X1 U694 ( .A(N413), .B(n608), .Y(n607) );
  OAI21X1 U696 ( .A(n467), .B(n889), .C(n609), .Y(n909) );
  NAND2X1 U697 ( .A(N412), .B(n608), .Y(n609) );
  OAI21X1 U699 ( .A(n467), .B(n888), .C(n611), .Y(n910) );
  NAND2X1 U700 ( .A(N411), .B(n608), .Y(n611) );
  OAI21X1 U702 ( .A(n467), .B(n887), .C(n613), .Y(n911) );
  NAND2X1 U703 ( .A(N410), .B(n608), .Y(n613) );
  OAI21X1 U705 ( .A(n467), .B(n886), .C(n615), .Y(n912) );
  NAND2X1 U706 ( .A(N409), .B(n608), .Y(n615) );
  OAI21X1 U708 ( .A(n467), .B(n885), .C(n617), .Y(n913) );
  NAND2X1 U709 ( .A(N408), .B(n608), .Y(n617) );
  OAI21X1 U711 ( .A(n467), .B(n884), .C(n619), .Y(n914) );
  NAND2X1 U712 ( .A(N414), .B(n608), .Y(n619) );
  OAI21X1 U714 ( .A(n467), .B(n401), .C(n620), .Y(n915) );
  NAND2X1 U715 ( .A(N407), .B(n608), .Y(n620) );
  NOR2X1 U716 ( .A(n457), .B(n210), .Y(n608) );
  NAND3X1 U721 ( .A(n5), .B(n197), .C(n621), .Y(n457) );
  NOR2X1 U722 ( .A(n506), .B(n497), .Y(n621) );
  NAND3X1 U723 ( .A(n8), .B(n581), .C(n622), .Y(n497) );
  NOR2X1 U724 ( .A(n302), .B(n246), .Y(n622) );
  NOR2X1 U727 ( .A(n116), .B(n499), .Y(n171) );
  NOR2X1 U731 ( .A(n485), .B(n162), .Y(n232) );
  NOR2X1 U732 ( .A(n183), .B(n110), .Y(n162) );
  OAI21X1 U733 ( .A(n116), .B(n625), .C(n512), .Y(n485) );
  OAI21X1 U735 ( .A(n170), .B(n605), .C(n562), .Y(n627) );
  NOR2X1 U737 ( .A(n111), .B(n605), .Y(n149) );
  NAND3X1 U738 ( .A(n628), .B(n604), .C(n592), .Y(n197) );
  XOR2X1 U739 ( .A(n4), .B(n218), .Y(n628) );
  NAND2X1 U743 ( .A(n483), .B(n516), .Y(n225) );
  OAI21X1 U745 ( .A(n111), .B(n602), .C(n601), .Y(n631) );
  NAND2X1 U746 ( .A(n606), .B(n177), .Y(n601) );
  NOR2X1 U748 ( .A(n598), .B(n241), .Y(n483) );
  OAI21X1 U750 ( .A(n110), .B(n111), .C(n633), .Y(n598) );
  NOR2X1 U751 ( .A(n600), .B(n118), .Y(n633) );
  NOR2X1 U752 ( .A(n183), .B(n116), .Y(n118) );
  NAND2X1 U754 ( .A(n67), .B(n4), .Y(n198) );
  NOR2X1 U755 ( .A(n314), .B(n540), .Y(n233) );
  NOR2X1 U757 ( .A(n273), .B(n575), .Y(n139) );
  NAND3X1 U759 ( .A(n142), .B(n592), .C(n4), .Y(n634) );
  NOR2X1 U760 ( .A(n623), .B(n605), .Y(n273) );
  OAI21X1 U762 ( .A(n170), .B(n110), .C(n557), .Y(n635) );
  NOR2X1 U764 ( .A(n111), .B(n116), .Y(n567) );
  NAND2X1 U765 ( .A(n571), .B(n610), .Y(n111) );
  NAND2X1 U766 ( .A(state[0]), .B(n522), .Y(n170) );
  NAND2X1 U767 ( .A(n518), .B(n501), .Y(n140) );
  AOI21X1 U769 ( .A(n183), .B(n625), .C(n605), .Y(n156) );
  NOR2X1 U771 ( .A(n614), .B(state[2]), .Y(n142) );
  NAND3X1 U772 ( .A(n4), .B(n555), .C(state[0]), .Y(n183) );
  NAND2X1 U774 ( .A(n172), .B(n603), .Y(n157) );
  NAND2X1 U780 ( .A(n555), .B(n161), .Y(n148) );
  NOR2X1 U781 ( .A(n595), .B(n594), .Y(n478) );
  NAND2X1 U783 ( .A(n240), .B(n188), .Y(n199) );
  NOR2X1 U784 ( .A(n110), .B(n115), .Y(n67) );
  NAND3X1 U785 ( .A(n152), .B(n564), .C(n528), .Y(n595) );
  NOR2X1 U787 ( .A(n116), .B(n623), .Y(n205) );
  NAND3X1 U788 ( .A(n612), .B(n555), .C(n4), .Y(n623) );
  NAND2X1 U790 ( .A(n604), .B(n614), .Y(n116) );
  NAND2X1 U792 ( .A(n569), .B(n606), .Y(n564) );
  NAND2X1 U794 ( .A(state[2]), .B(n614), .Y(n110) );
  NAND2X1 U797 ( .A(n571), .B(n4), .Y(n625) );
  NAND2X1 U799 ( .A(state[0]), .B(state[1]), .Y(n153) );
  NAND2X1 U801 ( .A(n592), .B(n188), .Y(n499) );
  NAND2X1 U804 ( .A(state[1]), .B(n612), .Y(n115) );
  NAND2X1 U806 ( .A(state[2]), .B(n218), .Y(n602) );
  NAND3X1 U807 ( .A(n639), .B(n641), .C(n640), .Y(N479) );
  NOR2X1 U808 ( .A(n643), .B(n642), .Y(n641) );
  OAI22X1 U809 ( .A(n785), .B(n212), .C(n870), .D(n645), .Y(n643) );
  OAI22X1 U812 ( .A(n769), .B(n646), .C(n777), .D(n647), .Y(n642) );
  AOI22X1 U815 ( .A(n947), .B(\keyTable[5][0] ), .C(n946), .D(\keyTable[4][0] ), .Y(n640) );
  AOI22X1 U816 ( .A(n949), .B(\keyTable[7][0] ), .C(\keyTable[6][0] ), .D(n948), .Y(n639) );
  NAND3X1 U817 ( .A(n652), .B(n653), .C(n654), .Y(N478) );
  NOR2X1 U818 ( .A(n655), .B(n656), .Y(n654) );
  OAI22X1 U819 ( .A(n786), .B(n212), .C(n869), .D(n645), .Y(n656) );
  OAI22X1 U822 ( .A(n770), .B(n646), .C(n778), .D(n647), .Y(n655) );
  AOI22X1 U825 ( .A(n947), .B(\keyTable[5][1] ), .C(n946), .D(\keyTable[4][1] ), .Y(n653) );
  AOI22X1 U826 ( .A(n949), .B(\keyTable[7][1] ), .C(n948), .D(\keyTable[6][1] ), .Y(n652) );
  NAND3X1 U827 ( .A(n657), .B(n658), .C(n659), .Y(N477) );
  NOR2X1 U828 ( .A(n660), .B(n661), .Y(n659) );
  OAI22X1 U829 ( .A(n787), .B(n212), .C(n868), .D(n645), .Y(n661) );
  OAI22X1 U832 ( .A(n771), .B(n646), .C(n779), .D(n647), .Y(n660) );
  AOI22X1 U835 ( .A(n947), .B(\keyTable[5][2] ), .C(n946), .D(\keyTable[4][2] ), .Y(n658) );
  AOI22X1 U836 ( .A(n949), .B(\keyTable[7][2] ), .C(n948), .D(\keyTable[6][2] ), .Y(n657) );
  NAND3X1 U837 ( .A(n662), .B(n663), .C(n664), .Y(N476) );
  NOR2X1 U838 ( .A(n665), .B(n666), .Y(n664) );
  OAI22X1 U839 ( .A(n788), .B(n212), .C(n867), .D(n645), .Y(n666) );
  OAI22X1 U842 ( .A(n772), .B(n646), .C(n780), .D(n647), .Y(n665) );
  AOI22X1 U845 ( .A(n947), .B(\keyTable[5][3] ), .C(n946), .D(\keyTable[4][3] ), .Y(n663) );
  AOI22X1 U846 ( .A(n949), .B(\keyTable[7][3] ), .C(n948), .D(\keyTable[6][3] ), .Y(n662) );
  NAND3X1 U847 ( .A(n667), .B(n668), .C(n669), .Y(N475) );
  NOR2X1 U848 ( .A(n670), .B(n671), .Y(n669) );
  OAI22X1 U849 ( .A(n789), .B(n212), .C(n866), .D(n645), .Y(n671) );
  OAI22X1 U852 ( .A(n773), .B(n646), .C(n781), .D(n647), .Y(n670) );
  AOI22X1 U855 ( .A(n947), .B(\keyTable[5][4] ), .C(n946), .D(\keyTable[4][4] ), .Y(n668) );
  AOI22X1 U856 ( .A(n949), .B(\keyTable[7][4] ), .C(n948), .D(\keyTable[6][4] ), .Y(n667) );
  NAND3X1 U857 ( .A(n672), .B(n673), .C(n674), .Y(N474) );
  NOR2X1 U858 ( .A(n675), .B(n676), .Y(n674) );
  OAI22X1 U859 ( .A(n790), .B(n212), .C(n865), .D(n645), .Y(n676) );
  OAI22X1 U862 ( .A(n774), .B(n646), .C(n782), .D(n647), .Y(n675) );
  AOI22X1 U865 ( .A(n947), .B(\keyTable[5][5] ), .C(n946), .D(\keyTable[4][5] ), .Y(n673) );
  AOI22X1 U866 ( .A(n949), .B(\keyTable[7][5] ), .C(n948), .D(\keyTable[6][5] ), .Y(n672) );
  NAND3X1 U867 ( .A(n677), .B(n678), .C(n679), .Y(N473) );
  NOR2X1 U868 ( .A(n680), .B(n681), .Y(n679) );
  OAI22X1 U869 ( .A(n791), .B(n212), .C(n864), .D(n645), .Y(n681) );
  OAI22X1 U872 ( .A(n775), .B(n237), .C(n783), .D(n647), .Y(n680) );
  AOI22X1 U875 ( .A(n947), .B(\keyTable[5][6] ), .C(n946), .D(\keyTable[4][6] ), .Y(n678) );
  AOI22X1 U876 ( .A(n949), .B(\keyTable[7][6] ), .C(n948), .D(\keyTable[6][6] ), .Y(n677) );
  NAND3X1 U877 ( .A(n682), .B(n683), .C(n684), .Y(N472) );
  NOR2X1 U878 ( .A(n685), .B(n686), .Y(n684) );
  OAI22X1 U879 ( .A(n871), .B(n212), .C(n883), .D(n645), .Y(n686) );
  NAND3X1 U880 ( .A(n950), .B(n945), .C(n951), .Y(n645) );
  NAND3X1 U882 ( .A(n950), .B(keyi[0]), .C(n945), .Y(n644) );
  OAI22X1 U884 ( .A(n776), .B(n237), .C(n784), .D(n647), .Y(n685) );
  NAND3X1 U885 ( .A(n951), .B(n945), .C(keyi[1]), .Y(n647) );
  NAND3X1 U887 ( .A(keyi[1]), .B(n230), .C(n945), .Y(n646) );
  AOI22X1 U890 ( .A(n947), .B(\keyTable[5][7] ), .C(n946), .D(\keyTable[4][7] ), .Y(n683) );
  NAND3X1 U892 ( .A(n951), .B(n228), .C(n235), .Y(n687) );
  NAND3X1 U894 ( .A(n228), .B(n230), .C(n235), .Y(n688) );
  AOI22X1 U896 ( .A(n949), .B(\keyTable[7][7] ), .C(n948), .D(\keyTable[6][7] ), .Y(n682) );
  NAND3X1 U898 ( .A(n951), .B(keyi[1]), .C(n235), .Y(n689) );
  NAND3X1 U901 ( .A(keyi[1]), .B(n230), .C(n235), .Y(n690) );
  OR2X2 U105 ( .A(n119), .B(n120), .Y(nextState[4]) );
  OR2X2 U134 ( .A(n162), .B(n575), .Y(n166) );
  AND2X2 U142 ( .A(n130), .B(n186), .Y(n159) );
  AND2X2 U635 ( .A(n507), .B(n564), .Y(n563) );
  AND2X2 U692 ( .A(n603), .B(n501), .Y(n123) );
  OR2X2 U761 ( .A(n140), .B(n635), .Y(n314) );
  OR2X2 U775 ( .A(n602), .B(n623), .Y(n603) );
  OR2X2 U800 ( .A(n602), .B(n499), .Y(n152) );
  KSA_1_DW01_add_0 add_377 ( .A(temp), .B(extratemp), .CI(1'b0), .SUM({N527, 
        N526, N525, N524, N523, N522, N521, N520}) );
  KSA_1_DW01_add_1 add_337 ( .A(intj), .B(DATA_IN), .CI(1'b0), .SUM({N519, 
        N518, N517, N516, N515, N514, N513, N512}) );
  KSA_1_DW01_inc_0 add_289 ( .A(si), .SUM({N431, N430, N429, N428, N427, N426, 
        N425, N424}) );
  KSA_1_DW01_inc_1 add_263 ( .A(prefillCounter), .SUM({N414, N413, N412, N411, 
        N410, N409, N408, N407}) );
  KSA_1_DW01_inc_2 r126 ( .A(inti), .SUM({N503, N502, N501, N500, N499, N498, 
        N497, N496}) );
  KSA_1_DW01_add_3 add_1_root_add_0_root_add_302_2 ( .A(DATA_IN), .B(sj), .CI(
        1'b0), .SUM({N456, N455, N454, N453, N452, N451, N450, N449}) );
  KSA_1_DW01_add_2 add_0_root_add_0_root_add_302_2 ( .A({N472, N473, N474, 
        N475, N476, N477, N478, N479}), .B({N456, N455, N454, N453, N452, N451, 
        N450, N449}), .CI(1'b0), .SUM({N487, N486, N485, N484, N483, N482, 
        N481, N480}) );
  TBUFX1 \nfaddr_tri[5]  ( .A(n703), .EN(n253), .Y(nfaddr[5]) );
  TBUFX1 \nfaddr_tri[0]  ( .A(n708), .EN(n253), .Y(nfaddr[0]) );
  TBUFX1 \nfaddr_tri[1]  ( .A(n707), .EN(n253), .Y(nfaddr[1]) );
  TBUFX1 \nfaddr_tri[2]  ( .A(n706), .EN(n253), .Y(nfaddr[2]) );
  TBUFX1 \nfaddr_tri[3]  ( .A(n705), .EN(n253), .Y(nfaddr[3]) );
  TBUFX1 \nfaddr_tri[4]  ( .A(n704), .EN(n253), .Y(nfaddr[4]) );
  TBUFX1 \nfaddr_tri[6]  ( .A(n702), .EN(n253), .Y(nfaddr[6]) );
  TBUFX1 \nfaddr_tri[7]  ( .A(n700), .EN(n253), .Y(nfaddr[7]) );
  TBUFX1 \nfdata_tri[0]  ( .A(n699), .EN(n581), .Y(nfdata[0]) );
  TBUFX1 \nfdata_tri[1]  ( .A(n698), .EN(n581), .Y(nfdata[1]) );
  TBUFX1 \nfdata_tri[2]  ( .A(n697), .EN(n581), .Y(nfdata[2]) );
  TBUFX1 \nfdata_tri[3]  ( .A(n696), .EN(n581), .Y(nfdata[3]) );
  TBUFX1 \nfdata_tri[4]  ( .A(n695), .EN(n581), .Y(nfdata[4]) );
  TBUFX1 \nfdata_tri[5]  ( .A(n694), .EN(n581), .Y(nfdata[5]) );
  TBUFX1 \nfdata_tri[6]  ( .A(n693), .EN(n581), .Y(nfdata[6]) );
  TBUFX1 \nfdata_tri[7]  ( .A(n691), .EN(n581), .Y(nfdata[7]) );
  DFFSR PDATA_READY_reg ( .D(n540), .CLK(CLK), .R(n292), .S(1'b1), .Q(
        PDATA_READY) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n292), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[4]  ( .D(nextState[4]), .CLK(CLK), .R(n292), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[3]  ( .D(nextState[3]), .CLK(CLK), .R(n292), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n292), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n292), .S(1'b1), .Q(
        state[0]) );
  DFFSR \si_reg[7]  ( .D(n900), .CLK(CLK), .R(n292), .S(1'b1), .Q(si[7]) );
  DFFSR \si_reg[6]  ( .D(n901), .CLK(CLK), .R(n292), .S(1'b1), .Q(si[6]) );
  DFFSR \si_reg[5]  ( .D(n902), .CLK(CLK), .R(n292), .S(1'b1), .Q(si[5]) );
  DFFSR \si_reg[4]  ( .D(n903), .CLK(CLK), .R(n292), .S(1'b1), .Q(si[4]) );
  DFFSR \si_reg[3]  ( .D(n904), .CLK(CLK), .R(n292), .S(1'b1), .Q(si[3]) );
  DFFSR \si_reg[2]  ( .D(n905), .CLK(CLK), .R(n292), .S(1'b1), .Q(si[2]) );
  DFFSR \si_reg[1]  ( .D(n906), .CLK(CLK), .R(n292), .S(1'b1), .Q(si[1]) );
  DFFSR \si_reg[0]  ( .D(n907), .CLK(CLK), .R(n292), .S(1'b1), .Q(si[0]) );
  DFFSR \sj_reg[4]  ( .D(n895), .CLK(CLK), .R(n292), .S(1'b1), .Q(sj[4]) );
  DFFSR \sj_reg[3]  ( .D(n894), .CLK(CLK), .R(n292), .S(1'b1), .Q(sj[3]) );
  DFFSR \sj_reg[2]  ( .D(n893), .CLK(CLK), .R(n292), .S(1'b1), .Q(sj[2]) );
  DFFSR \sj_reg[1]  ( .D(n892), .CLK(CLK), .R(n292), .S(1'b1), .Q(sj[1]) );
  DFFSR \sj_reg[0]  ( .D(n891), .CLK(CLK), .R(n292), .S(1'b1), .Q(sj[0]) );
  DFFSR \sj_reg[5]  ( .D(n896), .CLK(CLK), .R(n292), .S(1'b1), .Q(sj[5]) );
  DFFSR \currentProcessedData_reg[7]  ( .D(nextProcessedData[7]), .CLK(CLK), 
        .R(n292), .S(1'b1), .Q(currentProcessedData[7]) );
  DFFSR \currentProcessedData_reg[6]  ( .D(nextProcessedData[6]), .CLK(CLK), 
        .R(n292), .S(1'b1), .Q(currentProcessedData[6]) );
  DFFSR \currentProcessedData_reg[5]  ( .D(nextProcessedData[5]), .CLK(CLK), 
        .R(n292), .S(1'b1), .Q(currentProcessedData[5]) );
  DFFSR \currentProcessedData_reg[4]  ( .D(nextProcessedData[4]), .CLK(CLK), 
        .R(n292), .S(1'b1), .Q(currentProcessedData[4]) );
  DFFSR \currentProcessedData_reg[3]  ( .D(nextProcessedData[3]), .CLK(CLK), 
        .R(n292), .S(1'b1), .Q(currentProcessedData[3]) );
  DFFSR \currentProcessedData_reg[2]  ( .D(nextProcessedData[2]), .CLK(CLK), 
        .R(n292), .S(1'b1), .Q(currentProcessedData[2]) );
  DFFSR \currentProcessedData_reg[1]  ( .D(nextProcessedData[1]), .CLK(CLK), 
        .R(n292), .S(1'b1), .Q(currentProcessedData[1]) );
  DFFSR \currentProcessedData_reg[0]  ( .D(nextProcessedData[0]), .CLK(CLK), 
        .R(n292), .S(1'b1), .Q(currentProcessedData[0]) );
  DFFSR \sj_reg[6]  ( .D(n897), .CLK(CLK), .R(n292), .S(1'b1), .Q(sj[6]) );
  DFFSR \sj_reg[7]  ( .D(n898), .CLK(CLK), .R(n292), .S(1'b1), .Q(sj[7]) );
  BUFX4 U4 ( .A(n232), .Y(n3) );
  OR2X1 U11 ( .A(n602), .B(n170), .Y(n12) );
  INVX4 U16 ( .A(n7), .Y(n261) );
  INVX2 U21 ( .A(n688), .Y(n947) );
  INVX2 U26 ( .A(n687), .Y(n946) );
  INVX2 U31 ( .A(n602), .Y(n175) );
  INVX2 U36 ( .A(n12), .Y(n241) );
  INVX2 U41 ( .A(n255), .Y(n256) );
  INVX2 U45 ( .A(n477), .Y(n469) );
  BUFX2 U103 ( .A(state[4]), .Y(n4) );
  AND2X2 U107 ( .A(n233), .B(n9), .Y(n5) );
  AND2X2 U136 ( .A(n409), .B(n172), .Y(n6) );
  AND2X2 U141 ( .A(n233), .B(n520), .Y(n7) );
  INVX2 U144 ( .A(n10), .Y(n246) );
  OR2X2 U155 ( .A(n201), .B(n605), .Y(n8) );
  AND2X2 U157 ( .A(n504), .B(n478), .Y(n9) );
  OR2X2 U190 ( .A(n110), .B(n623), .Y(n10) );
  AND2X2 U194 ( .A(n162), .B(n469), .Y(n14) );
  INVX2 U198 ( .A(n258), .Y(n259) );
  INVX2 U199 ( .A(keyi[1]), .Y(n950) );
  INVX2 U201 ( .A(n8), .Y(n244) );
  AND2X2 U202 ( .A(n8), .B(n601), .Y(n15) );
  AND2X2 U204 ( .A(n529), .B(n528), .Y(n16) );
  INVX2 U205 ( .A(n249), .Y(n250) );
  INVX4 U207 ( .A(RST), .Y(n292) );
  INVX1 U281 ( .A(n241), .Y(n507) );
  BUFX4 U284 ( .A(n644), .Y(n212) );
  INVX1 U288 ( .A(n4), .Y(n161) );
  INVX1 U291 ( .A(n4), .Y(n610) );
  NAND2X1 U295 ( .A(n175), .B(n177), .Y(n172) );
  INVX1 U298 ( .A(n172), .Y(n127) );
  AND2X1 U302 ( .A(n522), .B(n612), .Y(n177) );
  BUFX2 U305 ( .A(n206), .Y(n180) );
  INVX2 U309 ( .A(n5), .Y(n185) );
  INVX2 U312 ( .A(n196), .Y(n484) );
  INVX1 U316 ( .A(n610), .Y(n187) );
  INVX2 U317 ( .A(n187), .Y(n188) );
  NAND3X1 U320 ( .A(n249), .B(n197), .C(n15), .Y(n196) );
  INVX1 U321 ( .A(n15), .Y(n252) );
  NAND2X1 U323 ( .A(n527), .B(n16), .Y(n526) );
  NAND2X1 U325 ( .A(n522), .B(n612), .Y(n201) );
  NAND2X1 U327 ( .A(n522), .B(n612), .Y(n203) );
  INVX2 U329 ( .A(n142), .Y(n605) );
  INVX2 U331 ( .A(n326), .Y(n297) );
  INVX2 U333 ( .A(n318), .Y(n300) );
  INVX2 U335 ( .A(n311), .Y(n305) );
  INVX2 U337 ( .A(n317), .Y(n302) );
  INVX2 U338 ( .A(n327), .Y(n295) );
  BUFX2 U341 ( .A(n265), .Y(n275) );
  BUFX2 U344 ( .A(n264), .Y(n270) );
  BUFX2 U347 ( .A(n264), .Y(n268) );
  BUFX2 U350 ( .A(n264), .Y(n271) );
  BUFX2 U353 ( .A(n265), .Y(n277) );
  BUFX2 U356 ( .A(n265), .Y(n280) );
  BUFX2 U359 ( .A(n267), .Y(n282) );
  BUFX2 U362 ( .A(n267), .Y(n285) );
  BUFX2 U365 ( .A(n267), .Y(n287) );
  BUFX2 U368 ( .A(n333), .Y(n329) );
  BUFX2 U371 ( .A(n335), .Y(n327) );
  BUFX2 U374 ( .A(n307), .Y(n326) );
  BUFX2 U377 ( .A(n335), .Y(n318) );
  BUFX2 U380 ( .A(n307), .Y(n317) );
  BUFX2 U383 ( .A(n337), .Y(n311) );
  BUFX2 U386 ( .A(n337), .Y(n307) );
  BUFX2 U389 ( .A(n333), .Y(n331) );
  INVX2 U392 ( .A(n171), .Y(n581) );
  INVX4 U395 ( .A(n6), .Y(n262) );
  NOR2X1 U398 ( .A(n477), .B(n478), .Y(n206) );
  BUFX2 U401 ( .A(n328), .Y(n265) );
  BUFX2 U404 ( .A(n328), .Y(n267) );
  BUFX2 U407 ( .A(n328), .Y(n264) );
  INVX2 U410 ( .A(n290), .Y(n335) );
  INVX2 U413 ( .A(n290), .Y(n333) );
  INVX2 U416 ( .A(n290), .Y(n337) );
  INVX2 U419 ( .A(n199), .Y(n594) );
  INVX2 U422 ( .A(n559), .Y(n407) );
  INVX2 U425 ( .A(n487), .Y(n258) );
  INVX2 U428 ( .A(n210), .Y(n247) );
  INVX2 U431 ( .A(n208), .Y(n253) );
  INVX2 U434 ( .A(n292), .Y(n290) );
  INVX2 U502 ( .A(n197), .Y(n572) );
  INVX2 U505 ( .A(n689), .Y(n948) );
  OR2X2 U508 ( .A(n506), .B(n593), .Y(n208) );
  OR2X2 U511 ( .A(n170), .B(n116), .Y(n210) );
  INVX2 U514 ( .A(n239), .Y(n240) );
  INVX2 U517 ( .A(n63), .Y(n249) );
  INVX2 U520 ( .A(n690), .Y(n949) );
  INVX2 U523 ( .A(n634), .Y(n575) );
  INVX2 U524 ( .A(keyi[2]), .Y(n945) );
  BUFX2 U525 ( .A(keyi[2]), .Y(n235) );
  BUFX2 U526 ( .A(n950), .Y(n228) );
  BUFX2 U529 ( .A(n532), .Y(n214) );
  BUFX2 U531 ( .A(n532), .Y(n216) );
  BUFX2 U533 ( .A(state[3]), .Y(n218) );
  INVX2 U535 ( .A(sj[0]), .Y(n220) );
  INVX2 U537 ( .A(keyi[0]), .Y(n951) );
  BUFX2 U539 ( .A(keyi[0]), .Y(n230) );
  BUFX2 U541 ( .A(n646), .Y(n237) );
  INVX2 U543 ( .A(n531), .Y(n255) );
  INVX1 U545 ( .A(n457), .Y(n467) );
  INVX2 U547 ( .A(n67), .Y(n239) );
  OR2X2 U549 ( .A(n407), .B(n938), .Y(n238) );
  NAND2X1 U554 ( .A(n238), .B(n558), .Y(n898) );
  INVX1 U558 ( .A(n110), .Y(n606) );
  INVX4 U562 ( .A(n526), .Y(n409) );
  NAND2X1 U565 ( .A(n357), .B(n924), .Y(n339) );
  OAI21X1 U568 ( .A(n924), .B(n357), .C(n339), .Y(N442) );
  NOR2X1 U571 ( .A(n339), .B(si[2]), .Y(n343) );
  AOI21X1 U574 ( .A(n339), .B(si[2]), .C(n343), .Y(n341) );
  NAND2X1 U577 ( .A(n343), .B(n355), .Y(n345) );
  OAI21X1 U580 ( .A(n343), .B(n355), .C(n345), .Y(N444) );
  NOR2X1 U584 ( .A(n345), .B(si[4]), .Y(n349) );
  AOI21X1 U585 ( .A(n345), .B(si[4]), .C(n349), .Y(n347) );
  NAND2X1 U586 ( .A(n349), .B(n927), .Y(n351) );
  OAI21X1 U588 ( .A(n349), .B(n927), .C(n351), .Y(N446) );
  XNOR2X1 U590 ( .A(si[6]), .B(n351), .Y(N447) );
  NOR2X1 U592 ( .A(si[6]), .B(n351), .Y(n353) );
  XOR2X1 U594 ( .A(si[7]), .B(n353), .Y(N448) );
  INVX2 U596 ( .A(si[3]), .Y(n355) );
  INVX2 U598 ( .A(si[1]), .Y(n357) );
  INVX2 U600 ( .A(n347), .Y(N445) );
  INVX2 U602 ( .A(n341), .Y(N443) );
  INVX2 U608 ( .A(KEY_ERROR), .Y(n359) );
  INVX2 U611 ( .A(BYTE_READY), .Y(n361) );
  INVX2 U614 ( .A(n130), .Y(n363) );
  INVX2 U617 ( .A(OPCODE[1]), .Y(n365) );
  INVX2 U620 ( .A(OPCODE[0]), .Y(n367) );
  INVX2 U623 ( .A(nextProcessedData[7]), .Y(n369) );
  INVX2 U626 ( .A(n316), .Y(n371) );
  INVX2 U627 ( .A(nextProcessedData[6]), .Y(n373) );
  INVX2 U629 ( .A(n325), .Y(n375) );
  INVX2 U630 ( .A(nextProcessedData[5]), .Y(n377) );
  INVX2 U636 ( .A(n324), .Y(n379) );
  INVX2 U640 ( .A(nextProcessedData[4]), .Y(n381) );
  INVX2 U642 ( .A(n323), .Y(n383) );
  INVX2 U644 ( .A(nextProcessedData[3]), .Y(n385) );
  INVX2 U645 ( .A(n322), .Y(n387) );
  INVX2 U648 ( .A(nextProcessedData[2]), .Y(n389) );
  INVX2 U651 ( .A(n321), .Y(n391) );
  INVX2 U658 ( .A(nextProcessedData[1]), .Y(n393) );
  INVX2 U661 ( .A(n320), .Y(n395) );
  INVX2 U670 ( .A(nextProcessedData[0]), .Y(n397) );
  INVX2 U671 ( .A(n319), .Y(n399) );
  INVX2 U674 ( .A(prefillCounter[0]), .Y(n401) );
  INVX2 U675 ( .A(nfdata[0]), .Y(n403) );
  INVX2 U676 ( .A(nfaddr[0]), .Y(n405) );
  INVX2 U680 ( .A(n539), .Y(n411) );
  INVX2 U682 ( .A(n538), .Y(n413) );
  INVX2 U683 ( .A(n537), .Y(n415) );
  INVX2 U687 ( .A(n536), .Y(n417) );
  INVX2 U688 ( .A(n535), .Y(n419) );
  INVX2 U689 ( .A(n534), .Y(n421) );
  INVX2 U691 ( .A(n533), .Y(n423) );
  INVX2 U695 ( .A(n530), .Y(n425) );
  INVX2 U698 ( .A(n508), .Y(n427) );
  INVX2 U701 ( .A(n502), .Y(n429) );
  INVX2 U704 ( .A(n570), .Y(n431) );
  INVX2 U707 ( .A(n590), .Y(n433) );
  INVX2 U710 ( .A(n596), .Y(n435) );
  INVX2 U713 ( .A(nfdata[7]), .Y(n437) );
  INVX2 U717 ( .A(nfdata[6]), .Y(n439) );
  INVX2 U718 ( .A(nfdata[5]), .Y(n441) );
  INVX2 U719 ( .A(nfdata[4]), .Y(n443) );
  INVX2 U720 ( .A(nfdata[3]), .Y(n445) );
  INVX2 U725 ( .A(nfdata[2]), .Y(n447) );
  INVX2 U726 ( .A(nfdata[1]), .Y(n449) );
  INVX2 U728 ( .A(n56), .Y(n451) );
  INVX2 U729 ( .A(n486), .Y(n453) );
  INVX2 U730 ( .A(n489), .Y(n455) );
  INVX2 U734 ( .A(n490), .Y(n458) );
  INVX2 U736 ( .A(n491), .Y(n459) );
  INVX2 U740 ( .A(n492), .Y(n461) );
  INVX2 U741 ( .A(n493), .Y(n462) );
  INVX2 U742 ( .A(n494), .Y(n463) );
  INVX2 U744 ( .A(n495), .Y(n465) );
  INVX2 U747 ( .A(nfaddr[1]), .Y(n471) );
  INVX2 U749 ( .A(nfaddr[2]), .Y(n473) );
  INVX2 U753 ( .A(nfaddr[3]), .Y(n475) );
  INVX2 U756 ( .A(nfaddr[4]), .Y(n480) );
  INVX2 U758 ( .A(nfaddr[5]), .Y(n482) );
  INVX2 U763 ( .A(nfaddr[6]), .Y(n488) );
  INVX2 U768 ( .A(nfaddr[7]), .Y(n498) );
  INVX2 U770 ( .A(n310), .Y(n500) );
  INVX2 U773 ( .A(n156), .Y(n501) );
  INVX2 U776 ( .A(n118), .Y(n503) );
  INVX2 U777 ( .A(n225), .Y(n504) );
  INVX2 U778 ( .A(n315), .Y(n505) );
  INVX2 U779 ( .A(n3), .Y(n506) );
  INVX2 U782 ( .A(n485), .Y(n509) );
  INVX2 U786 ( .A(n627), .Y(n512) );
  INVX2 U789 ( .A(n229), .Y(n514) );
  INVX2 U791 ( .A(n631), .Y(n516) );
  INVX2 U793 ( .A(n157), .Y(n518) );
  INVX2 U795 ( .A(n313), .Y(n520) );
  INVX2 U796 ( .A(n148), .Y(n522) );
  INVX2 U798 ( .A(n595), .Y(n524) );
  INVX2 U802 ( .A(n205), .Y(n528) );
  INVX2 U803 ( .A(n139), .Y(n540) );
  INVX2 U805 ( .A(n53), .Y(n541) );
  INVX2 U810 ( .A(n48), .Y(n542) );
  INVX2 U811 ( .A(n43), .Y(n543) );
  INVX2 U813 ( .A(n38), .Y(n545) );
  INVX2 U814 ( .A(n33), .Y(n547) );
  INVX2 U820 ( .A(n28), .Y(n549) );
  INVX2 U821 ( .A(n23), .Y(n551) );
  INVX2 U823 ( .A(n13), .Y(n553) );
  INVX2 U824 ( .A(state[1]), .Y(n555) );
  INVX2 U830 ( .A(n567), .Y(n557) );
  INVX2 U831 ( .A(n149), .Y(n562) );
  INVX2 U833 ( .A(n625), .Y(n569) );
  INVX2 U834 ( .A(n153), .Y(n571) );
  INVX2 U840 ( .A(n112), .Y(n577) );
  INVX2 U841 ( .A(n499), .Y(n579) );
  INVX2 U843 ( .A(n115), .Y(n592) );
  INVX2 U844 ( .A(n198), .Y(n600) );
  INVX2 U850 ( .A(state[2]), .Y(n604) );
  INVX2 U851 ( .A(state[0]), .Y(n612) );
  INVX2 U853 ( .A(state[3]), .Y(n614) );
  INVX2 U854 ( .A(\keyTable[7][0] ), .Y(n616) );
  INVX2 U860 ( .A(\keyTable[7][1] ), .Y(n618) );
  INVX2 U861 ( .A(\keyTable[7][2] ), .Y(n624) );
  INVX2 U863 ( .A(\keyTable[7][3] ), .Y(n626) );
  INVX2 U864 ( .A(\keyTable[7][4] ), .Y(n629) );
  INVX2 U870 ( .A(\keyTable[7][5] ), .Y(n630) );
  INVX2 U871 ( .A(\keyTable[7][6] ), .Y(n632) );
  INVX2 U873 ( .A(\keyTable[7][7] ), .Y(n636) );
  INVX2 U874 ( .A(\keyTable[6][0] ), .Y(n637) );
  INVX2 U881 ( .A(\keyTable[6][1] ), .Y(n638) );
  INVX2 U883 ( .A(\keyTable[6][2] ), .Y(n648) );
  INVX2 U886 ( .A(\keyTable[6][3] ), .Y(n649) );
  INVX2 U888 ( .A(\keyTable[6][4] ), .Y(n650) );
  INVX2 U889 ( .A(\keyTable[6][5] ), .Y(n651) );
  INVX2 U891 ( .A(\keyTable[6][6] ), .Y(n692) );
  INVX2 U893 ( .A(\keyTable[6][7] ), .Y(n701) );
  INVX2 U895 ( .A(\keyTable[5][0] ), .Y(n746) );
  INVX2 U897 ( .A(\keyTable[5][1] ), .Y(n748) );
  INVX2 U899 ( .A(\keyTable[5][2] ), .Y(n750) );
  INVX2 U900 ( .A(\keyTable[5][3] ), .Y(n752) );
  INVX2 U902 ( .A(\keyTable[5][4] ), .Y(n754) );
  INVX2 U903 ( .A(\keyTable[5][5] ), .Y(n756) );
  INVX2 U904 ( .A(\keyTable[5][6] ), .Y(n758) );
  INVX2 U905 ( .A(\keyTable[5][7] ), .Y(n760) );
  INVX2 U906 ( .A(\keyTable[4][0] ), .Y(n761) );
  INVX2 U907 ( .A(\keyTable[4][1] ), .Y(n762) );
  INVX2 U908 ( .A(\keyTable[4][2] ), .Y(n763) );
  INVX2 U909 ( .A(\keyTable[4][3] ), .Y(n764) );
  INVX2 U910 ( .A(\keyTable[4][4] ), .Y(n765) );
  INVX2 U911 ( .A(\keyTable[4][5] ), .Y(n766) );
  INVX2 U912 ( .A(\keyTable[4][6] ), .Y(n767) );
  INVX2 U913 ( .A(\keyTable[4][7] ), .Y(n768) );
  INVX2 U914 ( .A(\keyTable[3][0] ), .Y(n769) );
  INVX2 U915 ( .A(\keyTable[3][1] ), .Y(n770) );
  INVX2 U916 ( .A(\keyTable[3][2] ), .Y(n771) );
  INVX2 U917 ( .A(\keyTable[3][3] ), .Y(n772) );
  INVX2 U918 ( .A(\keyTable[3][4] ), .Y(n773) );
  INVX2 U919 ( .A(\keyTable[3][5] ), .Y(n774) );
  INVX2 U920 ( .A(\keyTable[3][6] ), .Y(n775) );
  INVX2 U921 ( .A(\keyTable[3][7] ), .Y(n776) );
  INVX2 U922 ( .A(\keyTable[2][0] ), .Y(n777) );
  INVX2 U923 ( .A(\keyTable[2][1] ), .Y(n778) );
  INVX2 U924 ( .A(\keyTable[2][2] ), .Y(n779) );
  INVX2 U925 ( .A(\keyTable[2][3] ), .Y(n780) );
  INVX2 U926 ( .A(\keyTable[2][4] ), .Y(n781) );
  INVX2 U927 ( .A(\keyTable[2][5] ), .Y(n782) );
  INVX2 U928 ( .A(\keyTable[2][6] ), .Y(n783) );
  INVX2 U929 ( .A(\keyTable[2][7] ), .Y(n784) );
  INVX2 U930 ( .A(\keyTable[1][0] ), .Y(n785) );
  INVX2 U931 ( .A(\keyTable[1][1] ), .Y(n786) );
  INVX2 U932 ( .A(\keyTable[1][2] ), .Y(n787) );
  INVX2 U933 ( .A(\keyTable[1][3] ), .Y(n788) );
  INVX2 U934 ( .A(\keyTable[1][4] ), .Y(n789) );
  INVX2 U935 ( .A(\keyTable[1][5] ), .Y(n790) );
  INVX2 U936 ( .A(\keyTable[1][6] ), .Y(n791) );
  INVX2 U937 ( .A(\keyTable[0][6] ), .Y(n864) );
  INVX2 U938 ( .A(\keyTable[0][5] ), .Y(n865) );
  INVX2 U939 ( .A(\keyTable[0][4] ), .Y(n866) );
  INVX2 U940 ( .A(\keyTable[0][3] ), .Y(n867) );
  INVX2 U941 ( .A(\keyTable[0][2] ), .Y(n868) );
  INVX2 U942 ( .A(\keyTable[0][1] ), .Y(n869) );
  INVX2 U943 ( .A(\keyTable[0][0] ), .Y(n870) );
  INVX2 U944 ( .A(\keyTable[1][7] ), .Y(n871) );
  INVX2 U945 ( .A(\keyTable[0][7] ), .Y(n883) );
  INVX2 U946 ( .A(prefillCounter[7]), .Y(n884) );
  INVX2 U947 ( .A(prefillCounter[1]), .Y(n885) );
  INVX2 U948 ( .A(prefillCounter[2]), .Y(n886) );
  INVX2 U949 ( .A(prefillCounter[3]), .Y(n887) );
  INVX2 U950 ( .A(prefillCounter[4]), .Y(n888) );
  INVX2 U951 ( .A(prefillCounter[5]), .Y(n889) );
  INVX2 U952 ( .A(prefillCounter[6]), .Y(n890) );
  INVX2 U953 ( .A(temp[7]), .Y(n916) );
  INVX2 U954 ( .A(temp[0]), .Y(n917) );
  INVX2 U955 ( .A(temp[1]), .Y(n918) );
  INVX2 U956 ( .A(temp[2]), .Y(n919) );
  INVX2 U957 ( .A(temp[3]), .Y(n920) );
  INVX2 U958 ( .A(temp[4]), .Y(n921) );
  INVX2 U959 ( .A(temp[5]), .Y(n922) );
  INVX2 U960 ( .A(temp[6]), .Y(n923) );
  INVX2 U961 ( .A(si[0]), .Y(n924) );
  INVX2 U962 ( .A(si[2]), .Y(n925) );
  INVX2 U963 ( .A(si[4]), .Y(n926) );
  INVX2 U964 ( .A(si[5]), .Y(n927) );
  INVX2 U965 ( .A(si[6]), .Y(n928) );
  INVX2 U966 ( .A(si[7]), .Y(n929) );
  INVX2 U967 ( .A(intj[7]), .Y(n930) );
  INVX2 U968 ( .A(intj[0]), .Y(n931) );
  INVX2 U969 ( .A(intj[1]), .Y(n932) );
  INVX2 U970 ( .A(intj[2]), .Y(n933) );
  INVX2 U971 ( .A(intj[3]), .Y(n934) );
  INVX2 U972 ( .A(intj[4]), .Y(n935) );
  INVX2 U973 ( .A(intj[5]), .Y(n936) );
  INVX2 U974 ( .A(intj[6]), .Y(n937) );
  INVX2 U975 ( .A(sj[7]), .Y(n938) );
  INVX2 U976 ( .A(sj[6]), .Y(n939) );
  INVX2 U977 ( .A(sj[5]), .Y(n940) );
  INVX2 U978 ( .A(sj[4]), .Y(n941) );
  INVX2 U979 ( .A(sj[3]), .Y(n942) );
  INVX2 U980 ( .A(sj[2]), .Y(n943) );
  INVX2 U981 ( .A(sj[1]), .Y(n944) );
  INVX2 U982 ( .A(currentProcessedData[0]), .Y(n952) );
  INVX2 U983 ( .A(currentProcessedData[1]), .Y(n953) );
  INVX2 U984 ( .A(currentProcessedData[2]), .Y(n954) );
  INVX2 U985 ( .A(currentProcessedData[3]), .Y(n955) );
  INVX2 U986 ( .A(currentProcessedData[4]), .Y(n956) );
  INVX2 U987 ( .A(currentProcessedData[5]), .Y(n957) );
  INVX2 U988 ( .A(currentProcessedData[6]), .Y(n958) );
  INVX2 U989 ( .A(currentProcessedData[7]), .Y(n959) );
  INVX2 U990 ( .A(faddr[7]), .Y(n960) );
  INVX2 U991 ( .A(faddr[6]), .Y(n961) );
  INVX2 U992 ( .A(faddr[5]), .Y(n962) );
  INVX2 U993 ( .A(faddr[4]), .Y(n963) );
  INVX2 U994 ( .A(faddr[3]), .Y(n964) );
  INVX2 U995 ( .A(faddr[2]), .Y(n965) );
  INVX2 U996 ( .A(faddr[1]), .Y(n966) );
  INVX2 U997 ( .A(faddr[0]), .Y(n967) );
  INVX2 U998 ( .A(fdata[7]), .Y(n968) );
  INVX2 U999 ( .A(fdata[6]), .Y(n969) );
  INVX2 U1000 ( .A(fdata[5]), .Y(n970) );
  INVX2 U1001 ( .A(fdata[4]), .Y(n971) );
  INVX2 U1002 ( .A(fdata[3]), .Y(n972) );
  INVX2 U1003 ( .A(fdata[2]), .Y(n973) );
  INVX2 U1004 ( .A(fdata[1]), .Y(n974) );
  INVX2 U1005 ( .A(fdata[0]), .Y(n975) );
endmodule


module uart_edge_detector_1 ( CLK, RST, SERIAL_IN, START_BIT );
  input CLK, RST, SERIAL_IN;
  output START_BIT;
  wire   Q_int, Q_int2, n2, n4;

  DFFSR Q_int_reg ( .D(SERIAL_IN), .CLK(CLK), .R(n2), .S(1'b1), .Q(Q_int) );
  NOR2X1 U7 ( .A(Q_int), .B(n4), .Y(START_BIT) );
  DFFSR Q_int2_reg ( .D(Q_int), .CLK(CLK), .R(n2), .S(1'b1), .Q(Q_int2) );
  INVX2 U4 ( .A(RST), .Y(n2) );
  INVX2 U6 ( .A(Q_int2), .Y(n4) );
endmodule


module uart_error_1 ( RST, CLK, RBUF_FULL, CHK_ERROR, OE );
  input RST, CLK, RBUF_FULL, CHK_ERROR;
  output OE;
  wire   OE_prime, n2;

  AND2X2 U5 ( .A(RBUF_FULL), .B(CHK_ERROR), .Y(OE_prime) );
  DFFSR OE_reg ( .D(OE_prime), .CLK(CLK), .R(n2), .S(1'b1), .Q(OE) );
  INVX2 U4 ( .A(RST), .Y(n2) );
endmodule


module uart_rcu_1 ( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT, RBUF_LOAD, 
        TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR );
  input CLK, RST, START_BIT, STOP_RCVING, SB_DETECT;
  output RBUF_LOAD, TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR;
  wire   timerRunning, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N99, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, \add_46/carry[7] ,
         \add_46/carry[6] , \add_46/carry[5] , \add_46/carry[4] ,
         \add_46/carry[3] , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47;
  wire   [2:0] state;
  wire   [7:0] count;
  wire   [7:0] nextCount;
  wire   [2:0] nextState;

  DFFSR \nextCount_reg[0]  ( .D(N31), .CLK(CLK), .R(1'b1), .S(n27), .Q(
        nextCount[0]) );
  AND2X2 U33 ( .A(N30), .B(timerRunning), .Y(N38) );
  AND2X2 U34 ( .A(N29), .B(timerRunning), .Y(N37) );
  AND2X2 U35 ( .A(N28), .B(timerRunning), .Y(N36) );
  AND2X2 U36 ( .A(N27), .B(timerRunning), .Y(N35) );
  AND2X2 U37 ( .A(N26), .B(timerRunning), .Y(N34) );
  AND2X2 U38 ( .A(N25), .B(timerRunning), .Y(N33) );
  AND2X2 U39 ( .A(N24), .B(timerRunning), .Y(N32) );
  OAI21X1 U54 ( .A(n49), .B(n43), .C(n50), .Y(n48) );
  OAI21X1 U55 ( .A(n44), .B(n42), .C(n43), .Y(n50) );
  NAND2X1 U56 ( .A(n51), .B(n52), .Y(n74) );
  OAI21X1 U57 ( .A(n53), .B(n54), .C(timerRunning), .Y(n52) );
  NAND2X1 U58 ( .A(n55), .B(n56), .Y(n54) );
  NAND2X1 U59 ( .A(n57), .B(n56), .Y(n75) );
  NAND3X1 U60 ( .A(n35), .B(n51), .C(CHK_ERROR), .Y(n57) );
  OAI21X1 U61 ( .A(n58), .B(n47), .C(n59), .Y(n76) );
  NAND2X1 U62 ( .A(n56), .B(n60), .Y(n58) );
  NAND2X1 U63 ( .A(n61), .B(n38), .Y(n56) );
  NAND3X1 U64 ( .A(n62), .B(n63), .C(n64), .Y(n77) );
  NAND3X1 U65 ( .A(n34), .B(n51), .C(SET_RBUF_FULL), .Y(n64) );
  NAND2X1 U66 ( .A(n60), .B(n63), .Y(n53) );
  NAND3X1 U67 ( .A(nextState[0]), .B(nextState[1]), .C(n61), .Y(n63) );
  NAND3X1 U68 ( .A(n36), .B(n38), .C(n61), .Y(n62) );
  OAI21X1 U69 ( .A(n65), .B(n45), .C(n51), .Y(n78) );
  OAI21X1 U70 ( .A(n65), .B(n46), .C(n51), .Y(n79) );
  NAND2X1 U71 ( .A(n60), .B(n59), .Y(n65) );
  NAND3X1 U72 ( .A(nextState[1]), .B(n36), .C(n39), .Y(n59) );
  NAND2X1 U73 ( .A(n66), .B(n55), .Y(n80) );
  NAND3X1 U74 ( .A(nextState[1]), .B(n36), .C(n61), .Y(n55) );
  NAND3X1 U75 ( .A(n60), .B(n51), .C(RBUF_LOAD), .Y(n66) );
  NAND3X1 U76 ( .A(nextState[0]), .B(n38), .C(n39), .Y(n51) );
  NAND3X1 U77 ( .A(n36), .B(n38), .C(n39), .Y(n60) );
  OAI21X1 U78 ( .A(n40), .B(n43), .C(n67), .Y(n61) );
  NAND3X1 U79 ( .A(state[0]), .B(n43), .C(state[1]), .Y(n67) );
  NAND2X1 U80 ( .A(n68), .B(n69), .Y(n49) );
  OAI21X1 U81 ( .A(n70), .B(n69), .C(n68), .Y(nextState[1]) );
  NOR2X1 U82 ( .A(N99), .B(state[2]), .Y(n70) );
  OAI21X1 U83 ( .A(state[2]), .B(n71), .C(n68), .Y(nextState[0]) );
  NAND2X1 U84 ( .A(state[1]), .B(n44), .Y(n68) );
  AOI21X1 U85 ( .A(START_BIT), .B(n44), .C(n72), .Y(n71) );
  OAI21X1 U86 ( .A(N99), .B(n69), .C(n73), .Y(n72) );
  NAND2X1 U87 ( .A(SB_DETECT), .B(state[1]), .Y(n73) );
  NAND2X1 U88 ( .A(state[0]), .B(n42), .Y(n69) );
  NAND2X1 U89 ( .A(n37), .B(timerRunning), .Y(N31) );
  DFFSR \count_reg[7]  ( .D(nextCount[7]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[7]) );
  DFFSR \count_reg[6]  ( .D(nextCount[6]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[6]) );
  DFFSR \count_reg[5]  ( .D(nextCount[5]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[5]) );
  DFFSR \count_reg[4]  ( .D(nextCount[4]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[4]) );
  DFFSR \count_reg[3]  ( .D(nextCount[3]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[3]) );
  DFFSR \count_reg[2]  ( .D(nextCount[2]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[1]  ( .D(nextCount[1]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[1]) );
  DFFSR \count_reg[0]  ( .D(nextCount[0]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[0]) );
  DFFSR \nextCount_reg[2]  ( .D(N33), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[2]) );
  DFFSR \nextCount_reg[1]  ( .D(N32), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[1]) );
  DFFSR \state_reg[2]  ( .D(n41), .CLK(CLK), .R(n27), .S(1'b1), .Q(state[2])
         );
  DFFSR \nextCount_reg[3]  ( .D(N34), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[3]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        state[1]) );
  DFFSR \nextCount_reg[4]  ( .D(N35), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[4]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        state[0]) );
  DFFSR \nextCount_reg[5]  ( .D(N36), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[5]) );
  DFFSR \nextCount_reg[6]  ( .D(N37), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[6]) );
  DFFSR RBUF_LOAD_reg ( .D(n80), .CLK(CLK), .R(n27), .S(1'b1), .Q(RBUF_LOAD)
         );
  DFFSR timerRunning_reg ( .D(n74), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        timerRunning) );
  DFFSR TIMER_TRIG_reg ( .D(n79), .CLK(CLK), .R(n27), .S(1'b1), .Q(TIMER_TRIG)
         );
  DFFSR SBC_CLR_reg ( .D(n78), .CLK(CLK), .R(n27), .S(1'b1), .Q(SBC_CLR) );
  DFFSR SBC_EN_reg ( .D(n76), .CLK(CLK), .R(n27), .S(1'b1), .Q(SBC_EN) );
  DFFSR \nextCount_reg[7]  ( .D(N38), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[7]) );
  DFFSR SET_RBUF_FULL_reg ( .D(n77), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        SET_RBUF_FULL) );
  DFFSR CHK_ERROR_reg ( .D(n75), .CLK(CLK), .R(n27), .S(1'b1), .Q(CHK_ERROR)
         );
  INVX4 U3 ( .A(RST), .Y(n27) );
  XOR2X1 U30 ( .A(count[7]), .B(\add_46/carry[7] ), .Y(N30) );
  AND2X1 U31 ( .A(count[6]), .B(\add_46/carry[6] ), .Y(\add_46/carry[7] ) );
  XOR2X1 U32 ( .A(\add_46/carry[6] ), .B(count[6]), .Y(N29) );
  AND2X1 U40 ( .A(count[5]), .B(\add_46/carry[5] ), .Y(\add_46/carry[6] ) );
  XOR2X1 U41 ( .A(\add_46/carry[5] ), .B(count[5]), .Y(N28) );
  AND2X1 U42 ( .A(count[4]), .B(\add_46/carry[4] ), .Y(\add_46/carry[5] ) );
  XOR2X1 U43 ( .A(\add_46/carry[4] ), .B(count[4]), .Y(N27) );
  AND2X1 U44 ( .A(count[3]), .B(\add_46/carry[3] ), .Y(\add_46/carry[4] ) );
  XOR2X1 U45 ( .A(\add_46/carry[3] ), .B(count[3]), .Y(N26) );
  AND2X1 U46 ( .A(count[2]), .B(count[1]), .Y(\add_46/carry[3] ) );
  XOR2X1 U47 ( .A(count[1]), .B(count[2]), .Y(N25) );
  INVX2 U48 ( .A(count[1]), .Y(N24) );
  OAI21X1 U49 ( .A(count[0]), .B(count[1]), .C(count[2]), .Y(n28) );
  NOR2X1 U50 ( .A(n33), .B(n28), .Y(n29) );
  OAI21X1 U51 ( .A(n29), .B(count[4]), .C(count[6]), .Y(n30) );
  OAI21X1 U52 ( .A(n32), .B(n30), .C(n31), .Y(N99) );
  INVX2 U53 ( .A(count[7]), .Y(n31) );
  INVX2 U90 ( .A(count[5]), .Y(n32) );
  INVX2 U91 ( .A(count[3]), .Y(n33) );
  INVX2 U92 ( .A(n53), .Y(n34) );
  INVX2 U93 ( .A(n58), .Y(n35) );
  INVX2 U94 ( .A(nextState[0]), .Y(n36) );
  INVX2 U95 ( .A(count[0]), .Y(n37) );
  INVX2 U96 ( .A(nextState[1]), .Y(n38) );
  INVX2 U97 ( .A(n61), .Y(n39) );
  INVX2 U98 ( .A(n49), .Y(n40) );
  INVX2 U99 ( .A(n48), .Y(n41) );
  INVX2 U100 ( .A(state[1]), .Y(n42) );
  INVX2 U101 ( .A(state[2]), .Y(n43) );
  INVX2 U102 ( .A(state[0]), .Y(n44) );
  INVX2 U103 ( .A(SBC_CLR), .Y(n45) );
  INVX2 U104 ( .A(TIMER_TRIG), .Y(n46) );
  INVX2 U105 ( .A(SBC_EN), .Y(n47) );
endmodule


module uart_rcv_buf_1 ( CLK, RST, LOAD_RBUF, LOAD_DATA, RCV_DATA );
  input [7:0] LOAD_DATA;
  output [7:0] RCV_DATA;
  input CLK, RST, LOAD_RBUF;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27;

  AOI22X1 U3 ( .A(n17), .B(LOAD_DATA[0]), .C(RCV_DATA[0]), .D(n27), .Y(n1) );
  AOI22X1 U5 ( .A(LOAD_DATA[1]), .B(n17), .C(RCV_DATA[1]), .D(n27), .Y(n3) );
  AOI22X1 U7 ( .A(LOAD_DATA[2]), .B(n17), .C(RCV_DATA[2]), .D(n27), .Y(n4) );
  AOI22X1 U9 ( .A(LOAD_DATA[3]), .B(n17), .C(RCV_DATA[3]), .D(n27), .Y(n5) );
  AOI22X1 U11 ( .A(LOAD_DATA[4]), .B(n17), .C(RCV_DATA[4]), .D(n27), .Y(n6) );
  AOI22X1 U13 ( .A(LOAD_DATA[5]), .B(n17), .C(RCV_DATA[5]), .D(n27), .Y(n7) );
  AOI22X1 U15 ( .A(LOAD_DATA[6]), .B(n17), .C(RCV_DATA[6]), .D(n27), .Y(n8) );
  AOI22X1 U18 ( .A(LOAD_DATA[7]), .B(n17), .C(RCV_DATA[7]), .D(n27), .Y(n9) );
  DFFSR \Q_int_reg[0]  ( .D(n26), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[0]) );
  DFFSR \Q_int_reg[7]  ( .D(n19), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[7]) );
  DFFSR \Q_int_reg[6]  ( .D(n20), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[6]) );
  DFFSR \Q_int_reg[5]  ( .D(n21), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[5]) );
  DFFSR \Q_int_reg[4]  ( .D(n22), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[4]) );
  DFFSR \Q_int_reg[2]  ( .D(n24), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[2]) );
  DFFSR \Q_int_reg[3]  ( .D(n23), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[3]) );
  DFFSR \Q_int_reg[1]  ( .D(n25), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[1]) );
  INVX2 U17 ( .A(RST), .Y(n18) );
  BUFX2 U19 ( .A(LOAD_RBUF), .Y(n17) );
  INVX2 U20 ( .A(n9), .Y(n19) );
  INVX2 U21 ( .A(n8), .Y(n20) );
  INVX2 U22 ( .A(n7), .Y(n21) );
  INVX2 U23 ( .A(n6), .Y(n22) );
  INVX2 U24 ( .A(n5), .Y(n23) );
  INVX2 U25 ( .A(n4), .Y(n24) );
  INVX2 U26 ( .A(n3), .Y(n25) );
  INVX2 U27 ( .A(n1), .Y(n26) );
  INVX2 U28 ( .A(n17), .Y(n27) );
endmodule


module uart_rcv_buf_full_1 ( CLK, RST, CLR_RBUF, SET_RBUF_FULL, RBUF_FULL );
  input CLK, RST, CLR_RBUF, SET_RBUF_FULL;
  output RBUF_FULL;
  wire   n1, n3;

  NOR2X1 U3 ( .A(RST), .B(CLR_RBUF), .Y(n1) );
  OR2X2 U4 ( .A(RBUF_FULL), .B(SET_RBUF_FULL), .Y(n3) );
  DFFSR Q_int_reg ( .D(n3), .CLK(CLK), .R(n1), .S(1'b1), .Q(RBUF_FULL) );
endmodule


module uart_sb_check_1 ( RST, CLK, SBC_CLR, SBC_EN, STOP_DATA, SB_DETECT, SBE
 );
  input [1:0] STOP_DATA;
  input RST, CLK, SBC_CLR, SBC_EN;
  output SB_DETECT, SBE;
  wire   SBE_prime, sb_detect_flag, n7, n8, n9, n3, n4, n5, n6;

  OR2X2 U6 ( .A(SBC_CLR), .B(STOP_DATA[0]), .Y(n7) );
  NOR2X1 U10 ( .A(n7), .B(n8), .Y(sb_detect_flag) );
  NAND2X1 U11 ( .A(STOP_DATA[1]), .B(SBC_EN), .Y(n8) );
  NOR2X1 U12 ( .A(n6), .B(n9), .Y(SBE_prime) );
  OAI21X1 U13 ( .A(STOP_DATA[0]), .B(n4), .C(n5), .Y(n9) );
  DFFSR SBE_reg ( .D(SBE_prime), .CLK(CLK), .R(n3), .S(1'b1), .Q(SBE) );
  DFFSR SB_DETECT_reg ( .D(sb_detect_flag), .CLK(CLK), .R(n3), .S(1'b1), .Q(
        SB_DETECT) );
  INVX2 U5 ( .A(RST), .Y(n3) );
  INVX2 U7 ( .A(STOP_DATA[1]), .Y(n4) );
  INVX2 U8 ( .A(SBC_CLR), .Y(n5) );
  INVX2 U9 ( .A(SBC_EN), .Y(n6) );
endmodule


module uart_sr_10bit_1 ( CLK, RST, SHIFT_STROBE, SERIAL_IN, LOAD_DATA, 
        STOP_DATA );
  output [7:0] LOAD_DATA;
  output [1:0] STOP_DATA;
  input CLK, RST, SHIFT_STROBE, SERIAL_IN;
  wire   n3, n12, n14, n16, n18, n20, n22, n24, n26, n28, n30, n33, n13, n15,
         n17, n19, n21, n23, n25, n27, n29, n31, n32;

  OAI21X1 U2 ( .A(n32), .B(n13), .C(n3), .Y(n14) );
  NAND2X1 U3 ( .A(LOAD_DATA[0]), .B(n13), .Y(n3) );
  OAI22X1 U4 ( .A(n13), .B(n31), .C(SHIFT_STROBE), .D(n32), .Y(n16) );
  OAI22X1 U6 ( .A(n13), .B(n29), .C(SHIFT_STROBE), .D(n31), .Y(n18) );
  OAI22X1 U8 ( .A(n13), .B(n27), .C(SHIFT_STROBE), .D(n29), .Y(n20) );
  OAI22X1 U10 ( .A(n13), .B(n25), .C(SHIFT_STROBE), .D(n27), .Y(n22) );
  OAI22X1 U12 ( .A(n13), .B(n23), .C(SHIFT_STROBE), .D(n25), .Y(n24) );
  OAI22X1 U14 ( .A(n13), .B(n21), .C(SHIFT_STROBE), .D(n23), .Y(n26) );
  OAI22X1 U16 ( .A(n13), .B(n19), .C(SHIFT_STROBE), .D(n21), .Y(n28) );
  OAI22X1 U18 ( .A(n13), .B(n17), .C(SHIFT_STROBE), .D(n19), .Y(n30) );
  OAI21X1 U22 ( .A(SHIFT_STROBE), .B(n17), .C(n12), .Y(n33) );
  NAND2X1 U23 ( .A(SERIAL_IN), .B(SHIFT_STROBE), .Y(n12) );
  DFFSR \present_val_reg[9]  ( .D(n33), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        STOP_DATA[1]) );
  DFFSR \present_val_reg[8]  ( .D(n30), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        STOP_DATA[0]) );
  DFFSR \present_val_reg[7]  ( .D(n28), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[7]) );
  DFFSR \present_val_reg[6]  ( .D(n26), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[6]) );
  DFFSR \present_val_reg[5]  ( .D(n24), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[5]) );
  DFFSR \present_val_reg[4]  ( .D(n22), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[4]) );
  DFFSR \present_val_reg[3]  ( .D(n20), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[3]) );
  DFFSR \present_val_reg[2]  ( .D(n18), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[2]) );
  DFFSR \present_val_reg[1]  ( .D(n16), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[1]) );
  DFFSR \present_val_reg[0]  ( .D(n14), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[0]) );
  INVX2 U24 ( .A(RST), .Y(n15) );
  INVX2 U25 ( .A(SHIFT_STROBE), .Y(n13) );
  INVX2 U26 ( .A(STOP_DATA[1]), .Y(n17) );
  INVX2 U27 ( .A(STOP_DATA[0]), .Y(n19) );
  INVX2 U28 ( .A(LOAD_DATA[7]), .Y(n21) );
  INVX2 U29 ( .A(LOAD_DATA[6]), .Y(n23) );
  INVX2 U30 ( .A(LOAD_DATA[5]), .Y(n25) );
  INVX2 U31 ( .A(LOAD_DATA[4]), .Y(n27) );
  INVX2 U32 ( .A(LOAD_DATA[3]), .Y(n29) );
  INVX2 U33 ( .A(LOAD_DATA[2]), .Y(n31) );
  INVX2 U34 ( .A(LOAD_DATA[1]), .Y(n32) );
endmodule


module keyreg_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n9), .YC(carry[2]), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(A[3]), .B(B[3]), .Y(n1) );
  XOR2X1 U2 ( .A(n1), .B(carry[3]), .Y(SUM[3]) );
  NAND2X1 U3 ( .A(A[3]), .B(B[3]), .Y(n2) );
  NAND2X1 U4 ( .A(A[3]), .B(carry[3]), .Y(n3) );
  NAND2X1 U5 ( .A(B[3]), .B(carry[3]), .Y(n4) );
  NAND3X1 U6 ( .A(n2), .B(n3), .C(n4), .Y(carry[4]) );
  XOR2X1 U7 ( .A(A[4]), .B(B[4]), .Y(n5) );
  XOR2X1 U8 ( .A(n5), .B(carry[4]), .Y(SUM[4]) );
  NAND2X1 U9 ( .A(A[4]), .B(B[4]), .Y(n6) );
  NAND2X1 U10 ( .A(A[4]), .B(carry[4]), .Y(n7) );
  NAND2X1 U11 ( .A(B[4]), .B(carry[4]), .Y(n8) );
  NAND3X1 U12 ( .A(n6), .B(n7), .C(n8), .Y(carry[5]) );
  AND2X2 U13 ( .A(B[0]), .B(A[0]), .Y(n9) );
  XOR2X1 U14 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module keyreg_1 ( CLK, RST, SBE, OE, RBUF_FULL, RCV_DATA, PLAINKEY, KEY_ERROR, 
        PROG_ERROR, CLR_RBUFF, PARITY_ERROR );
  input [7:0] RCV_DATA;
  output [63:0] PLAINKEY;
  input CLK, RST, SBE, OE, RBUF_FULL;
  output KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR;
  wire   parityError, nextParityError, N694, N1792, N1793, N1794, N1795, N1796,
         N1797, N1798, N1799, n12, n13, n15, n18, n22, n24, n26, n28, n30, n32,
         n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60,
         n62, n64, n66, n68, n70, n72, n74, n76, n78, n80, n82, n84, n86, n88,
         n90, n92, n94, n96, n98, n100, n102, n104, n106, n108, n110, n112,
         n114, n116, n118, n120, n122, n124, n126, n128, n130, n132, n134,
         n136, n138, n140, n142, n144, n146, n148, n152, n155, n157, n159,
         n162, n163, n164, n167, n169, n170, n171, n174, n176, n179, n182,
         n190, n191, n194, n196, n198, n199, n200, n201, n202, n204, n211,
         n212, n213, n214, n215, n216, n218, n220, n235, n236, n237, n238,
         n239, n246, n251, n252, n253, n254, n256, n272, n273, n274, n276,
         n283, n288, n290, n292, n293, n294, n306, n307, n308, n309, n310,
         n318, n323, n325, n328, n329, n341, n342, n349, n354, n356, n358,
         n359, n371, n372, n379, n384, n386, n388, n389, n401, n402, n403,
         n410, n415, n417, n420, n421, n433, n434, n442, n447, n449, n451,
         n463, n464, n470, n475, n477, n478, n490, n491, n497, n502, n504,
         n505, n517, n518, n524, n529, n531, n532, n544, n545, n546, n553,
         n558, n560, n562, n574, n575, n581, n586, n588, n589, n601, n602,
         n608, n613, n615, n616, n628, n629, n635, n640, n642, n643, n655,
         n656, n664, n669, n671, n673, n685, n686, n692, n697, n699, n700,
         n712, n713, n719, n724, n726, n727, n739, n740, n746, n751, n753,
         n754, n766, n767, n768, n775, n780, n782, n784, n796, n797, n803,
         n808, n810, n811, n823, n824, n830, n835, n837, n838, n850, n851,
         n857, n862, n864, n865, n877, n878, n886, n891, n893, n895, n907,
         n908, n914, n919, n921, n922, n934, n935, n941, n946, n948, n949,
         n961, n962, n968, n973, n975, n976, n988, n989, n990, n1002, n1004,
         n1006, n1011, n1018, n1019, n1031, n1033, n1034, n1038, n1046, n1047,
         n1062, n1063, n1077, n1078, n1089, n1090, n1101, n1103, n1104, n1105,
         n1106, n1107, n1108, n1143, n1144, n1160, n1178, n1186, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n14, n16, n17, n19, n20,
         n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47,
         n49, n51, n53, n55, n57, n59, n61, n63, n65, n67, n69, n83, n85, n87,
         n89, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109, n111,
         n113, n115, n117, n119, n121, n123, n125, n127, n129, n131, n133,
         n135, n137, n139, n141, n143, n145, n147, n149, n150, n151, n153,
         n154, n156, n158, n160, n161, n165, n166, n168, n172, n173, n175,
         n177, n178, n180, n181, n183, n184, n185, n186, n187, n188, n189,
         n192, n193, n195, n197, n203, n205, n206, n207, n208, n209, n210,
         n217, n219, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n240, n241, n242, n243, n244, n245,
         n247, n248, n249, n250, n255, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n275, n277,
         n278, n279, n280, n281, n282, n284, n285, n286, n287, n289, n291,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n311, n312, n313, n314, n315, n316, n317, n319, n320, n321, n322,
         n324, n326, n327, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n343, n344, n345, n346, n347, n348, n350, n351,
         n352, n353, n355, n357, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n373, n374, n375, n376, n377, n378, n380,
         n381, n382, n383, n385, n387, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n404, n405, n406, n407, n408, n409,
         n411, n412, n413, n414, n416, n418, n419, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n435, n436, n437, n438,
         n439, n440, n441, n443, n444, n445, n446, n448, n450, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n465, n466,
         n467, n468, n469, n471, n472, n473, n474, n476, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n492, n493, n494,
         n495, n496, n498, n499, n500, n501, n503, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n519, n520, n521, n522,
         n523, n525, n526, n527, n528, n530, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n547, n548, n549, n550, n551,
         n552, n554, n555, n556, n557, n559, n561, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n576, n577, n578, n579,
         n580, n582, n583, n584, n585, n587, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n603, n604, n605, n606, n607,
         n609, n610, n611, n612, n614, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n630, n631, n632, n633, n634, n636,
         n637, n638, n639, n641, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n657, n658, n659, n660, n661, n662, n663,
         n665, n666, n667, n668, n670, n672, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n687, n688, n689, n690, n691,
         n693, n694, n695, n696, n698, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n714, n715, n716, n717, n718, n720,
         n721, n722, n723, n725, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n741, n742, n743, n744, n745, n747, n748,
         n749, n750, n752, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n769, n770, n771, n772, n773, n774, n776, n777,
         n778, n779, n781, n783, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n798, n799, n800, n801, n802, n804, n805,
         n806, n807, n809, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n825, n826, n827, n828, n829, n831, n832, n833,
         n834, n836, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n852, n853, n854, n855, n856, n858, n859, n860, n861,
         n863, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n879, n880, n881, n882, n883, n884, n885, n887, n888, n889,
         n890, n892, n894, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n909, n910, n911, n912, n913, n915, n916, n917,
         n918, n920, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n936, n937, n938, n939, n940, n942, n943, n944, n945,
         n947, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n963, n964, n965, n966, n967, n969, n970, n971, n972, n974,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1003, n1005, n1007, n1008, n1009, n1010, n1012, n1013, n1014, n1015,
         n1016, n1017, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1032, n1035, n1036, n1037, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1102, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579;
  wire   [3:0] state;
  wire   [3:0] keyCount;
  wire   [7:0] address;
  wire   [63:0] currentPlainKey;
  wire   [7:0] parityAccumulator;

  DFFPOSX1 \keyCount_reg[0]  ( .D(n1356), .CLK(CLK), .Q(keyCount[0]) );
  DFFPOSX1 \keyCount_reg[2]  ( .D(n1349), .CLK(CLK), .Q(keyCount[2]) );
  DFFPOSX1 \keyCount_reg[3]  ( .D(n1355), .CLK(CLK), .Q(keyCount[3]) );
  DFFPOSX1 \parityAccumulator_reg[0]  ( .D(n1348), .CLK(CLK), .Q(
        parityAccumulator[0]) );
  DFFPOSX1 \parityAccumulator_reg[1]  ( .D(n1347), .CLK(CLK), .Q(
        parityAccumulator[1]) );
  DFFPOSX1 \parityAccumulator_reg[2]  ( .D(n1346), .CLK(CLK), .Q(
        parityAccumulator[2]) );
  DFFPOSX1 \parityAccumulator_reg[3]  ( .D(n1345), .CLK(CLK), .Q(
        parityAccumulator[3]) );
  DFFPOSX1 \parityAccumulator_reg[4]  ( .D(n1344), .CLK(CLK), .Q(
        parityAccumulator[4]) );
  DFFPOSX1 \parityAccumulator_reg[5]  ( .D(n1343), .CLK(CLK), .Q(
        parityAccumulator[5]) );
  DFFPOSX1 \parityAccumulator_reg[6]  ( .D(n1342), .CLK(CLK), .Q(
        parityAccumulator[6]) );
  DFFPOSX1 \parityAccumulator_reg[7]  ( .D(n1341), .CLK(CLK), .Q(
        parityAccumulator[7]) );
  DFFPOSX1 \keyCount_reg[1]  ( .D(n1350), .CLK(CLK), .Q(keyCount[1]) );
  DFFPOSX1 \address_reg[7]  ( .D(n1340), .CLK(CLK), .Q(address[7]) );
  DFFPOSX1 \address_reg[6]  ( .D(n1339), .CLK(CLK), .Q(address[6]) );
  DFFPOSX1 \address_reg[5]  ( .D(n1338), .CLK(CLK), .Q(address[5]) );
  DFFPOSX1 \address_reg[4]  ( .D(n1337), .CLK(CLK), .Q(address[4]) );
  DFFPOSX1 \address_reg[3]  ( .D(n1336), .CLK(CLK), .Q(address[3]) );
  DFFPOSX1 \address_reg[2]  ( .D(n1335), .CLK(CLK), .Q(address[2]) );
  DFFPOSX1 \address_reg[1]  ( .D(n1334), .CLK(CLK), .Q(address[1]) );
  DFFPOSX1 \address_reg[0]  ( .D(n1333), .CLK(CLK), .Q(address[0]) );
  DFFPOSX1 \currentPlainKey_reg[63]  ( .D(n1269), .CLK(CLK), .Q(
        currentPlainKey[63]) );
  DFFPOSX1 \currentPlainKey_reg[62]  ( .D(n1270), .CLK(CLK), .Q(
        currentPlainKey[62]) );
  DFFPOSX1 \currentPlainKey_reg[61]  ( .D(n1271), .CLK(CLK), .Q(
        currentPlainKey[61]) );
  DFFPOSX1 \currentPlainKey_reg[60]  ( .D(n1272), .CLK(CLK), .Q(
        currentPlainKey[60]) );
  DFFPOSX1 \currentPlainKey_reg[59]  ( .D(n1273), .CLK(CLK), .Q(
        currentPlainKey[59]) );
  DFFPOSX1 \currentPlainKey_reg[58]  ( .D(n1274), .CLK(CLK), .Q(
        currentPlainKey[58]) );
  DFFPOSX1 \currentPlainKey_reg[57]  ( .D(n1275), .CLK(CLK), .Q(
        currentPlainKey[57]) );
  DFFPOSX1 \currentPlainKey_reg[56]  ( .D(n1276), .CLK(CLK), .Q(
        currentPlainKey[56]) );
  DFFPOSX1 \currentPlainKey_reg[55]  ( .D(n1277), .CLK(CLK), .Q(
        currentPlainKey[55]) );
  DFFPOSX1 \currentPlainKey_reg[54]  ( .D(n1278), .CLK(CLK), .Q(
        currentPlainKey[54]) );
  DFFPOSX1 \currentPlainKey_reg[53]  ( .D(n1279), .CLK(CLK), .Q(
        currentPlainKey[53]) );
  DFFPOSX1 \currentPlainKey_reg[52]  ( .D(n1280), .CLK(CLK), .Q(
        currentPlainKey[52]) );
  DFFPOSX1 \currentPlainKey_reg[51]  ( .D(n1281), .CLK(CLK), .Q(
        currentPlainKey[51]) );
  DFFPOSX1 \currentPlainKey_reg[50]  ( .D(n1282), .CLK(CLK), .Q(
        currentPlainKey[50]) );
  DFFPOSX1 \currentPlainKey_reg[49]  ( .D(n1283), .CLK(CLK), .Q(
        currentPlainKey[49]) );
  DFFPOSX1 \currentPlainKey_reg[48]  ( .D(n1284), .CLK(CLK), .Q(
        currentPlainKey[48]) );
  DFFPOSX1 \currentPlainKey_reg[47]  ( .D(n1285), .CLK(CLK), .Q(
        currentPlainKey[47]) );
  DFFPOSX1 \currentPlainKey_reg[46]  ( .D(n1286), .CLK(CLK), .Q(
        currentPlainKey[46]) );
  DFFPOSX1 \currentPlainKey_reg[45]  ( .D(n1287), .CLK(CLK), .Q(
        currentPlainKey[45]) );
  DFFPOSX1 \currentPlainKey_reg[44]  ( .D(n1288), .CLK(CLK), .Q(
        currentPlainKey[44]) );
  DFFPOSX1 \currentPlainKey_reg[43]  ( .D(n1289), .CLK(CLK), .Q(
        currentPlainKey[43]) );
  DFFPOSX1 \currentPlainKey_reg[42]  ( .D(n1290), .CLK(CLK), .Q(
        currentPlainKey[42]) );
  DFFPOSX1 \currentPlainKey_reg[41]  ( .D(n1291), .CLK(CLK), .Q(
        currentPlainKey[41]) );
  DFFPOSX1 \currentPlainKey_reg[40]  ( .D(n1292), .CLK(CLK), .Q(
        currentPlainKey[40]) );
  DFFPOSX1 \currentPlainKey_reg[39]  ( .D(n1293), .CLK(CLK), .Q(
        currentPlainKey[39]) );
  DFFPOSX1 \currentPlainKey_reg[38]  ( .D(n1294), .CLK(CLK), .Q(
        currentPlainKey[38]) );
  DFFPOSX1 \currentPlainKey_reg[37]  ( .D(n1295), .CLK(CLK), .Q(
        currentPlainKey[37]) );
  DFFPOSX1 \currentPlainKey_reg[36]  ( .D(n1296), .CLK(CLK), .Q(
        currentPlainKey[36]) );
  DFFPOSX1 \currentPlainKey_reg[35]  ( .D(n1297), .CLK(CLK), .Q(
        currentPlainKey[35]) );
  DFFPOSX1 \currentPlainKey_reg[34]  ( .D(n1298), .CLK(CLK), .Q(
        currentPlainKey[34]) );
  DFFPOSX1 \currentPlainKey_reg[33]  ( .D(n1299), .CLK(CLK), .Q(
        currentPlainKey[33]) );
  DFFPOSX1 \currentPlainKey_reg[32]  ( .D(n1300), .CLK(CLK), .Q(
        currentPlainKey[32]) );
  DFFPOSX1 \currentPlainKey_reg[31]  ( .D(n1301), .CLK(CLK), .Q(
        currentPlainKey[31]) );
  DFFPOSX1 \currentPlainKey_reg[30]  ( .D(n1302), .CLK(CLK), .Q(
        currentPlainKey[30]) );
  DFFPOSX1 \currentPlainKey_reg[29]  ( .D(n1303), .CLK(CLK), .Q(
        currentPlainKey[29]) );
  DFFPOSX1 \currentPlainKey_reg[28]  ( .D(n1304), .CLK(CLK), .Q(
        currentPlainKey[28]) );
  DFFPOSX1 \currentPlainKey_reg[27]  ( .D(n1305), .CLK(CLK), .Q(
        currentPlainKey[27]) );
  DFFPOSX1 \currentPlainKey_reg[26]  ( .D(n1306), .CLK(CLK), .Q(
        currentPlainKey[26]) );
  DFFPOSX1 \currentPlainKey_reg[25]  ( .D(n1307), .CLK(CLK), .Q(
        currentPlainKey[25]) );
  DFFPOSX1 \currentPlainKey_reg[24]  ( .D(n1308), .CLK(CLK), .Q(
        currentPlainKey[24]) );
  DFFPOSX1 \currentPlainKey_reg[23]  ( .D(n1309), .CLK(CLK), .Q(
        currentPlainKey[23]) );
  DFFPOSX1 \currentPlainKey_reg[22]  ( .D(n1310), .CLK(CLK), .Q(
        currentPlainKey[22]) );
  DFFPOSX1 \currentPlainKey_reg[21]  ( .D(n1311), .CLK(CLK), .Q(
        currentPlainKey[21]) );
  DFFPOSX1 \currentPlainKey_reg[20]  ( .D(n1312), .CLK(CLK), .Q(
        currentPlainKey[20]) );
  DFFPOSX1 \currentPlainKey_reg[19]  ( .D(n1313), .CLK(CLK), .Q(
        currentPlainKey[19]) );
  DFFPOSX1 \currentPlainKey_reg[18]  ( .D(n1314), .CLK(CLK), .Q(
        currentPlainKey[18]) );
  DFFPOSX1 \currentPlainKey_reg[17]  ( .D(n1315), .CLK(CLK), .Q(
        currentPlainKey[17]) );
  DFFPOSX1 \currentPlainKey_reg[16]  ( .D(n1316), .CLK(CLK), .Q(
        currentPlainKey[16]) );
  DFFPOSX1 \currentPlainKey_reg[15]  ( .D(n1317), .CLK(CLK), .Q(
        currentPlainKey[15]) );
  DFFPOSX1 \currentPlainKey_reg[14]  ( .D(n1318), .CLK(CLK), .Q(
        currentPlainKey[14]) );
  DFFPOSX1 \currentPlainKey_reg[13]  ( .D(n1319), .CLK(CLK), .Q(
        currentPlainKey[13]) );
  DFFPOSX1 \currentPlainKey_reg[12]  ( .D(n1320), .CLK(CLK), .Q(
        currentPlainKey[12]) );
  DFFPOSX1 \currentPlainKey_reg[11]  ( .D(n1321), .CLK(CLK), .Q(
        currentPlainKey[11]) );
  DFFPOSX1 \currentPlainKey_reg[10]  ( .D(n1322), .CLK(CLK), .Q(
        currentPlainKey[10]) );
  DFFPOSX1 \currentPlainKey_reg[9]  ( .D(n1323), .CLK(CLK), .Q(
        currentPlainKey[9]) );
  DFFPOSX1 \currentPlainKey_reg[8]  ( .D(n1324), .CLK(CLK), .Q(
        currentPlainKey[8]) );
  DFFPOSX1 \currentPlainKey_reg[7]  ( .D(n1325), .CLK(CLK), .Q(
        currentPlainKey[7]) );
  DFFPOSX1 \currentPlainKey_reg[6]  ( .D(n1326), .CLK(CLK), .Q(
        currentPlainKey[6]) );
  DFFPOSX1 \currentPlainKey_reg[5]  ( .D(n1327), .CLK(CLK), .Q(
        currentPlainKey[5]) );
  DFFPOSX1 \currentPlainKey_reg[4]  ( .D(n1328), .CLK(CLK), .Q(
        currentPlainKey[4]) );
  DFFPOSX1 \currentPlainKey_reg[3]  ( .D(n1329), .CLK(CLK), .Q(
        currentPlainKey[3]) );
  DFFPOSX1 \currentPlainKey_reg[2]  ( .D(n1330), .CLK(CLK), .Q(
        currentPlainKey[2]) );
  DFFPOSX1 \currentPlainKey_reg[1]  ( .D(n1331), .CLK(CLK), .Q(
        currentPlainKey[1]) );
  DFFPOSX1 \currentPlainKey_reg[0]  ( .D(n1332), .CLK(CLK), .Q(
        currentPlainKey[0]) );
  DFFPOSX1 \PLAINKEY_reg[63]  ( .D(n1260), .CLK(CLK), .Q(PLAINKEY[63]) );
  DFFPOSX1 \PLAINKEY_reg[62]  ( .D(n1259), .CLK(CLK), .Q(PLAINKEY[62]) );
  DFFPOSX1 \PLAINKEY_reg[61]  ( .D(n1258), .CLK(CLK), .Q(PLAINKEY[61]) );
  DFFPOSX1 \PLAINKEY_reg[60]  ( .D(n1257), .CLK(CLK), .Q(PLAINKEY[60]) );
  DFFPOSX1 \PLAINKEY_reg[59]  ( .D(n1256), .CLK(CLK), .Q(PLAINKEY[59]) );
  DFFPOSX1 \PLAINKEY_reg[58]  ( .D(n1255), .CLK(CLK), .Q(PLAINKEY[58]) );
  DFFPOSX1 \PLAINKEY_reg[57]  ( .D(n1254), .CLK(CLK), .Q(PLAINKEY[57]) );
  DFFPOSX1 \PLAINKEY_reg[56]  ( .D(n1253), .CLK(CLK), .Q(PLAINKEY[56]) );
  DFFPOSX1 \PLAINKEY_reg[55]  ( .D(n1252), .CLK(CLK), .Q(PLAINKEY[55]) );
  DFFPOSX1 \PLAINKEY_reg[54]  ( .D(n1251), .CLK(CLK), .Q(PLAINKEY[54]) );
  DFFPOSX1 \PLAINKEY_reg[53]  ( .D(n1250), .CLK(CLK), .Q(PLAINKEY[53]) );
  DFFPOSX1 \PLAINKEY_reg[52]  ( .D(n1249), .CLK(CLK), .Q(PLAINKEY[52]) );
  DFFPOSX1 \PLAINKEY_reg[51]  ( .D(n1248), .CLK(CLK), .Q(PLAINKEY[51]) );
  DFFPOSX1 \PLAINKEY_reg[50]  ( .D(n1247), .CLK(CLK), .Q(PLAINKEY[50]) );
  DFFPOSX1 \PLAINKEY_reg[49]  ( .D(n1246), .CLK(CLK), .Q(PLAINKEY[49]) );
  DFFPOSX1 \PLAINKEY_reg[48]  ( .D(n1245), .CLK(CLK), .Q(PLAINKEY[48]) );
  DFFPOSX1 \PLAINKEY_reg[47]  ( .D(n1244), .CLK(CLK), .Q(PLAINKEY[47]) );
  DFFPOSX1 \PLAINKEY_reg[46]  ( .D(n1243), .CLK(CLK), .Q(PLAINKEY[46]) );
  DFFPOSX1 \PLAINKEY_reg[45]  ( .D(n1242), .CLK(CLK), .Q(PLAINKEY[45]) );
  DFFPOSX1 \PLAINKEY_reg[44]  ( .D(n1241), .CLK(CLK), .Q(PLAINKEY[44]) );
  DFFPOSX1 \PLAINKEY_reg[43]  ( .D(n1240), .CLK(CLK), .Q(PLAINKEY[43]) );
  DFFPOSX1 \PLAINKEY_reg[42]  ( .D(n1239), .CLK(CLK), .Q(PLAINKEY[42]) );
  DFFPOSX1 \PLAINKEY_reg[41]  ( .D(n1238), .CLK(CLK), .Q(PLAINKEY[41]) );
  DFFPOSX1 \PLAINKEY_reg[40]  ( .D(n1237), .CLK(CLK), .Q(PLAINKEY[40]) );
  DFFPOSX1 \PLAINKEY_reg[39]  ( .D(n1236), .CLK(CLK), .Q(PLAINKEY[39]) );
  DFFPOSX1 \PLAINKEY_reg[38]  ( .D(n1235), .CLK(CLK), .Q(PLAINKEY[38]) );
  DFFPOSX1 \PLAINKEY_reg[37]  ( .D(n1234), .CLK(CLK), .Q(PLAINKEY[37]) );
  DFFPOSX1 \PLAINKEY_reg[36]  ( .D(n1233), .CLK(CLK), .Q(PLAINKEY[36]) );
  DFFPOSX1 \PLAINKEY_reg[35]  ( .D(n1232), .CLK(CLK), .Q(PLAINKEY[35]) );
  DFFPOSX1 \PLAINKEY_reg[34]  ( .D(n1231), .CLK(CLK), .Q(PLAINKEY[34]) );
  DFFPOSX1 \PLAINKEY_reg[33]  ( .D(n1230), .CLK(CLK), .Q(PLAINKEY[33]) );
  DFFPOSX1 \PLAINKEY_reg[32]  ( .D(n1229), .CLK(CLK), .Q(PLAINKEY[32]) );
  DFFPOSX1 \PLAINKEY_reg[31]  ( .D(n1228), .CLK(CLK), .Q(PLAINKEY[31]) );
  DFFPOSX1 \PLAINKEY_reg[30]  ( .D(n1227), .CLK(CLK), .Q(PLAINKEY[30]) );
  DFFPOSX1 \PLAINKEY_reg[29]  ( .D(n1226), .CLK(CLK), .Q(PLAINKEY[29]) );
  DFFPOSX1 \PLAINKEY_reg[28]  ( .D(n1225), .CLK(CLK), .Q(PLAINKEY[28]) );
  DFFPOSX1 \PLAINKEY_reg[27]  ( .D(n1224), .CLK(CLK), .Q(PLAINKEY[27]) );
  DFFPOSX1 \PLAINKEY_reg[26]  ( .D(n1223), .CLK(CLK), .Q(PLAINKEY[26]) );
  DFFPOSX1 \PLAINKEY_reg[25]  ( .D(n1222), .CLK(CLK), .Q(PLAINKEY[25]) );
  DFFPOSX1 \PLAINKEY_reg[24]  ( .D(n1221), .CLK(CLK), .Q(PLAINKEY[24]) );
  DFFPOSX1 \PLAINKEY_reg[23]  ( .D(n1220), .CLK(CLK), .Q(PLAINKEY[23]) );
  DFFPOSX1 \PLAINKEY_reg[22]  ( .D(n1219), .CLK(CLK), .Q(PLAINKEY[22]) );
  DFFPOSX1 \PLAINKEY_reg[21]  ( .D(n1218), .CLK(CLK), .Q(PLAINKEY[21]) );
  DFFPOSX1 \PLAINKEY_reg[20]  ( .D(n1217), .CLK(CLK), .Q(PLAINKEY[20]) );
  DFFPOSX1 \PLAINKEY_reg[19]  ( .D(n1216), .CLK(CLK), .Q(PLAINKEY[19]) );
  DFFPOSX1 \PLAINKEY_reg[18]  ( .D(n1215), .CLK(CLK), .Q(PLAINKEY[18]) );
  DFFPOSX1 \PLAINKEY_reg[17]  ( .D(n1214), .CLK(CLK), .Q(PLAINKEY[17]) );
  DFFPOSX1 \PLAINKEY_reg[16]  ( .D(n1213), .CLK(CLK), .Q(PLAINKEY[16]) );
  DFFPOSX1 \PLAINKEY_reg[15]  ( .D(n1212), .CLK(CLK), .Q(PLAINKEY[15]) );
  DFFPOSX1 \PLAINKEY_reg[14]  ( .D(n1211), .CLK(CLK), .Q(PLAINKEY[14]) );
  DFFPOSX1 \PLAINKEY_reg[13]  ( .D(n1210), .CLK(CLK), .Q(PLAINKEY[13]) );
  DFFPOSX1 \PLAINKEY_reg[12]  ( .D(n1209), .CLK(CLK), .Q(PLAINKEY[12]) );
  DFFPOSX1 \PLAINKEY_reg[11]  ( .D(n1208), .CLK(CLK), .Q(PLAINKEY[11]) );
  DFFPOSX1 \PLAINKEY_reg[10]  ( .D(n1207), .CLK(CLK), .Q(PLAINKEY[10]) );
  DFFPOSX1 \PLAINKEY_reg[9]  ( .D(n1206), .CLK(CLK), .Q(PLAINKEY[9]) );
  DFFPOSX1 \PLAINKEY_reg[8]  ( .D(n1205), .CLK(CLK), .Q(PLAINKEY[8]) );
  DFFPOSX1 \PLAINKEY_reg[7]  ( .D(n1204), .CLK(CLK), .Q(PLAINKEY[7]) );
  DFFPOSX1 \PLAINKEY_reg[6]  ( .D(n1203), .CLK(CLK), .Q(PLAINKEY[6]) );
  DFFPOSX1 \PLAINKEY_reg[5]  ( .D(n1202), .CLK(CLK), .Q(PLAINKEY[5]) );
  DFFPOSX1 \PLAINKEY_reg[4]  ( .D(n1201), .CLK(CLK), .Q(PLAINKEY[4]) );
  DFFPOSX1 \PLAINKEY_reg[3]  ( .D(n1200), .CLK(CLK), .Q(PLAINKEY[3]) );
  DFFPOSX1 \PLAINKEY_reg[2]  ( .D(n1199), .CLK(CLK), .Q(PLAINKEY[2]) );
  DFFPOSX1 \PLAINKEY_reg[1]  ( .D(n1198), .CLK(CLK), .Q(PLAINKEY[1]) );
  DFFPOSX1 \PLAINKEY_reg[0]  ( .D(n1197), .CLK(CLK), .Q(PLAINKEY[0]) );
  NAND3X1 U9 ( .A(parityAccumulator[7]), .B(parityAccumulator[6]), .C(n15), 
        .Y(n13) );
  NOR2X1 U10 ( .A(n1490), .B(n1491), .Y(n15) );
  NAND3X1 U11 ( .A(parityAccumulator[3]), .B(parityAccumulator[2]), .C(n18), 
        .Y(n12) );
  NOR2X1 U12 ( .A(n1486), .B(n1487), .Y(n18) );
  OAI21X1 U13 ( .A(n227), .B(n1573), .C(n22), .Y(n1197) );
  NAND2X1 U14 ( .A(PLAINKEY[0]), .B(n231), .Y(n22) );
  OAI21X1 U15 ( .A(n227), .B(n1572), .C(n24), .Y(n1198) );
  NAND2X1 U16 ( .A(PLAINKEY[1]), .B(RST), .Y(n24) );
  OAI21X1 U17 ( .A(n227), .B(n1571), .C(n26), .Y(n1199) );
  NAND2X1 U18 ( .A(PLAINKEY[2]), .B(RST), .Y(n26) );
  OAI21X1 U19 ( .A(n227), .B(n1570), .C(n28), .Y(n1200) );
  NAND2X1 U20 ( .A(PLAINKEY[3]), .B(RST), .Y(n28) );
  OAI21X1 U21 ( .A(n227), .B(n1569), .C(n30), .Y(n1201) );
  NAND2X1 U22 ( .A(PLAINKEY[4]), .B(n231), .Y(n30) );
  OAI21X1 U24 ( .A(n227), .B(n1568), .C(n32), .Y(n1202) );
  NAND2X1 U25 ( .A(PLAINKEY[5]), .B(n232), .Y(n32) );
  OAI21X1 U27 ( .A(n227), .B(n1567), .C(n34), .Y(n1203) );
  NAND2X1 U28 ( .A(PLAINKEY[6]), .B(n233), .Y(n34) );
  OAI21X1 U30 ( .A(n227), .B(n1566), .C(n36), .Y(n1204) );
  NAND2X1 U31 ( .A(PLAINKEY[7]), .B(RST), .Y(n36) );
  OAI21X1 U33 ( .A(n227), .B(n1565), .C(n38), .Y(n1205) );
  NAND2X1 U34 ( .A(PLAINKEY[8]), .B(n231), .Y(n38) );
  OAI21X1 U36 ( .A(n228), .B(n1564), .C(n40), .Y(n1206) );
  NAND2X1 U37 ( .A(PLAINKEY[9]), .B(n232), .Y(n40) );
  OAI21X1 U39 ( .A(n228), .B(n1563), .C(n42), .Y(n1207) );
  NAND2X1 U40 ( .A(PLAINKEY[10]), .B(n233), .Y(n42) );
  OAI21X1 U42 ( .A(n228), .B(n1562), .C(n44), .Y(n1208) );
  NAND2X1 U43 ( .A(PLAINKEY[11]), .B(n233), .Y(n44) );
  OAI21X1 U45 ( .A(n228), .B(n1561), .C(n46), .Y(n1209) );
  NAND2X1 U46 ( .A(PLAINKEY[12]), .B(n233), .Y(n46) );
  OAI21X1 U48 ( .A(n228), .B(n1560), .C(n48), .Y(n1210) );
  NAND2X1 U49 ( .A(PLAINKEY[13]), .B(n233), .Y(n48) );
  OAI21X1 U51 ( .A(n228), .B(n1559), .C(n50), .Y(n1211) );
  NAND2X1 U52 ( .A(PLAINKEY[14]), .B(n233), .Y(n50) );
  OAI21X1 U54 ( .A(n228), .B(n1558), .C(n52), .Y(n1212) );
  NAND2X1 U55 ( .A(PLAINKEY[15]), .B(n233), .Y(n52) );
  OAI21X1 U57 ( .A(n229), .B(n1557), .C(n54), .Y(n1213) );
  NAND2X1 U58 ( .A(PLAINKEY[16]), .B(n233), .Y(n54) );
  OAI21X1 U60 ( .A(n229), .B(n1556), .C(n56), .Y(n1214) );
  NAND2X1 U61 ( .A(PLAINKEY[17]), .B(n233), .Y(n56) );
  OAI21X1 U63 ( .A(n229), .B(n1555), .C(n58), .Y(n1215) );
  NAND2X1 U64 ( .A(PLAINKEY[18]), .B(n233), .Y(n58) );
  OAI21X1 U66 ( .A(n229), .B(n1554), .C(n60), .Y(n1216) );
  NAND2X1 U67 ( .A(PLAINKEY[19]), .B(n233), .Y(n60) );
  OAI21X1 U69 ( .A(n229), .B(n1553), .C(n62), .Y(n1217) );
  NAND2X1 U70 ( .A(PLAINKEY[20]), .B(n233), .Y(n62) );
  OAI21X1 U72 ( .A(n229), .B(n1552), .C(n64), .Y(n1218) );
  NAND2X1 U73 ( .A(PLAINKEY[21]), .B(n233), .Y(n64) );
  OAI21X1 U75 ( .A(n229), .B(n1551), .C(n66), .Y(n1219) );
  NAND2X1 U76 ( .A(PLAINKEY[22]), .B(n233), .Y(n66) );
  OAI21X1 U78 ( .A(n230), .B(n1550), .C(n68), .Y(n1220) );
  NAND2X1 U79 ( .A(PLAINKEY[23]), .B(n233), .Y(n68) );
  OAI21X1 U81 ( .A(n229), .B(n1549), .C(n70), .Y(n1221) );
  NAND2X1 U82 ( .A(PLAINKEY[24]), .B(n233), .Y(n70) );
  OAI21X1 U84 ( .A(n228), .B(n1548), .C(n72), .Y(n1222) );
  NAND2X1 U85 ( .A(PLAINKEY[25]), .B(n233), .Y(n72) );
  OAI21X1 U87 ( .A(n230), .B(n1547), .C(n74), .Y(n1223) );
  NAND2X1 U88 ( .A(PLAINKEY[26]), .B(n233), .Y(n74) );
  OAI21X1 U90 ( .A(n230), .B(n1546), .C(n76), .Y(n1224) );
  NAND2X1 U91 ( .A(PLAINKEY[27]), .B(n233), .Y(n76) );
  OAI21X1 U93 ( .A(n229), .B(n1545), .C(n78), .Y(n1225) );
  NAND2X1 U94 ( .A(PLAINKEY[28]), .B(n233), .Y(n78) );
  OAI21X1 U96 ( .A(n230), .B(n1544), .C(n80), .Y(n1226) );
  NAND2X1 U97 ( .A(PLAINKEY[29]), .B(n232), .Y(n80) );
  OAI21X1 U99 ( .A(n230), .B(n1543), .C(n82), .Y(n1227) );
  NAND2X1 U100 ( .A(PLAINKEY[30]), .B(n232), .Y(n82) );
  OAI21X1 U102 ( .A(n229), .B(n1542), .C(n84), .Y(n1228) );
  NAND2X1 U103 ( .A(PLAINKEY[31]), .B(n232), .Y(n84) );
  OAI21X1 U105 ( .A(RST), .B(n1541), .C(n86), .Y(n1229) );
  NAND2X1 U106 ( .A(PLAINKEY[32]), .B(n232), .Y(n86) );
  OAI21X1 U108 ( .A(n230), .B(n1540), .C(n88), .Y(n1230) );
  NAND2X1 U109 ( .A(PLAINKEY[33]), .B(n232), .Y(n88) );
  OAI21X1 U111 ( .A(n233), .B(n1539), .C(n90), .Y(n1231) );
  NAND2X1 U112 ( .A(PLAINKEY[34]), .B(n232), .Y(n90) );
  OAI21X1 U114 ( .A(n230), .B(n1538), .C(n92), .Y(n1232) );
  NAND2X1 U115 ( .A(PLAINKEY[35]), .B(n232), .Y(n92) );
  OAI21X1 U117 ( .A(n230), .B(n1537), .C(n94), .Y(n1233) );
  NAND2X1 U118 ( .A(PLAINKEY[36]), .B(n232), .Y(n94) );
  OAI21X1 U120 ( .A(n231), .B(n1536), .C(n96), .Y(n1234) );
  NAND2X1 U121 ( .A(PLAINKEY[37]), .B(n232), .Y(n96) );
  OAI21X1 U123 ( .A(n227), .B(n1535), .C(n98), .Y(n1235) );
  NAND2X1 U124 ( .A(PLAINKEY[38]), .B(n232), .Y(n98) );
  OAI21X1 U126 ( .A(n230), .B(n1534), .C(n100), .Y(n1236) );
  NAND2X1 U127 ( .A(PLAINKEY[39]), .B(n232), .Y(n100) );
  OAI21X1 U129 ( .A(n229), .B(n1533), .C(n102), .Y(n1237) );
  NAND2X1 U130 ( .A(PLAINKEY[40]), .B(n232), .Y(n102) );
  OAI21X1 U132 ( .A(n230), .B(n1532), .C(n104), .Y(n1238) );
  NAND2X1 U133 ( .A(PLAINKEY[41]), .B(n232), .Y(n104) );
  OAI21X1 U135 ( .A(n230), .B(n1531), .C(n106), .Y(n1239) );
  NAND2X1 U136 ( .A(PLAINKEY[42]), .B(n232), .Y(n106) );
  OAI21X1 U138 ( .A(RST), .B(n1530), .C(n108), .Y(n1240) );
  NAND2X1 U139 ( .A(PLAINKEY[43]), .B(n232), .Y(n108) );
  OAI21X1 U141 ( .A(n228), .B(n1529), .C(n110), .Y(n1241) );
  NAND2X1 U142 ( .A(PLAINKEY[44]), .B(n231), .Y(n110) );
  OAI21X1 U144 ( .A(n228), .B(n1528), .C(n112), .Y(n1242) );
  NAND2X1 U145 ( .A(PLAINKEY[45]), .B(n231), .Y(n112) );
  OAI21X1 U147 ( .A(n232), .B(n1527), .C(n114), .Y(n1243) );
  NAND2X1 U148 ( .A(PLAINKEY[46]), .B(n232), .Y(n114) );
  OAI21X1 U150 ( .A(n228), .B(n1526), .C(n116), .Y(n1244) );
  NAND2X1 U151 ( .A(PLAINKEY[47]), .B(n231), .Y(n116) );
  OAI21X1 U153 ( .A(n230), .B(n1525), .C(n118), .Y(n1245) );
  NAND2X1 U154 ( .A(PLAINKEY[48]), .B(n231), .Y(n118) );
  OAI21X1 U156 ( .A(n230), .B(n1524), .C(n120), .Y(n1246) );
  NAND2X1 U157 ( .A(PLAINKEY[49]), .B(n231), .Y(n120) );
  OAI21X1 U159 ( .A(n230), .B(n1523), .C(n122), .Y(n1247) );
  NAND2X1 U160 ( .A(PLAINKEY[50]), .B(n231), .Y(n122) );
  OAI21X1 U162 ( .A(n229), .B(n1522), .C(n124), .Y(n1248) );
  NAND2X1 U163 ( .A(PLAINKEY[51]), .B(n231), .Y(n124) );
  OAI21X1 U165 ( .A(n230), .B(n1521), .C(n126), .Y(n1249) );
  NAND2X1 U166 ( .A(PLAINKEY[52]), .B(n231), .Y(n126) );
  OAI21X1 U168 ( .A(n229), .B(n1520), .C(n128), .Y(n1250) );
  NAND2X1 U169 ( .A(PLAINKEY[53]), .B(n231), .Y(n128) );
  OAI21X1 U171 ( .A(n229), .B(n1519), .C(n130), .Y(n1251) );
  NAND2X1 U172 ( .A(PLAINKEY[54]), .B(n231), .Y(n130) );
  OAI21X1 U174 ( .A(n228), .B(n1518), .C(n132), .Y(n1252) );
  NAND2X1 U175 ( .A(PLAINKEY[55]), .B(n232), .Y(n132) );
  OAI21X1 U177 ( .A(n229), .B(n1517), .C(n134), .Y(n1253) );
  NAND2X1 U178 ( .A(PLAINKEY[56]), .B(n231), .Y(n134) );
  OAI21X1 U180 ( .A(n228), .B(n1516), .C(n136), .Y(n1254) );
  NAND2X1 U181 ( .A(PLAINKEY[57]), .B(n231), .Y(n136) );
  OAI21X1 U183 ( .A(n228), .B(n1515), .C(n138), .Y(n1255) );
  NAND2X1 U184 ( .A(PLAINKEY[58]), .B(n231), .Y(n138) );
  OAI21X1 U186 ( .A(n228), .B(n1514), .C(n140), .Y(n1256) );
  NAND2X1 U187 ( .A(PLAINKEY[59]), .B(n231), .Y(n140) );
  OAI21X1 U188 ( .A(n227), .B(n1513), .C(n142), .Y(n1257) );
  NAND2X1 U189 ( .A(PLAINKEY[60]), .B(n231), .Y(n142) );
  OAI21X1 U191 ( .A(n227), .B(n1512), .C(n144), .Y(n1258) );
  NAND2X1 U192 ( .A(PLAINKEY[61]), .B(n231), .Y(n144) );
  OAI21X1 U194 ( .A(n227), .B(n1511), .C(n146), .Y(n1259) );
  NAND2X1 U195 ( .A(PLAINKEY[62]), .B(n231), .Y(n146) );
  OAI21X1 U196 ( .A(n227), .B(n1510), .C(n148), .Y(n1260) );
  NAND2X1 U197 ( .A(PLAINKEY[63]), .B(n232), .Y(n148) );
  OAI21X1 U202 ( .A(n1449), .B(n162), .C(n157), .Y(n155) );
  AOI22X1 U203 ( .A(n163), .B(n164), .C(n1498), .D(n1576), .Y(n162) );
  OAI22X1 U205 ( .A(RCV_DATA[3]), .B(n167), .C(n1499), .D(n169), .Y(n163) );
  AOI22X1 U206 ( .A(n170), .B(n171), .C(n1500), .D(n1578), .Y(n169) );
  OAI22X1 U208 ( .A(n174), .B(n1501), .C(RCV_DATA[1]), .D(n176), .Y(n170) );
  NAND2X1 U210 ( .A(n33), .B(n14), .Y(n176) );
  AOI22X1 U211 ( .A(n179), .B(n156), .C(n1507), .D(n1510), .Y(n174) );
  NOR2X1 U213 ( .A(n182), .B(n149), .Y(n179) );
  OAI22X1 U220 ( .A(n157), .B(n1575), .C(n159), .D(n1576), .Y(n191) );
  OAI21X1 U221 ( .A(n164), .B(n1577), .C(n194), .Y(n190) );
  AOI22X1 U222 ( .A(RCV_DATA[2]), .B(n1499), .C(n1496), .D(n196), .Y(n194) );
  OAI21X1 U223 ( .A(n171), .B(n226), .C(n198), .Y(n196) );
  NAND2X1 U224 ( .A(n199), .B(n171), .Y(n198) );
  OAI21X1 U225 ( .A(n182), .B(n200), .C(n201), .Y(n199) );
  OAI21X1 U226 ( .A(n202), .B(n182), .C(currentPlainKey[62]), .Y(n201) );
  NAND2X1 U227 ( .A(n31), .B(n14), .Y(n171) );
  OAI21X1 U233 ( .A(n212), .B(n213), .C(n152), .Y(n211) );
  OAI22X1 U234 ( .A(n157), .B(n1576), .C(n164), .D(n1578), .Y(n213) );
  OAI21X1 U235 ( .A(n214), .B(n204), .C(n215), .Y(n212) );
  AOI22X1 U236 ( .A(n225), .B(n1499), .C(RCV_DATA[3]), .D(n1449), .Y(n215) );
  NAND2X1 U238 ( .A(n216), .B(n167), .Y(n204) );
  NAND2X1 U239 ( .A(n29), .B(n14), .Y(n167) );
  AOI22X1 U240 ( .A(n218), .B(n158), .C(currentPlainKey[61]), .D(n1506), .Y(
        n214) );
  NOR2X1 U242 ( .A(n182), .B(n220), .Y(n218) );
  OAI21X1 U252 ( .A(n182), .B(n236), .C(n237), .Y(n235) );
  OAI21X1 U253 ( .A(n238), .B(n182), .C(currentPlainKey[60]), .Y(n237) );
  OAI21X1 U264 ( .A(n157), .B(n1578), .C(n252), .Y(n251) );
  AOI22X1 U265 ( .A(n239), .B(n253), .C(n225), .D(n1449), .Y(n252) );
  OAI22X1 U266 ( .A(n254), .B(n1514), .C(n156), .D(n1505), .Y(n253) );
  NOR2X1 U270 ( .A(n182), .B(n256), .Y(n254) );
  NOR2X1 U271 ( .A(n1449), .B(n1497), .Y(n239) );
  OAI22X1 U284 ( .A(n157), .B(n226), .C(n1497), .D(n273), .Y(n272) );
  AOI22X1 U285 ( .A(n274), .B(n158), .C(currentPlainKey[58]), .D(n1504), .Y(
        n273) );
  NOR2X1 U287 ( .A(n182), .B(n276), .Y(n274) );
  AOI22X1 U300 ( .A(n290), .B(n152), .C(n225), .D(n1450), .Y(n288) );
  OAI21X1 U303 ( .A(n182), .B(n292), .C(n293), .Y(n290) );
  OAI21X1 U304 ( .A(n294), .B(n182), .C(currentPlainKey[57]), .Y(n293) );
  OAI21X1 U314 ( .A(n182), .B(n307), .C(n308), .Y(n306) );
  OAI21X1 U315 ( .A(n309), .B(n182), .C(currentPlainKey[56]), .Y(n308) );
  NAND2X1 U316 ( .A(address[3]), .B(n310), .Y(n182) );
  AOI22X1 U330 ( .A(n325), .B(n246), .C(n1451), .D(n225), .Y(n323) );
  OAI21X1 U333 ( .A(n173), .B(n328), .C(n329), .Y(n325) );
  OAI21X1 U334 ( .A(n149), .B(n173), .C(currentPlainKey[55]), .Y(n329) );
  OAI21X1 U344 ( .A(n200), .B(n173), .C(n342), .Y(n341) );
  OAI21X1 U345 ( .A(n202), .B(n173), .C(currentPlainKey[54]), .Y(n342) );
  AOI22X1 U359 ( .A(n356), .B(n283), .C(n1452), .D(RCV_DATA[1]), .Y(n354) );
  OAI21X1 U362 ( .A(n173), .B(n358), .C(n359), .Y(n356) );
  OAI21X1 U363 ( .A(n220), .B(n173), .C(currentPlainKey[53]), .Y(n359) );
  OAI21X1 U373 ( .A(n236), .B(n173), .C(n372), .Y(n371) );
  OAI21X1 U374 ( .A(n238), .B(n173), .C(currentPlainKey[52]), .Y(n372) );
  AOI22X1 U388 ( .A(n386), .B(n318), .C(n1453), .D(n225), .Y(n384) );
  OAI21X1 U391 ( .A(n173), .B(n388), .C(n389), .Y(n386) );
  OAI21X1 U392 ( .A(n256), .B(n173), .C(currentPlainKey[51]), .Y(n389) );
  OAI21X1 U402 ( .A(n173), .B(n402), .C(n403), .Y(n401) );
  OAI21X1 U403 ( .A(n276), .B(n173), .C(currentPlainKey[50]), .Y(n403) );
  AOI22X1 U417 ( .A(n417), .B(n349), .C(n1454), .D(RCV_DATA[1]), .Y(n415) );
  OAI21X1 U422 ( .A(n292), .B(n173), .C(n421), .Y(n417) );
  OAI21X1 U423 ( .A(n294), .B(n173), .C(currentPlainKey[49]), .Y(n421) );
  OAI21X1 U433 ( .A(n307), .B(n173), .C(n434), .Y(n433) );
  OAI21X1 U434 ( .A(n309), .B(n173), .C(currentPlainKey[48]), .Y(n434) );
  AOI22X1 U449 ( .A(n449), .B(n379), .C(n1455), .D(n225), .Y(n447) );
  OAI21X1 U452 ( .A(n328), .B(n172), .C(n451), .Y(n449) );
  OAI21X1 U453 ( .A(n149), .B(n172), .C(currentPlainKey[47]), .Y(n451) );
  OAI21X1 U463 ( .A(n200), .B(n172), .C(n464), .Y(n463) );
  OAI21X1 U464 ( .A(n202), .B(n172), .C(currentPlainKey[46]), .Y(n464) );
  AOI22X1 U478 ( .A(n477), .B(n410), .C(n1456), .D(RCV_DATA[1]), .Y(n475) );
  OAI21X1 U481 ( .A(n358), .B(n172), .C(n478), .Y(n477) );
  OAI21X1 U482 ( .A(n220), .B(n172), .C(currentPlainKey[45]), .Y(n478) );
  OAI21X1 U492 ( .A(n236), .B(n172), .C(n491), .Y(n490) );
  OAI21X1 U493 ( .A(n238), .B(n172), .C(currentPlainKey[44]), .Y(n491) );
  AOI22X1 U507 ( .A(n504), .B(n442), .C(n1457), .D(n225), .Y(n502) );
  OAI21X1 U510 ( .A(n388), .B(n172), .C(n505), .Y(n504) );
  OAI21X1 U511 ( .A(n256), .B(n172), .C(currentPlainKey[43]), .Y(n505) );
  OAI21X1 U521 ( .A(n402), .B(n172), .C(n518), .Y(n517) );
  OAI21X1 U522 ( .A(n276), .B(n172), .C(currentPlainKey[42]), .Y(n518) );
  AOI22X1 U536 ( .A(n531), .B(n470), .C(n1458), .D(n225), .Y(n529) );
  OAI21X1 U539 ( .A(n292), .B(n172), .C(n532), .Y(n531) );
  OAI21X1 U540 ( .A(n294), .B(n172), .C(currentPlainKey[41]), .Y(n532) );
  OAI21X1 U550 ( .A(n307), .B(n172), .C(n545), .Y(n544) );
  OAI21X1 U551 ( .A(n309), .B(n172), .C(currentPlainKey[40]), .Y(n545) );
  AOI22X1 U566 ( .A(n560), .B(n497), .C(n1459), .D(n225), .Y(n558) );
  OAI21X1 U569 ( .A(n328), .B(n168), .C(n562), .Y(n560) );
  OAI21X1 U570 ( .A(n149), .B(n168), .C(currentPlainKey[39]), .Y(n562) );
  OAI21X1 U580 ( .A(n200), .B(n168), .C(n575), .Y(n574) );
  OAI21X1 U581 ( .A(n202), .B(n168), .C(currentPlainKey[38]), .Y(n575) );
  AOI22X1 U595 ( .A(n588), .B(n524), .C(n1460), .D(RCV_DATA[1]), .Y(n586) );
  OAI21X1 U598 ( .A(n358), .B(n168), .C(n589), .Y(n588) );
  OAI21X1 U599 ( .A(n220), .B(n168), .C(currentPlainKey[37]), .Y(n589) );
  OAI21X1 U609 ( .A(n236), .B(n168), .C(n602), .Y(n601) );
  OAI21X1 U610 ( .A(n238), .B(n168), .C(currentPlainKey[36]), .Y(n602) );
  AOI22X1 U624 ( .A(n615), .B(n553), .C(n1461), .D(n225), .Y(n613) );
  OAI21X1 U627 ( .A(n388), .B(n168), .C(n616), .Y(n615) );
  OAI21X1 U628 ( .A(n256), .B(n168), .C(currentPlainKey[35]), .Y(n616) );
  OAI21X1 U638 ( .A(n402), .B(n168), .C(n629), .Y(n628) );
  OAI21X1 U639 ( .A(n276), .B(n168), .C(currentPlainKey[34]), .Y(n629) );
  AOI22X1 U653 ( .A(n642), .B(n581), .C(n1462), .D(n225), .Y(n640) );
  OAI21X1 U658 ( .A(n292), .B(n168), .C(n643), .Y(n642) );
  OAI21X1 U659 ( .A(n294), .B(n168), .C(currentPlainKey[33]), .Y(n643) );
  OAI21X1 U669 ( .A(n307), .B(n168), .C(n656), .Y(n655) );
  OAI21X1 U670 ( .A(n309), .B(n168), .C(currentPlainKey[32]), .Y(n656) );
  NOR2X1 U672 ( .A(n1508), .B(address[4]), .Y(n546) );
  AOI22X1 U686 ( .A(n671), .B(n608), .C(n1463), .D(n225), .Y(n669) );
  OAI21X1 U689 ( .A(n328), .B(n166), .C(n673), .Y(n671) );
  OAI21X1 U690 ( .A(n149), .B(n166), .C(currentPlainKey[31]), .Y(n673) );
  OAI21X1 U700 ( .A(n200), .B(n166), .C(n686), .Y(n685) );
  OAI21X1 U701 ( .A(n202), .B(n166), .C(currentPlainKey[30]), .Y(n686) );
  AOI22X1 U715 ( .A(n699), .B(n635), .C(n1464), .D(n225), .Y(n697) );
  OAI21X1 U718 ( .A(n358), .B(n166), .C(n700), .Y(n699) );
  OAI21X1 U719 ( .A(n220), .B(n166), .C(currentPlainKey[29]), .Y(n700) );
  OAI21X1 U729 ( .A(n236), .B(n166), .C(n713), .Y(n712) );
  OAI21X1 U730 ( .A(n238), .B(n166), .C(currentPlainKey[28]), .Y(n713) );
  AOI22X1 U744 ( .A(n726), .B(n664), .C(n1465), .D(n225), .Y(n724) );
  OAI21X1 U747 ( .A(n388), .B(n166), .C(n727), .Y(n726) );
  OAI21X1 U748 ( .A(n256), .B(n166), .C(currentPlainKey[27]), .Y(n727) );
  OAI21X1 U758 ( .A(n402), .B(n166), .C(n740), .Y(n739) );
  OAI21X1 U759 ( .A(n276), .B(n166), .C(currentPlainKey[26]), .Y(n740) );
  AOI22X1 U773 ( .A(n753), .B(n692), .C(n1466), .D(n225), .Y(n751) );
  OAI21X1 U776 ( .A(n292), .B(n166), .C(n754), .Y(n753) );
  OAI21X1 U777 ( .A(n294), .B(n166), .C(currentPlainKey[25]), .Y(n754) );
  OAI21X1 U787 ( .A(n307), .B(n166), .C(n767), .Y(n766) );
  OAI21X1 U788 ( .A(n309), .B(n166), .C(currentPlainKey[24]), .Y(n767) );
  AOI22X1 U803 ( .A(n782), .B(n719), .C(n1467), .D(n225), .Y(n780) );
  OAI21X1 U806 ( .A(n328), .B(n165), .C(n784), .Y(n782) );
  OAI21X1 U807 ( .A(n149), .B(n165), .C(currentPlainKey[23]), .Y(n784) );
  OAI21X1 U817 ( .A(n200), .B(n165), .C(n797), .Y(n796) );
  OAI21X1 U818 ( .A(n202), .B(n165), .C(currentPlainKey[22]), .Y(n797) );
  AOI22X1 U832 ( .A(n810), .B(n746), .C(n1468), .D(n225), .Y(n808) );
  OAI21X1 U835 ( .A(n358), .B(n165), .C(n811), .Y(n810) );
  OAI21X1 U836 ( .A(n220), .B(n165), .C(currentPlainKey[21]), .Y(n811) );
  OAI21X1 U846 ( .A(n236), .B(n165), .C(n824), .Y(n823) );
  OAI21X1 U847 ( .A(n238), .B(n165), .C(currentPlainKey[20]), .Y(n824) );
  AOI22X1 U861 ( .A(n837), .B(n775), .C(n1469), .D(n225), .Y(n835) );
  OAI21X1 U864 ( .A(n388), .B(n165), .C(n838), .Y(n837) );
  OAI21X1 U865 ( .A(n256), .B(n165), .C(currentPlainKey[19]), .Y(n838) );
  OAI21X1 U875 ( .A(n402), .B(n165), .C(n851), .Y(n850) );
  OAI21X1 U876 ( .A(n276), .B(n165), .C(currentPlainKey[18]), .Y(n851) );
  AOI22X1 U890 ( .A(n864), .B(n803), .C(n1470), .D(n225), .Y(n862) );
  OAI21X1 U895 ( .A(n292), .B(n165), .C(n865), .Y(n864) );
  OAI21X1 U896 ( .A(n294), .B(n165), .C(currentPlainKey[17]), .Y(n865) );
  OAI21X1 U906 ( .A(n307), .B(n165), .C(n878), .Y(n877) );
  OAI21X1 U907 ( .A(n309), .B(n165), .C(currentPlainKey[16]), .Y(n878) );
  NOR2X1 U909 ( .A(n1509), .B(address[5]), .Y(n768) );
  AOI22X1 U923 ( .A(n893), .B(n830), .C(n1471), .D(n225), .Y(n891) );
  OAI21X1 U926 ( .A(n328), .B(n161), .C(n895), .Y(n893) );
  OAI21X1 U927 ( .A(n149), .B(n161), .C(currentPlainKey[15]), .Y(n895) );
  OAI21X1 U937 ( .A(n200), .B(n161), .C(n908), .Y(n907) );
  OAI21X1 U938 ( .A(n202), .B(n161), .C(currentPlainKey[14]), .Y(n908) );
  AOI22X1 U952 ( .A(n921), .B(n857), .C(n1472), .D(n225), .Y(n919) );
  OAI21X1 U955 ( .A(n358), .B(n161), .C(n922), .Y(n921) );
  OAI21X1 U956 ( .A(n220), .B(n161), .C(currentPlainKey[13]), .Y(n922) );
  OAI21X1 U966 ( .A(n236), .B(n161), .C(n935), .Y(n934) );
  OAI21X1 U967 ( .A(n238), .B(n161), .C(currentPlainKey[12]), .Y(n935) );
  AOI22X1 U981 ( .A(n948), .B(n886), .C(n1473), .D(n225), .Y(n946) );
  OAI21X1 U984 ( .A(n388), .B(n161), .C(n949), .Y(n948) );
  OAI21X1 U985 ( .A(n256), .B(n161), .C(currentPlainKey[11]), .Y(n949) );
  OAI21X1 U995 ( .A(n402), .B(n161), .C(n962), .Y(n961) );
  OAI21X1 U996 ( .A(n276), .B(n161), .C(currentPlainKey[10]), .Y(n962) );
  AOI22X1 U1010 ( .A(n975), .B(n914), .C(n1474), .D(n225), .Y(n973) );
  OAI21X1 U1014 ( .A(n292), .B(n161), .C(n976), .Y(n975) );
  OAI21X1 U1015 ( .A(n294), .B(n161), .C(currentPlainKey[9]), .Y(n976) );
  OAI21X1 U1025 ( .A(n307), .B(n161), .C(n989), .Y(n988) );
  OAI21X1 U1026 ( .A(n309), .B(n161), .C(currentPlainKey[8]), .Y(n989) );
  AOI22X1 U1041 ( .A(n1004), .B(n941), .C(n1475), .D(n225), .Y(n1002) );
  OAI21X1 U1044 ( .A(n328), .B(n160), .C(n1006), .Y(n1004) );
  OAI21X1 U1045 ( .A(n149), .B(n160), .C(currentPlainKey[7]), .Y(n1006) );
  NAND2X1 U1046 ( .A(n158), .B(n16), .Y(n328) );
  OAI21X1 U1057 ( .A(n200), .B(n160), .C(n1019), .Y(n1018) );
  OAI21X1 U1058 ( .A(n202), .B(n160), .C(currentPlainKey[6]), .Y(n1019) );
  NAND2X1 U1059 ( .A(n158), .B(n147), .Y(n200) );
  AOI22X1 U1074 ( .A(n1033), .B(n968), .C(n1476), .D(n225), .Y(n1031) );
  OAI21X1 U1077 ( .A(n358), .B(n160), .C(n1034), .Y(n1033) );
  OAI21X1 U1078 ( .A(n220), .B(n160), .C(currentPlainKey[5]), .Y(n1034) );
  NAND2X1 U1079 ( .A(n158), .B(n1478), .Y(n358) );
  OAI21X1 U1090 ( .A(n236), .B(n160), .C(n1047), .Y(n1046) );
  OAI21X1 U1091 ( .A(n238), .B(n160), .C(currentPlainKey[4]), .Y(n1047) );
  NAND2X1 U1092 ( .A(n158), .B(n150), .Y(n236) );
  OAI21X1 U1111 ( .A(n388), .B(n160), .C(n1063), .Y(n1062) );
  OAI21X1 U1112 ( .A(n256), .B(n160), .C(currentPlainKey[3]), .Y(n1063) );
  NAND2X1 U1113 ( .A(n158), .B(n1481), .Y(n388) );
  OAI21X1 U1126 ( .A(n402), .B(n160), .C(n1078), .Y(n1077) );
  OAI21X1 U1127 ( .A(n276), .B(n160), .C(currentPlainKey[2]), .Y(n1078) );
  NAND2X1 U1128 ( .A(n158), .B(n151), .Y(n402) );
  NOR2X1 U1154 ( .A(address[6]), .B(address[7]), .Y(n420) );
  OAI21X1 U1155 ( .A(n292), .B(n160), .C(n1090), .Y(n1089) );
  OAI21X1 U1156 ( .A(n294), .B(n160), .C(currentPlainKey[1]), .Y(n1090) );
  NAND2X1 U1157 ( .A(n158), .B(n143), .Y(n292) );
  AOI22X1 U1182 ( .A(n21), .B(n1576), .C(n1103), .D(n1104), .Y(n1101) );
  AOI21X1 U1183 ( .A(n1105), .B(n1038), .C(n21), .Y(n1104) );
  OAI21X1 U1184 ( .A(n226), .B(n1011), .C(n1106), .Y(n1105) );
  NAND2X1 U1185 ( .A(n25), .B(n1107), .Y(n1106) );
  OAI21X1 U1186 ( .A(n307), .B(n160), .C(n1108), .Y(n1107) );
  OAI21X1 U1187 ( .A(n309), .B(n160), .C(currentPlainKey[0]), .Y(n1108) );
  NOR2X1 U1189 ( .A(address[4]), .B(address[5]), .Y(n990) );
  NAND2X1 U1190 ( .A(n158), .B(n1477), .Y(n307) );
  AOI22X1 U1199 ( .A(n1479), .B(RCV_DATA[2]), .C(n1502), .D(RCV_DATA[3]), .Y(
        n1103) );
  NOR2X1 U1220 ( .A(n1508), .B(n1509), .Y(n310) );
  OAI21X1 U1273 ( .A(n1480), .B(n1484), .C(n1143), .Y(n1349) );
  NAND3X1 U1274 ( .A(keyCount[0]), .B(n1484), .C(n1144), .Y(n1143) );
  NAND2X1 U1305 ( .A(n1579), .B(n1574), .Y(n1178) );
  NAND3X1 U1314 ( .A(keyCount[2]), .B(keyCount[1]), .C(n1186), .Y(n1160) );
  NOR2X1 U1315 ( .A(keyCount[3]), .B(n1483), .Y(n1186) );
  AND2X2 U254 ( .A(n239), .B(n164), .Y(n216) );
  keyreg_1_DW01_add_0 r577 ( .A(parityAccumulator), .B({RCV_DATA[7:1], n158}), 
        .CI(1'b0), .SUM({N1799, N1798, N1797, N1796, N1795, N1794, N1793, 
        N1792}) );
  DFFSR \state_reg[3]  ( .D(n1354), .CLK(CLK), .R(n243), .S(1'b1), .Q(state[3]) );
  DFFSR \state_reg[2]  ( .D(n1352), .CLK(CLK), .R(n243), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[0]  ( .D(n1353), .CLK(CLK), .R(n243), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[1]  ( .D(n1351), .CLK(CLK), .R(n243), .S(1'b1), .Q(state[1]) );
  DFFSR parityError_reg ( .D(nextParityError), .CLK(CLK), .R(n243), .S(1'b1), 
        .Q(parityError) );
  DFFSR PARITY_ERROR_reg ( .D(nextParityError), .CLK(CLK), .R(n243), .S(1'b1), 
        .Q(PARITY_ERROR) );
  INVX4 U3 ( .A(n327), .Y(n1363) );
  BUFX4 U4 ( .A(n1363), .Y(n210) );
  BUFX4 U5 ( .A(n1363), .Y(n209) );
  BUFX4 U7 ( .A(n1363), .Y(n217) );
  INVX1 U8 ( .A(n1367), .Y(n1) );
  INVX1 U23 ( .A(n1367), .Y(n2) );
  INVX1 U26 ( .A(n1367), .Y(n4) );
  INVX8 U29 ( .A(n1174), .Y(n1367) );
  INVX2 U32 ( .A(n1172), .Y(n1184) );
  BUFX2 U35 ( .A(n1184), .Y(n195) );
  BUFX2 U38 ( .A(n1417), .Y(n89) );
  BUFX2 U41 ( .A(n1370), .Y(n224) );
  BUFX2 U44 ( .A(n1370), .Y(n219) );
  INVX2 U47 ( .A(n1409), .Y(n5) );
  INVX2 U50 ( .A(n5), .Y(n6) );
  INVX1 U53 ( .A(n5), .Y(n7) );
  AND2X2 U56 ( .A(n105), .B(n1482), .Y(n8) );
  AND2X2 U59 ( .A(n107), .B(n1482), .Y(n9) );
  AND2X2 U62 ( .A(n109), .B(n1482), .Y(n10) );
  AND2X2 U65 ( .A(n14), .B(n1482), .Y(n11) );
  INVX2 U68 ( .A(n139), .Y(n141) );
  AND2X2 U71 ( .A(n310), .B(n420), .Y(n14) );
  AND2X2 U74 ( .A(n65), .B(address[0]), .Y(n16) );
  INVX2 U77 ( .A(n95), .Y(n178) );
  INVX2 U80 ( .A(n178), .Y(n177) );
  NAND2X1 U83 ( .A(n177), .B(RCV_DATA[3]), .Y(n17) );
  AND2X2 U86 ( .A(n131), .B(n141), .Y(n19) );
  AND2X2 U89 ( .A(n1481), .B(address[3]), .Y(n20) );
  AND2X2 U92 ( .A(n271), .B(n29), .Y(n21) );
  AND2X2 U95 ( .A(n271), .B(n20), .Y(n23) );
  INVX2 U98 ( .A(n189), .Y(n185) );
  INVX2 U101 ( .A(n189), .Y(n186) );
  INVX2 U104 ( .A(n131), .Y(n133) );
  AND2X2 U107 ( .A(n300), .B(n1011), .Y(n25) );
  AND2X2 U110 ( .A(n151), .B(address[3]), .Y(n27) );
  AND2X2 U113 ( .A(n150), .B(address[3]), .Y(n29) );
  AND2X2 U116 ( .A(n1478), .B(address[3]), .Y(n31) );
  AND2X2 U119 ( .A(n147), .B(address[3]), .Y(n33) );
  AND2X2 U122 ( .A(n16), .B(address[3]), .Y(n35) );
  AND2X2 U125 ( .A(n1477), .B(address[3]), .Y(n37) );
  AND2X2 U128 ( .A(n319), .B(n347), .Y(n39) );
  AND2X2 U131 ( .A(n410), .B(n1016), .Y(n41) );
  AND2X2 U134 ( .A(n470), .B(n955), .Y(n43) );
  AND2X2 U137 ( .A(n914), .B(n460), .Y(n45) );
  AND2X2 U140 ( .A(n857), .B(n522), .Y(n47) );
  AND2X2 U143 ( .A(n692), .B(n707), .Y(n49) );
  AND2X2 U146 ( .A(n635), .B(n770), .Y(n51) );
  AND2X2 U149 ( .A(n968), .B(n397), .Y(n53) );
  AND2X2 U152 ( .A(n803), .B(n584), .Y(n55) );
  AND2X2 U155 ( .A(n746), .B(n647), .Y(n57) );
  AND2X2 U158 ( .A(n581), .B(n831), .Y(n59) );
  AND2X2 U161 ( .A(n524), .B(n892), .Y(n61) );
  AND2X2 U164 ( .A(n349), .B(n1074), .Y(n63) );
  AND2X2 U167 ( .A(address[1]), .B(address[2]), .Y(n65) );
  AND2X2 U170 ( .A(n216), .B(n235), .Y(n67) );
  AND2X2 U173 ( .A(n271), .B(n27), .Y(n69) );
  INVX1 U198 ( .A(n332), .Y(n333) );
  AND2X2 U199 ( .A(n85), .B(RCV_DATA[1]), .Y(n99) );
  AND2X1 U200 ( .A(n117), .B(n19), .Y(n83) );
  INVX1 U201 ( .A(n83), .Y(n1432) );
  BUFX2 U204 ( .A(n177), .Y(n85) );
  BUFX4 U207 ( .A(n177), .Y(n87) );
  AND2X2 U209 ( .A(n91), .B(n1263), .Y(n1164) );
  NOR2X1 U212 ( .A(n1162), .B(n1450), .Y(n91) );
  INVX2 U214 ( .A(n226), .Y(n225) );
  BUFX2 U215 ( .A(n17), .Y(n97) );
  INVX2 U216 ( .A(n184), .Y(n180) );
  INVX2 U217 ( .A(n1387), .Y(n93) );
  AND2X2 U218 ( .A(n101), .B(n1425), .Y(n95) );
  INVX1 U219 ( .A(n95), .Y(n1364) );
  INVX2 U228 ( .A(n178), .Y(n175) );
  INVX4 U229 ( .A(n153), .Y(n1136) );
  INVX2 U230 ( .A(n156), .Y(n158) );
  AND2X1 U231 ( .A(n177), .B(RCV_DATA[2]), .Y(n119) );
  INVX2 U232 ( .A(n240), .Y(n230) );
  INVX2 U237 ( .A(n240), .Y(n229) );
  INVX2 U241 ( .A(n234), .Y(n228) );
  INVX2 U243 ( .A(n234), .Y(n227) );
  INVX2 U244 ( .A(n241), .Y(n231) );
  INVX2 U245 ( .A(n241), .Y(n232) );
  INVX2 U246 ( .A(n242), .Y(n233) );
  INVX2 U247 ( .A(n208), .Y(n207) );
  BUFX2 U248 ( .A(n243), .Y(n241) );
  BUFX2 U249 ( .A(n241), .Y(n240) );
  BUFX2 U250 ( .A(n242), .Y(n234) );
  BUFX2 U251 ( .A(n243), .Y(n242) );
  INVX2 U255 ( .A(n99), .Y(n154) );
  INVX2 U256 ( .A(n99), .Y(n153) );
  INVX2 U257 ( .A(n208), .Y(n206) );
  INVX2 U258 ( .A(n208), .Y(n205) );
  INVX2 U259 ( .A(RST), .Y(n243) );
  BUFX2 U260 ( .A(n1370), .Y(n221) );
  BUFX2 U261 ( .A(n1370), .Y(n222) );
  BUFX2 U262 ( .A(n1370), .Y(n223) );
  INVX2 U263 ( .A(n184), .Y(n181) );
  BUFX2 U267 ( .A(n1184), .Y(n197) );
  BUFX2 U268 ( .A(n1184), .Y(n193) );
  BUFX2 U269 ( .A(n1184), .Y(n192) );
  AND2X2 U272 ( .A(n269), .B(n1419), .Y(n101) );
  INVX2 U273 ( .A(n184), .Y(n183) );
  INVX2 U274 ( .A(n188), .Y(n187) );
  BUFX2 U275 ( .A(n1184), .Y(n203) );
  INVX2 U276 ( .A(n103), .Y(n160) );
  INVX2 U277 ( .A(n111), .Y(n173) );
  INVX2 U278 ( .A(n113), .Y(n165) );
  INVX2 U279 ( .A(n115), .Y(n168) );
  INVX2 U280 ( .A(n17), .Y(n184) );
  BUFX2 U281 ( .A(n119), .Y(n188) );
  AND2X2 U282 ( .A(n990), .B(n1482), .Y(n103) );
  AND2X2 U283 ( .A(n546), .B(n420), .Y(n105) );
  AND2X2 U286 ( .A(n990), .B(n420), .Y(n107) );
  AND2X2 U288 ( .A(n768), .B(n420), .Y(n109) );
  INVX2 U289 ( .A(n202), .Y(n147) );
  AND2X2 U290 ( .A(n310), .B(n1482), .Y(n111) );
  AND2X2 U291 ( .A(n768), .B(n1482), .Y(n113) );
  AND2X2 U292 ( .A(n546), .B(n1482), .Y(n115) );
  INVX2 U293 ( .A(n121), .Y(n161) );
  INVX2 U294 ( .A(n123), .Y(n166) );
  INVX2 U295 ( .A(n125), .Y(n172) );
  INVX2 U296 ( .A(RCV_DATA[1]), .Y(n226) );
  AND2X2 U297 ( .A(state[1]), .B(n1417), .Y(n117) );
  INVX2 U298 ( .A(RCV_DATA[0]), .Y(n156) );
  INVX2 U299 ( .A(n294), .Y(n143) );
  INVX2 U301 ( .A(n238), .Y(n150) );
  INVX2 U302 ( .A(n276), .Y(n151) );
  INVX2 U305 ( .A(n16), .Y(n149) );
  AND2X2 U306 ( .A(n990), .B(address[3]), .Y(n121) );
  AND2X2 U307 ( .A(n768), .B(address[3]), .Y(n123) );
  AND2X2 U308 ( .A(n546), .B(address[3]), .Y(n125) );
  BUFX2 U309 ( .A(n101), .Y(n208) );
  AND2X2 U310 ( .A(n259), .B(n129), .Y(n127) );
  BUFX2 U311 ( .A(n1430), .Y(n129) );
  AND2X1 U312 ( .A(n129), .B(n93), .Y(n1423) );
  INVX2 U313 ( .A(state[2]), .Y(n131) );
  NOR2X1 U317 ( .A(state[1]), .B(n141), .Y(n135) );
  INVX1 U318 ( .A(n135), .Y(n1413) );
  INVX1 U319 ( .A(state[1]), .Y(n250) );
  INVX2 U320 ( .A(n188), .Y(n137) );
  INVX2 U321 ( .A(state[0]), .Y(n139) );
  INVX1 U322 ( .A(n7), .Y(n1397) );
  INVX1 U323 ( .A(n7), .Y(n1406) );
  INVX1 U324 ( .A(n7), .Y(n1395) );
  INVX1 U325 ( .A(n7), .Y(n1403) );
  INVX1 U326 ( .A(n7), .Y(n1401) );
  INVX1 U327 ( .A(n7), .Y(n1399) );
  INVX1 U328 ( .A(n7), .Y(n1408) );
  BUFX2 U329 ( .A(n119), .Y(n189) );
  INVX1 U331 ( .A(n1429), .Y(n249) );
  INVX1 U332 ( .A(n1431), .Y(n1387) );
  INVX2 U335 ( .A(n6), .Y(n145) );
  NAND2X1 U336 ( .A(address[0]), .B(address[1]), .Y(n244) );
  OR2X2 U337 ( .A(address[2]), .B(n244), .Y(n256) );
  INVX2 U338 ( .A(n256), .Y(n1481) );
  NAND2X1 U339 ( .A(n20), .B(n14), .Y(n164) );
  INVX2 U340 ( .A(address[2]), .Y(n267) );
  INVX2 U341 ( .A(address[1]), .Y(n266) );
  NAND3X1 U342 ( .A(address[0]), .B(n267), .C(n266), .Y(n294) );
  NAND2X1 U343 ( .A(n143), .B(address[3]), .Y(n278) );
  INVX2 U346 ( .A(n278), .Y(n925) );
  NAND2X1 U347 ( .A(n925), .B(n14), .Y(n157) );
  INVX2 U348 ( .A(state[3]), .Y(n1417) );
  NAND3X1 U349 ( .A(n117), .B(n139), .C(n131), .Y(n1442) );
  NAND3X1 U350 ( .A(n133), .B(n141), .C(n117), .Y(n1416) );
  NAND2X1 U351 ( .A(n1442), .B(n1416), .Y(CLR_RBUFF) );
  NAND3X1 U352 ( .A(n135), .B(n133), .C(n89), .Y(n245) );
  INVX2 U353 ( .A(n245), .Y(PROG_ERROR) );
  NAND2X1 U354 ( .A(n135), .B(n131), .Y(n1429) );
  OAI21X1 U355 ( .A(state[3]), .B(n1429), .C(n1432), .Y(n248) );
  NAND3X1 U356 ( .A(n117), .B(n133), .C(n139), .Y(n1430) );
  NAND2X1 U357 ( .A(n1430), .B(n245), .Y(n247) );
  NOR3X1 U358 ( .A(CLR_RBUFF), .B(n248), .C(n247), .Y(n1374) );
  NAND2X1 U360 ( .A(state[3]), .B(n249), .Y(n1431) );
  NAND3X1 U361 ( .A(n141), .B(n250), .C(n1417), .Y(n255) );
  INVX2 U364 ( .A(n255), .Y(n257) );
  NAND2X1 U365 ( .A(n257), .B(n133), .Y(n1419) );
  INVX2 U366 ( .A(n1419), .Y(n1439) );
  NAND2X1 U367 ( .A(n257), .B(n131), .Y(n259) );
  INVX2 U368 ( .A(n259), .Y(n1386) );
  AOI21X1 U369 ( .A(n1439), .B(parityError), .C(n1386), .Y(n258) );
  NAND3X1 U370 ( .A(n1374), .B(n1431), .C(n258), .Y(KEY_ERROR) );
  NOR2X1 U371 ( .A(PROG_ERROR), .B(n227), .Y(n261) );
  NAND2X1 U372 ( .A(n259), .B(n1430), .Y(n1424) );
  NOR2X1 U375 ( .A(n83), .B(n1424), .Y(n260) );
  NAND3X1 U376 ( .A(n261), .B(n1431), .C(n260), .Y(n1409) );
  NAND2X1 U377 ( .A(n145), .B(n1416), .Y(n1446) );
  INVX2 U378 ( .A(n1446), .Y(n269) );
  INVX2 U379 ( .A(n1442), .Y(n1425) );
  NAND2X1 U380 ( .A(n269), .B(n1425), .Y(n1448) );
  NOR2X1 U381 ( .A(n1494), .B(n1448), .Y(n1144) );
  NAND2X1 U382 ( .A(keyCount[1]), .B(keyCount[0]), .Y(n262) );
  NAND2X1 U383 ( .A(n1425), .B(n262), .Y(n263) );
  NAND2X1 U384 ( .A(n269), .B(n263), .Y(n1443) );
  INVX2 U385 ( .A(n1443), .Y(n1480) );
  INVX2 U386 ( .A(address[0]), .Y(n268) );
  NAND2X1 U387 ( .A(n65), .B(n268), .Y(n202) );
  NAND3X1 U389 ( .A(address[6]), .B(address[7]), .C(n310), .Y(n277) );
  INVX2 U390 ( .A(n277), .Y(n271) );
  NAND2X1 U393 ( .A(n271), .B(n33), .Y(n300) );
  INVX2 U394 ( .A(n300), .Y(n1479) );
  NAND2X1 U395 ( .A(address[0]), .B(address[2]), .Y(n264) );
  OR2X2 U396 ( .A(address[1]), .B(n264), .Y(n220) );
  INVX2 U397 ( .A(n220), .Y(n1478) );
  NAND2X1 U398 ( .A(n271), .B(n31), .Y(n1038) );
  INVX2 U399 ( .A(n1038), .Y(n1502) );
  NOR2X1 U400 ( .A(address[2]), .B(address[0]), .Y(n265) );
  NAND2X1 U401 ( .A(n265), .B(n266), .Y(n309) );
  INVX2 U404 ( .A(n309), .Y(n1477) );
  INVX2 U405 ( .A(address[3]), .Y(n1482) );
  NAND2X1 U406 ( .A(n271), .B(n35), .Y(n1011) );
  NAND3X1 U407 ( .A(address[2]), .B(n268), .C(n266), .Y(n238) );
  INVX2 U408 ( .A(RCV_DATA[4]), .Y(n1576) );
  NAND3X1 U409 ( .A(address[1]), .B(n268), .C(n267), .Y(n276) );
  NAND2X1 U410 ( .A(n9), .B(n150), .Y(n968) );
  INVX2 U411 ( .A(n968), .Y(n1476) );
  NAND2X1 U412 ( .A(n9), .B(n147), .Y(n941) );
  INVX2 U413 ( .A(n941), .Y(n1475) );
  NAND2X1 U414 ( .A(n107), .B(n37), .Y(n914) );
  INVX2 U415 ( .A(n914), .Y(n1474) );
  NAND2X1 U416 ( .A(n107), .B(n27), .Y(n886) );
  INVX2 U418 ( .A(n886), .Y(n1473) );
  NAND2X1 U419 ( .A(n107), .B(n29), .Y(n857) );
  INVX2 U420 ( .A(n857), .Y(n1472) );
  NAND2X1 U421 ( .A(n107), .B(n33), .Y(n830) );
  INVX2 U424 ( .A(n830), .Y(n1471) );
  NAND2X1 U425 ( .A(n10), .B(n1477), .Y(n803) );
  INVX2 U426 ( .A(n803), .Y(n1470) );
  NAND2X1 U427 ( .A(n10), .B(n151), .Y(n775) );
  INVX2 U428 ( .A(n775), .Y(n1469) );
  NAND2X1 U429 ( .A(n10), .B(n150), .Y(n746) );
  INVX2 U430 ( .A(n746), .Y(n1468) );
  NAND2X1 U431 ( .A(n10), .B(n147), .Y(n719) );
  INVX2 U432 ( .A(n719), .Y(n1467) );
  NAND2X1 U435 ( .A(n109), .B(n37), .Y(n692) );
  INVX2 U436 ( .A(n692), .Y(n1466) );
  NAND2X1 U437 ( .A(n109), .B(n27), .Y(n664) );
  INVX2 U438 ( .A(n664), .Y(n1465) );
  NAND2X1 U439 ( .A(n109), .B(n29), .Y(n635) );
  INVX2 U440 ( .A(n635), .Y(n1464) );
  NAND2X1 U441 ( .A(n109), .B(n33), .Y(n608) );
  INVX2 U442 ( .A(n608), .Y(n1463) );
  NAND2X1 U443 ( .A(n8), .B(n1477), .Y(n581) );
  INVX2 U444 ( .A(n581), .Y(n1462) );
  NAND2X1 U445 ( .A(n8), .B(n151), .Y(n553) );
  INVX2 U446 ( .A(n553), .Y(n1461) );
  NAND2X1 U447 ( .A(n8), .B(n150), .Y(n524) );
  INVX2 U448 ( .A(n524), .Y(n1460) );
  NAND2X1 U450 ( .A(n8), .B(n147), .Y(n497) );
  INVX2 U451 ( .A(n497), .Y(n1459) );
  NAND2X1 U454 ( .A(n105), .B(n37), .Y(n470) );
  INVX2 U455 ( .A(n470), .Y(n1458) );
  NAND2X1 U456 ( .A(n105), .B(n27), .Y(n442) );
  INVX2 U457 ( .A(n442), .Y(n1457) );
  NAND2X1 U458 ( .A(n29), .B(n105), .Y(n410) );
  INVX2 U459 ( .A(n410), .Y(n1456) );
  NAND2X1 U460 ( .A(n33), .B(n105), .Y(n379) );
  INVX2 U461 ( .A(n379), .Y(n1455) );
  NAND2X1 U462 ( .A(n11), .B(n1477), .Y(n349) );
  INVX2 U465 ( .A(n349), .Y(n1454) );
  NAND2X1 U466 ( .A(n11), .B(n151), .Y(n318) );
  INVX2 U467 ( .A(n318), .Y(n1453) );
  NAND2X1 U468 ( .A(n11), .B(n150), .Y(n283) );
  INVX2 U469 ( .A(n283), .Y(n1452) );
  NAND2X1 U470 ( .A(n11), .B(n147), .Y(n246) );
  INVX2 U471 ( .A(n246), .Y(n1451) );
  NAND2X1 U472 ( .A(n37), .B(n14), .Y(n152) );
  INVX2 U473 ( .A(n152), .Y(n1450) );
  NAND2X1 U474 ( .A(n14), .B(n27), .Y(n159) );
  INVX2 U475 ( .A(n159), .Y(n1449) );
  INVX2 U476 ( .A(RCV_DATA[2]), .Y(n1578) );
  INVX2 U477 ( .A(RCV_DATA[3]), .Y(n1577) );
  INVX2 U479 ( .A(RCV_DATA[5]), .Y(n1575) );
  INVX2 U480 ( .A(currentPlainKey[3]), .Y(n1570) );
  INVX2 U483 ( .A(currentPlainKey[2]), .Y(n1571) );
  INVX2 U484 ( .A(currentPlainKey[1]), .Y(n1572) );
  NAND2X1 U485 ( .A(n207), .B(currentPlainKey[0]), .Y(n282) );
  NAND2X1 U486 ( .A(n175), .B(RCV_DATA[5]), .Y(n1174) );
  OAI21X1 U487 ( .A(n23), .B(n1364), .C(n2), .Y(n270) );
  OAI21X1 U488 ( .A(n1101), .B(n23), .C(n270), .Y(n275) );
  NAND2X1 U489 ( .A(RCV_DATA[6]), .B(n85), .Y(n327) );
  MUX2X1 U490 ( .B(n275), .A(n327), .S(n69), .Y(n280) );
  NAND2X1 U491 ( .A(RCV_DATA[7]), .B(n175), .Y(n1358) );
  INVX2 U494 ( .A(n1358), .Y(n1370) );
  NOR2X1 U495 ( .A(n278), .B(n277), .Y(n279) );
  MUX2X1 U496 ( .B(n280), .A(n222), .S(n279), .Y(n281) );
  NAND2X1 U497 ( .A(n282), .B(n281), .Y(n1332) );
  NAND2X1 U498 ( .A(n207), .B(currentPlainKey[1]), .Y(n299) );
  INVX2 U499 ( .A(n1089), .Y(n284) );
  NAND2X1 U500 ( .A(n9), .B(n1477), .Y(n319) );
  INVX2 U501 ( .A(n319), .Y(n382) );
  MUX2X1 U502 ( .B(n284), .A(n226), .S(n382), .Y(n286) );
  NOR2X1 U503 ( .A(n1578), .B(n1011), .Y(n285) );
  AOI21X1 U504 ( .A(n25), .B(n286), .C(n285), .Y(n287) );
  NOR2X1 U505 ( .A(n287), .B(n1364), .Y(n289) );
  AOI21X1 U506 ( .A(n1479), .B(n184), .C(n289), .Y(n291) );
  NAND2X1 U508 ( .A(n177), .B(RCV_DATA[4]), .Y(n1172) );
  MUX2X1 U509 ( .B(n291), .A(n1172), .S(n1502), .Y(n295) );
  MUX2X1 U512 ( .B(n295), .A(n1367), .S(n21), .Y(n296) );
  MUX2X1 U513 ( .B(n296), .A(n327), .S(n23), .Y(n297) );
  MUX2X1 U514 ( .B(n297), .A(n224), .S(n69), .Y(n298) );
  NAND2X1 U515 ( .A(n299), .B(n298), .Y(n1331) );
  NAND2X1 U516 ( .A(n207), .B(currentPlainKey[2]), .Y(n315) );
  NOR2X1 U517 ( .A(n1172), .B(n300), .Y(n311) );
  NAND2X1 U518 ( .A(n9), .B(n143), .Y(n347) );
  NAND2X1 U519 ( .A(n39), .B(n87), .Y(n336) );
  INVX2 U520 ( .A(n1077), .Y(n301) );
  OAI22X1 U523 ( .A(n153), .B(n347), .C(n336), .D(n301), .Y(n303) );
  OAI22X1 U524 ( .A(n1011), .B(n17), .C(n137), .D(n319), .Y(n302) );
  AOI21X1 U525 ( .A(n25), .B(n303), .C(n302), .Y(n304) );
  MUX2X1 U526 ( .B(n304), .A(n1), .S(n1502), .Y(n305) );
  NOR2X1 U527 ( .A(n311), .B(n305), .Y(n312) );
  MUX2X1 U528 ( .B(n312), .A(n327), .S(n21), .Y(n313) );
  MUX2X1 U529 ( .B(n313), .A(n224), .S(n23), .Y(n314) );
  NAND2X1 U530 ( .A(n315), .B(n314), .Y(n1330) );
  NAND2X1 U531 ( .A(n207), .B(currentPlainKey[3]), .Y(n334) );
  NAND2X1 U532 ( .A(n1479), .B(n1367), .Y(n326) );
  INVX2 U533 ( .A(n336), .Y(n316) );
  NAND2X1 U534 ( .A(n1062), .B(n316), .Y(n317) );
  NAND2X1 U535 ( .A(n9), .B(n151), .Y(n348) );
  INVX2 U537 ( .A(n348), .Y(n427) );
  MUX2X1 U538 ( .B(n317), .A(n154), .S(n427), .Y(n321) );
  OAI22X1 U541 ( .A(n97), .B(n319), .C(n137), .D(n347), .Y(n320) );
  OAI21X1 U542 ( .A(n321), .B(n320), .C(n25), .Y(n324) );
  INVX2 U543 ( .A(n1011), .Y(n377) );
  NAND2X1 U544 ( .A(n195), .B(n377), .Y(n322) );
  NAND3X1 U545 ( .A(n326), .B(n324), .C(n322), .Y(n330) );
  MUX2X1 U546 ( .B(n330), .A(n217), .S(n1502), .Y(n331) );
  MUX2X1 U547 ( .B(n331), .A(n1358), .S(n21), .Y(n332) );
  NAND2X1 U548 ( .A(n334), .B(n333), .Y(n1329) );
  AOI22X1 U549 ( .A(currentPlainKey[4]), .B(n207), .C(n1479), .D(n209), .Y(
        n346) );
  NAND2X1 U552 ( .A(n382), .B(n192), .Y(n343) );
  OAI22X1 U553 ( .A(n181), .B(n347), .C(n186), .D(n348), .Y(n338) );
  NAND2X1 U554 ( .A(n9), .B(n1481), .Y(n387) );
  NAND2X1 U555 ( .A(n348), .B(n387), .Y(n367) );
  INVX2 U556 ( .A(n367), .Y(n425) );
  NAND2X1 U557 ( .A(n1046), .B(n425), .Y(n335) );
  OAI22X1 U558 ( .A(n153), .B(n387), .C(n336), .D(n335), .Y(n337) );
  OAI21X1 U559 ( .A(n338), .B(n337), .C(n25), .Y(n340) );
  NAND2X1 U560 ( .A(n1367), .B(n377), .Y(n339) );
  NAND3X1 U561 ( .A(n343), .B(n340), .C(n339), .Y(n344) );
  MUX2X1 U562 ( .B(n344), .A(n224), .S(n1502), .Y(n345) );
  NAND2X1 U563 ( .A(n346), .B(n345), .Y(n1328) );
  NAND2X1 U564 ( .A(n1479), .B(n224), .Y(n365) );
  INVX2 U565 ( .A(n347), .Y(n408) );
  NAND2X1 U567 ( .A(n408), .B(n192), .Y(n360) );
  NOR2X1 U568 ( .A(n180), .B(n348), .Y(n353) );
  INVX2 U571 ( .A(n1031), .Y(n350) );
  NAND3X1 U572 ( .A(n425), .B(n87), .C(n350), .Y(n351) );
  OAI21X1 U573 ( .A(n186), .B(n387), .C(n351), .Y(n352) );
  OAI21X1 U574 ( .A(n353), .B(n352), .C(n39), .Y(n357) );
  NAND2X1 U575 ( .A(n382), .B(n1367), .Y(n355) );
  NAND3X1 U576 ( .A(n360), .B(n357), .C(n355), .Y(n361) );
  NAND2X1 U577 ( .A(n25), .B(n361), .Y(n364) );
  AND2X2 U578 ( .A(currentPlainKey[5]), .B(n207), .Y(n362) );
  AOI21X1 U579 ( .A(n217), .B(n377), .C(n362), .Y(n363) );
  NAND3X1 U582 ( .A(n365), .B(n364), .C(n363), .Y(n1327) );
  AOI22X1 U583 ( .A(currentPlainKey[6]), .B(n206), .C(n382), .D(n209), .Y(n381) );
  NAND2X1 U584 ( .A(n408), .B(n1367), .Y(n376) );
  NAND2X1 U585 ( .A(n9), .B(n1478), .Y(n397) );
  INVX2 U586 ( .A(n397), .Y(n471) );
  NAND2X1 U587 ( .A(n471), .B(n1136), .Y(n369) );
  NAND2X1 U588 ( .A(n53), .B(n87), .Y(n399) );
  INVX2 U589 ( .A(n399), .Y(n366) );
  NAND2X1 U590 ( .A(n1018), .B(n366), .Y(n368) );
  AOI21X1 U591 ( .A(n369), .B(n368), .C(n367), .Y(n373) );
  OAI22X1 U592 ( .A(n181), .B(n387), .C(n968), .D(n185), .Y(n370) );
  OAI21X1 U593 ( .A(n373), .B(n370), .C(n39), .Y(n375) );
  NAND2X1 U594 ( .A(n427), .B(n192), .Y(n374) );
  NAND3X1 U596 ( .A(n376), .B(n375), .C(n374), .Y(n378) );
  MUX2X1 U597 ( .B(n378), .A(n224), .S(n377), .Y(n380) );
  NAND2X1 U600 ( .A(n381), .B(n380), .Y(n1326) );
  AOI22X1 U601 ( .A(currentPlainKey[7]), .B(n206), .C(n382), .D(n219), .Y(n396) );
  NAND2X1 U602 ( .A(n427), .B(n1367), .Y(n392) );
  NOR2X1 U603 ( .A(n968), .B(n183), .Y(n385) );
  OAI22X1 U604 ( .A(n187), .B(n397), .C(n1002), .D(n399), .Y(n383) );
  OAI21X1 U605 ( .A(n385), .B(n383), .C(n425), .Y(n391) );
  INVX2 U606 ( .A(n387), .Y(n443) );
  NAND2X1 U607 ( .A(n443), .B(n192), .Y(n390) );
  NAND3X1 U608 ( .A(n392), .B(n391), .C(n390), .Y(n393) );
  NAND2X1 U611 ( .A(n39), .B(n393), .Y(n395) );
  NAND2X1 U612 ( .A(n408), .B(n209), .Y(n394) );
  NAND3X1 U613 ( .A(n396), .B(n395), .C(n394), .Y(n1325) );
  AOI22X1 U614 ( .A(currentPlainKey[8]), .B(n207), .C(n427), .D(n209), .Y(n412) );
  NAND2X1 U615 ( .A(n203), .B(n1476), .Y(n407) );
  OAI22X1 U616 ( .A(n181), .B(n397), .C(n941), .D(n185), .Y(n404) );
  NAND2X1 U617 ( .A(n9), .B(n16), .Y(n452) );
  NAND2X1 U618 ( .A(n941), .B(n452), .Y(n432) );
  INVX2 U619 ( .A(n432), .Y(n486) );
  NAND2X1 U620 ( .A(n988), .B(n486), .Y(n398) );
  OAI22X1 U621 ( .A(n153), .B(n452), .C(n399), .D(n398), .Y(n400) );
  OAI21X1 U622 ( .A(n404), .B(n400), .C(n425), .Y(n406) );
  NAND2X1 U623 ( .A(n443), .B(n1367), .Y(n405) );
  NAND3X1 U625 ( .A(n407), .B(n406), .C(n405), .Y(n409) );
  MUX2X1 U626 ( .B(n409), .A(n224), .S(n408), .Y(n411) );
  NAND2X1 U629 ( .A(n412), .B(n411), .Y(n1324) );
  NAND2X1 U630 ( .A(n443), .B(n209), .Y(n430) );
  NAND2X1 U631 ( .A(n471), .B(n192), .Y(n423) );
  NOR2X1 U632 ( .A(n941), .B(n183), .Y(n418) );
  INVX2 U633 ( .A(n973), .Y(n413) );
  NAND3X1 U634 ( .A(n486), .B(n87), .C(n413), .Y(n414) );
  OAI21X1 U635 ( .A(n187), .B(n452), .C(n414), .Y(n416) );
  OAI21X1 U636 ( .A(n418), .B(n416), .C(n53), .Y(n422) );
  NAND2X1 U637 ( .A(n1367), .B(n1476), .Y(n419) );
  NAND3X1 U640 ( .A(n423), .B(n422), .C(n419), .Y(n424) );
  NAND2X1 U641 ( .A(n425), .B(n424), .Y(n429) );
  AND2X2 U642 ( .A(currentPlainKey[9]), .B(n205), .Y(n426) );
  AOI21X1 U643 ( .A(n427), .B(n221), .C(n426), .Y(n428) );
  NAND3X1 U644 ( .A(n430), .B(n429), .C(n428), .Y(n1323) );
  AOI22X1 U645 ( .A(currentPlainKey[10]), .B(n207), .C(n209), .D(n1476), .Y(
        n446) );
  NAND2X1 U646 ( .A(n203), .B(n1475), .Y(n441) );
  NAND2X1 U647 ( .A(n107), .B(n925), .Y(n460) );
  INVX2 U648 ( .A(n460), .Y(n534) );
  NAND2X1 U649 ( .A(n534), .B(n1136), .Y(n436) );
  NAND2X1 U650 ( .A(n45), .B(n87), .Y(n462) );
  INVX2 U651 ( .A(n462), .Y(n431) );
  NAND2X1 U652 ( .A(n961), .B(n431), .Y(n435) );
  AOI21X1 U654 ( .A(n436), .B(n435), .C(n432), .Y(n438) );
  OAI22X1 U655 ( .A(n181), .B(n452), .C(n914), .D(n185), .Y(n437) );
  OAI21X1 U656 ( .A(n438), .B(n437), .C(n53), .Y(n440) );
  NAND2X1 U657 ( .A(n471), .B(n1367), .Y(n439) );
  NAND3X1 U660 ( .A(n441), .B(n440), .C(n439), .Y(n444) );
  MUX2X1 U661 ( .B(n444), .A(n224), .S(n443), .Y(n445) );
  NAND2X1 U662 ( .A(n446), .B(n445), .Y(n1322) );
  AOI22X1 U663 ( .A(currentPlainKey[11]), .B(n206), .C(n219), .D(n1476), .Y(
        n459) );
  NAND2X1 U664 ( .A(n1367), .B(n1475), .Y(n455) );
  NOR2X1 U665 ( .A(n914), .B(n183), .Y(n450) );
  OAI22X1 U666 ( .A(n187), .B(n460), .C(n946), .D(n462), .Y(n448) );
  OAI21X1 U667 ( .A(n450), .B(n448), .C(n486), .Y(n454) );
  INVX2 U668 ( .A(n452), .Y(n506) );
  NAND2X1 U671 ( .A(n506), .B(n192), .Y(n453) );
  NAND3X1 U673 ( .A(n455), .B(n454), .C(n453), .Y(n456) );
  NAND2X1 U674 ( .A(n53), .B(n456), .Y(n458) );
  NAND2X1 U675 ( .A(n471), .B(n209), .Y(n457) );
  NAND3X1 U676 ( .A(n459), .B(n458), .C(n457), .Y(n1321) );
  AOI22X1 U677 ( .A(currentPlainKey[12]), .B(n207), .C(n209), .D(n1475), .Y(
        n474) );
  NAND2X1 U678 ( .A(n203), .B(n1474), .Y(n469) );
  OAI22X1 U679 ( .A(n180), .B(n460), .C(n886), .D(n185), .Y(n466) );
  NAND2X1 U680 ( .A(n107), .B(n20), .Y(n512) );
  NAND2X1 U681 ( .A(n886), .B(n512), .Y(n494) );
  INVX2 U682 ( .A(n494), .Y(n549) );
  NAND2X1 U683 ( .A(n934), .B(n549), .Y(n461) );
  OAI22X1 U684 ( .A(n153), .B(n512), .C(n462), .D(n461), .Y(n465) );
  OAI21X1 U685 ( .A(n466), .B(n465), .C(n486), .Y(n468) );
  NAND2X1 U687 ( .A(n506), .B(n1367), .Y(n467) );
  NAND3X1 U688 ( .A(n469), .B(n468), .C(n467), .Y(n472) );
  MUX2X1 U691 ( .B(n472), .A(n224), .S(n471), .Y(n473) );
  NAND2X1 U692 ( .A(n474), .B(n473), .Y(n1320) );
  NAND2X1 U693 ( .A(n506), .B(n209), .Y(n492) );
  NAND2X1 U694 ( .A(n534), .B(n192), .Y(n484) );
  NOR2X1 U695 ( .A(n886), .B(n183), .Y(n481) );
  INVX2 U696 ( .A(n919), .Y(n476) );
  NAND3X1 U697 ( .A(n549), .B(n175), .C(n476), .Y(n479) );
  OAI21X1 U698 ( .A(n187), .B(n512), .C(n479), .Y(n480) );
  OAI21X1 U699 ( .A(n481), .B(n480), .C(n45), .Y(n483) );
  NAND2X1 U702 ( .A(n1367), .B(n1474), .Y(n482) );
  NAND3X1 U703 ( .A(n484), .B(n483), .C(n482), .Y(n485) );
  NAND2X1 U704 ( .A(n486), .B(n485), .Y(n489) );
  AND2X2 U705 ( .A(currentPlainKey[13]), .B(n207), .Y(n487) );
  AOI21X1 U706 ( .A(n221), .B(n1475), .C(n487), .Y(n488) );
  NAND3X1 U707 ( .A(n492), .B(n489), .C(n488), .Y(n1319) );
  AOI22X1 U708 ( .A(currentPlainKey[14]), .B(n207), .C(n209), .D(n1474), .Y(
        n509) );
  NAND2X1 U709 ( .A(n203), .B(n1473), .Y(n503) );
  NAND2X1 U710 ( .A(n107), .B(n31), .Y(n522) );
  INVX2 U711 ( .A(n522), .Y(n595) );
  NAND2X1 U712 ( .A(n595), .B(n1136), .Y(n496) );
  NAND2X1 U713 ( .A(n47), .B(n85), .Y(n525) );
  INVX2 U714 ( .A(n525), .Y(n493) );
  NAND2X1 U716 ( .A(n907), .B(n493), .Y(n495) );
  AOI21X1 U717 ( .A(n496), .B(n495), .C(n494), .Y(n499) );
  OAI22X1 U720 ( .A(n97), .B(n512), .C(n857), .D(n185), .Y(n498) );
  OAI21X1 U721 ( .A(n499), .B(n498), .C(n45), .Y(n501) );
  NAND2X1 U722 ( .A(n534), .B(n1367), .Y(n500) );
  NAND3X1 U723 ( .A(n503), .B(n501), .C(n500), .Y(n507) );
  MUX2X1 U724 ( .B(n507), .A(n224), .S(n506), .Y(n508) );
  NAND2X1 U725 ( .A(n509), .B(n508), .Y(n1318) );
  AOI22X1 U726 ( .A(currentPlainKey[15]), .B(n206), .C(n219), .D(n1474), .Y(
        n521) );
  NAND2X1 U727 ( .A(n1367), .B(n1473), .Y(n515) );
  NOR2X1 U728 ( .A(n857), .B(n181), .Y(n511) );
  OAI22X1 U731 ( .A(n187), .B(n522), .C(n891), .D(n525), .Y(n510) );
  OAI21X1 U732 ( .A(n511), .B(n510), .C(n549), .Y(n514) );
  INVX2 U733 ( .A(n512), .Y(n567) );
  NAND2X1 U734 ( .A(n567), .B(n192), .Y(n513) );
  NAND3X1 U735 ( .A(n515), .B(n514), .C(n513), .Y(n516) );
  NAND2X1 U736 ( .A(n45), .B(n516), .Y(n520) );
  NAND2X1 U737 ( .A(n534), .B(n209), .Y(n519) );
  NAND3X1 U738 ( .A(n521), .B(n520), .C(n519), .Y(n1317) );
  AOI22X1 U739 ( .A(currentPlainKey[16]), .B(n206), .C(n210), .D(n1473), .Y(
        n537) );
  NAND2X1 U740 ( .A(n203), .B(n1472), .Y(n533) );
  OAI22X1 U741 ( .A(n97), .B(n522), .C(n830), .D(n186), .Y(n527) );
  NAND2X1 U742 ( .A(n107), .B(n35), .Y(n573) );
  NAND2X1 U743 ( .A(n830), .B(n573), .Y(n556) );
  INVX2 U745 ( .A(n556), .Y(n610) );
  NAND2X1 U746 ( .A(n877), .B(n610), .Y(n523) );
  OAI22X1 U749 ( .A(n154), .B(n573), .C(n525), .D(n523), .Y(n526) );
  OAI21X1 U750 ( .A(n527), .B(n526), .C(n549), .Y(n530) );
  NAND2X1 U751 ( .A(n567), .B(n1367), .Y(n528) );
  NAND3X1 U752 ( .A(n533), .B(n530), .C(n528), .Y(n535) );
  MUX2X1 U753 ( .B(n535), .A(n224), .S(n534), .Y(n536) );
  NAND2X1 U754 ( .A(n537), .B(n536), .Y(n1316) );
  NAND2X1 U755 ( .A(n567), .B(n209), .Y(n554) );
  NAND2X1 U756 ( .A(n595), .B(n192), .Y(n547) );
  NOR2X1 U757 ( .A(n830), .B(n181), .Y(n541) );
  INVX2 U760 ( .A(n862), .Y(n538) );
  NAND3X1 U761 ( .A(n610), .B(n87), .C(n538), .Y(n539) );
  OAI21X1 U762 ( .A(n186), .B(n573), .C(n539), .Y(n540) );
  OAI21X1 U763 ( .A(n541), .B(n540), .C(n47), .Y(n543) );
  NAND2X1 U764 ( .A(n1367), .B(n1472), .Y(n542) );
  NAND3X1 U765 ( .A(n547), .B(n543), .C(n542), .Y(n548) );
  NAND2X1 U766 ( .A(n549), .B(n548), .Y(n552) );
  AND2X2 U767 ( .A(currentPlainKey[17]), .B(n207), .Y(n550) );
  AOI21X1 U768 ( .A(n221), .B(n1473), .C(n550), .Y(n551) );
  NAND3X1 U769 ( .A(n554), .B(n552), .C(n551), .Y(n1315) );
  AOI22X1 U770 ( .A(currentPlainKey[18]), .B(n206), .C(n209), .D(n1472), .Y(
        n570) );
  NAND2X1 U771 ( .A(n203), .B(n1471), .Y(n566) );
  NAND2X1 U772 ( .A(n10), .B(n143), .Y(n584) );
  INVX2 U774 ( .A(n584), .Y(n657) );
  NAND2X1 U775 ( .A(n657), .B(n1136), .Y(n559) );
  NAND2X1 U778 ( .A(n55), .B(n87), .Y(n587) );
  INVX2 U779 ( .A(n587), .Y(n555) );
  NAND2X1 U780 ( .A(n850), .B(n555), .Y(n557) );
  AOI21X1 U781 ( .A(n559), .B(n557), .C(n556), .Y(n563) );
  OAI22X1 U782 ( .A(n180), .B(n573), .C(n803), .D(n185), .Y(n561) );
  OAI21X1 U783 ( .A(n563), .B(n561), .C(n47), .Y(n565) );
  NAND2X1 U784 ( .A(n595), .B(n1367), .Y(n564) );
  NAND3X1 U785 ( .A(n566), .B(n565), .C(n564), .Y(n568) );
  MUX2X1 U786 ( .B(n568), .A(n223), .S(n567), .Y(n569) );
  NAND2X1 U789 ( .A(n570), .B(n569), .Y(n1314) );
  AOI22X1 U790 ( .A(currentPlainKey[19]), .B(n206), .C(n219), .D(n1472), .Y(
        n583) );
  NAND2X1 U791 ( .A(n1367), .B(n1471), .Y(n578) );
  NOR2X1 U792 ( .A(n803), .B(n181), .Y(n572) );
  OAI22X1 U793 ( .A(n187), .B(n584), .C(n835), .D(n587), .Y(n571) );
  OAI21X1 U794 ( .A(n572), .B(n571), .C(n610), .Y(n577) );
  INVX2 U795 ( .A(n573), .Y(n627) );
  NAND2X1 U796 ( .A(n627), .B(n193), .Y(n576) );
  NAND3X1 U797 ( .A(n578), .B(n577), .C(n576), .Y(n579) );
  NAND2X1 U798 ( .A(n47), .B(n579), .Y(n582) );
  NAND2X1 U799 ( .A(n595), .B(n210), .Y(n580) );
  NAND3X1 U800 ( .A(n583), .B(n582), .C(n580), .Y(n1313) );
  AOI22X1 U801 ( .A(currentPlainKey[20]), .B(n206), .C(n210), .D(n1471), .Y(
        n598) );
  NAND2X1 U802 ( .A(n203), .B(n1470), .Y(n594) );
  OAI22X1 U804 ( .A(n180), .B(n584), .C(n775), .D(n186), .Y(n591) );
  NAND2X1 U805 ( .A(n10), .B(n1481), .Y(n636) );
  NAND2X1 U808 ( .A(n775), .B(n636), .Y(n619) );
  INVX2 U809 ( .A(n619), .Y(n672) );
  NAND2X1 U810 ( .A(n823), .B(n672), .Y(n585) );
  OAI22X1 U811 ( .A(n154), .B(n636), .C(n587), .D(n585), .Y(n590) );
  OAI21X1 U812 ( .A(n591), .B(n590), .C(n610), .Y(n593) );
  NAND2X1 U813 ( .A(n627), .B(n1367), .Y(n592) );
  NAND3X1 U814 ( .A(n594), .B(n593), .C(n592), .Y(n596) );
  MUX2X1 U815 ( .B(n596), .A(n223), .S(n595), .Y(n597) );
  NAND2X1 U816 ( .A(n598), .B(n597), .Y(n1312) );
  NAND2X1 U819 ( .A(n627), .B(n209), .Y(n617) );
  NAND2X1 U820 ( .A(n657), .B(n193), .Y(n607) );
  NOR2X1 U821 ( .A(n775), .B(n181), .Y(n604) );
  INVX2 U822 ( .A(n808), .Y(n599) );
  NAND3X1 U823 ( .A(n672), .B(n87), .C(n599), .Y(n600) );
  OAI21X1 U824 ( .A(n187), .B(n636), .C(n600), .Y(n603) );
  OAI21X1 U825 ( .A(n604), .B(n603), .C(n55), .Y(n606) );
  NAND2X1 U826 ( .A(n1367), .B(n1470), .Y(n605) );
  NAND3X1 U827 ( .A(n607), .B(n606), .C(n605), .Y(n609) );
  NAND2X1 U828 ( .A(n610), .B(n609), .Y(n614) );
  AND2X2 U829 ( .A(currentPlainKey[21]), .B(n207), .Y(n611) );
  AOI21X1 U830 ( .A(n221), .B(n1471), .C(n611), .Y(n612) );
  NAND3X1 U831 ( .A(n617), .B(n614), .C(n612), .Y(n1311) );
  AOI22X1 U833 ( .A(currentPlainKey[22]), .B(n206), .C(n210), .D(n1470), .Y(
        n632) );
  NAND2X1 U834 ( .A(n197), .B(n1469), .Y(n626) );
  NAND2X1 U837 ( .A(n10), .B(n1478), .Y(n647) );
  INVX2 U838 ( .A(n647), .Y(n717) );
  NAND2X1 U839 ( .A(n717), .B(n1136), .Y(n621) );
  NAND2X1 U840 ( .A(n57), .B(n85), .Y(n649) );
  INVX2 U841 ( .A(n649), .Y(n618) );
  NAND2X1 U842 ( .A(n796), .B(n618), .Y(n620) );
  AOI21X1 U843 ( .A(n621), .B(n620), .C(n619), .Y(n623) );
  OAI22X1 U844 ( .A(n180), .B(n636), .C(n746), .D(n186), .Y(n622) );
  OAI21X1 U845 ( .A(n623), .B(n622), .C(n55), .Y(n625) );
  NAND2X1 U848 ( .A(n657), .B(n1367), .Y(n624) );
  NAND3X1 U849 ( .A(n626), .B(n625), .C(n624), .Y(n630) );
  MUX2X1 U850 ( .B(n630), .A(n223), .S(n627), .Y(n631) );
  NAND2X1 U851 ( .A(n632), .B(n631), .Y(n1310) );
  AOI22X1 U852 ( .A(currentPlainKey[23]), .B(n206), .C(n219), .D(n1470), .Y(
        n646) );
  NAND2X1 U853 ( .A(n1367), .B(n1469), .Y(n639) );
  NOR2X1 U854 ( .A(n746), .B(n181), .Y(n634) );
  OAI22X1 U855 ( .A(n187), .B(n647), .C(n780), .D(n649), .Y(n633) );
  OAI21X1 U856 ( .A(n634), .B(n633), .C(n672), .Y(n638) );
  INVX2 U857 ( .A(n636), .Y(n689) );
  NAND2X1 U858 ( .A(n689), .B(n193), .Y(n637) );
  NAND3X1 U859 ( .A(n639), .B(n638), .C(n637), .Y(n641) );
  NAND2X1 U860 ( .A(n55), .B(n641), .Y(n645) );
  NAND2X1 U862 ( .A(n657), .B(n1363), .Y(n644) );
  NAND3X1 U863 ( .A(n646), .B(n645), .C(n644), .Y(n1309) );
  AOI22X1 U866 ( .A(currentPlainKey[24]), .B(n206), .C(n210), .D(n1469), .Y(
        n660) );
  NAND2X1 U867 ( .A(n197), .B(n1468), .Y(n654) );
  OAI22X1 U868 ( .A(n97), .B(n647), .C(n719), .D(n186), .Y(n651) );
  NAND2X1 U869 ( .A(n10), .B(n16), .Y(n696) );
  NAND2X1 U870 ( .A(n719), .B(n696), .Y(n679) );
  INVX2 U871 ( .A(n679), .Y(n733) );
  NAND2X1 U872 ( .A(n766), .B(n733), .Y(n648) );
  OAI22X1 U873 ( .A(n154), .B(n696), .C(n649), .D(n648), .Y(n650) );
  OAI21X1 U874 ( .A(n651), .B(n650), .C(n672), .Y(n653) );
  NAND2X1 U877 ( .A(n689), .B(n1367), .Y(n652) );
  NAND3X1 U878 ( .A(n654), .B(n653), .C(n652), .Y(n658) );
  MUX2X1 U879 ( .B(n658), .A(n223), .S(n657), .Y(n659) );
  NAND2X1 U880 ( .A(n660), .B(n659), .Y(n1308) );
  NAND2X1 U881 ( .A(n689), .B(n217), .Y(n677) );
  NAND2X1 U882 ( .A(n717), .B(n193), .Y(n668) );
  NOR2X1 U883 ( .A(n719), .B(n181), .Y(n665) );
  INVX2 U884 ( .A(n751), .Y(n661) );
  NAND3X1 U885 ( .A(n733), .B(n175), .C(n661), .Y(n662) );
  OAI21X1 U886 ( .A(n187), .B(n696), .C(n662), .Y(n663) );
  OAI21X1 U887 ( .A(n665), .B(n663), .C(n57), .Y(n667) );
  NAND2X1 U888 ( .A(n1367), .B(n1468), .Y(n666) );
  NAND3X1 U889 ( .A(n668), .B(n667), .C(n666), .Y(n670) );
  NAND2X1 U891 ( .A(n672), .B(n670), .Y(n676) );
  AND2X2 U892 ( .A(currentPlainKey[25]), .B(n206), .Y(n674) );
  AOI21X1 U893 ( .A(n221), .B(n1469), .C(n674), .Y(n675) );
  NAND3X1 U894 ( .A(n677), .B(n676), .C(n675), .Y(n1307) );
  AOI22X1 U897 ( .A(currentPlainKey[26]), .B(n206), .C(n210), .D(n1468), .Y(
        n693) );
  NAND2X1 U898 ( .A(n197), .B(n1467), .Y(n688) );
  NAND2X1 U899 ( .A(n109), .B(n925), .Y(n707) );
  INVX2 U900 ( .A(n707), .Y(n779) );
  NAND2X1 U901 ( .A(n779), .B(n1136), .Y(n681) );
  NAND2X1 U902 ( .A(n49), .B(n87), .Y(n709) );
  INVX2 U903 ( .A(n709), .Y(n678) );
  NAND2X1 U904 ( .A(n739), .B(n678), .Y(n680) );
  AOI21X1 U905 ( .A(n681), .B(n680), .C(n679), .Y(n683) );
  OAI22X1 U908 ( .A(n97), .B(n696), .C(n692), .D(n186), .Y(n682) );
  OAI21X1 U910 ( .A(n683), .B(n682), .C(n57), .Y(n687) );
  NAND2X1 U911 ( .A(n717), .B(n1367), .Y(n684) );
  NAND3X1 U912 ( .A(n688), .B(n687), .C(n684), .Y(n690) );
  MUX2X1 U913 ( .B(n690), .A(n223), .S(n689), .Y(n691) );
  NAND2X1 U914 ( .A(n693), .B(n691), .Y(n1306) );
  AOI22X1 U915 ( .A(currentPlainKey[27]), .B(n206), .C(n219), .D(n1468), .Y(
        n706) );
  NAND2X1 U916 ( .A(n1367), .B(n1467), .Y(n702) );
  NOR2X1 U917 ( .A(n692), .B(n183), .Y(n695) );
  OAI22X1 U918 ( .A(n137), .B(n707), .C(n724), .D(n709), .Y(n694) );
  OAI21X1 U919 ( .A(n695), .B(n694), .C(n733), .Y(n701) );
  INVX2 U920 ( .A(n696), .Y(n750) );
  NAND2X1 U921 ( .A(n750), .B(n192), .Y(n698) );
  NAND3X1 U922 ( .A(n702), .B(n701), .C(n698), .Y(n703) );
  NAND2X1 U924 ( .A(n57), .B(n703), .Y(n705) );
  NAND2X1 U925 ( .A(n717), .B(n217), .Y(n704) );
  NAND3X1 U928 ( .A(n706), .B(n705), .C(n704), .Y(n1305) );
  AOI22X1 U929 ( .A(currentPlainKey[28]), .B(n205), .C(n210), .D(n1467), .Y(
        n721) );
  NAND2X1 U930 ( .A(n197), .B(n1466), .Y(n716) );
  OAI22X1 U931 ( .A(n180), .B(n707), .C(n664), .D(n186), .Y(n711) );
  NAND2X1 U932 ( .A(n109), .B(n20), .Y(n759) );
  NAND2X1 U933 ( .A(n664), .B(n759), .Y(n741) );
  INVX2 U934 ( .A(n741), .Y(n794) );
  NAND2X1 U935 ( .A(n712), .B(n794), .Y(n708) );
  OAI22X1 U936 ( .A(n154), .B(n759), .C(n709), .D(n708), .Y(n710) );
  OAI21X1 U939 ( .A(n711), .B(n710), .C(n733), .Y(n715) );
  NAND2X1 U940 ( .A(n750), .B(n1367), .Y(n714) );
  NAND3X1 U941 ( .A(n716), .B(n715), .C(n714), .Y(n718) );
  MUX2X1 U942 ( .B(n718), .A(n223), .S(n717), .Y(n720) );
  NAND2X1 U943 ( .A(n721), .B(n720), .Y(n1304) );
  NAND2X1 U944 ( .A(n750), .B(n217), .Y(n737) );
  NAND2X1 U945 ( .A(n779), .B(n193), .Y(n731) );
  NOR2X1 U946 ( .A(n664), .B(n181), .Y(n728) );
  INVX2 U947 ( .A(n697), .Y(n722) );
  NAND3X1 U948 ( .A(n794), .B(n85), .C(n722), .Y(n723) );
  OAI21X1 U949 ( .A(n187), .B(n759), .C(n723), .Y(n725) );
  OAI21X1 U950 ( .A(n728), .B(n725), .C(n49), .Y(n730) );
  NAND2X1 U951 ( .A(n1367), .B(n1466), .Y(n729) );
  NAND3X1 U953 ( .A(n731), .B(n730), .C(n729), .Y(n732) );
  NAND2X1 U954 ( .A(n733), .B(n732), .Y(n736) );
  AND2X2 U957 ( .A(currentPlainKey[29]), .B(n207), .Y(n734) );
  AOI21X1 U958 ( .A(n221), .B(n1467), .C(n734), .Y(n735) );
  NAND3X1 U959 ( .A(n737), .B(n736), .C(n735), .Y(n1303) );
  AOI22X1 U960 ( .A(currentPlainKey[30]), .B(n205), .C(n217), .D(n1466), .Y(
        n756) );
  NAND2X1 U961 ( .A(n197), .B(n1465), .Y(n749) );
  NAND2X1 U962 ( .A(n109), .B(n31), .Y(n770) );
  INVX2 U963 ( .A(n770), .Y(n842) );
  NAND2X1 U964 ( .A(n842), .B(n1136), .Y(n743) );
  NAND2X1 U965 ( .A(n51), .B(n87), .Y(n772) );
  INVX2 U968 ( .A(n772), .Y(n738) );
  NAND2X1 U969 ( .A(n685), .B(n738), .Y(n742) );
  AOI21X1 U970 ( .A(n743), .B(n742), .C(n741), .Y(n745) );
  OAI22X1 U971 ( .A(n180), .B(n759), .C(n635), .D(n185), .Y(n744) );
  OAI21X1 U972 ( .A(n745), .B(n744), .C(n49), .Y(n748) );
  NAND2X1 U973 ( .A(n779), .B(n1367), .Y(n747) );
  NAND3X1 U974 ( .A(n749), .B(n748), .C(n747), .Y(n752) );
  MUX2X1 U975 ( .B(n752), .A(n223), .S(n750), .Y(n755) );
  NAND2X1 U976 ( .A(n756), .B(n755), .Y(n1302) );
  AOI22X1 U977 ( .A(currentPlainKey[31]), .B(n205), .C(n219), .D(n1466), .Y(
        n769) );
  NAND2X1 U978 ( .A(n1367), .B(n1465), .Y(n762) );
  NOR2X1 U979 ( .A(n635), .B(n181), .Y(n758) );
  OAI22X1 U980 ( .A(n137), .B(n770), .C(n669), .D(n772), .Y(n757) );
  OAI21X1 U982 ( .A(n758), .B(n757), .C(n794), .Y(n761) );
  INVX2 U983 ( .A(n759), .Y(n814) );
  NAND2X1 U986 ( .A(n814), .B(n195), .Y(n760) );
  NAND3X1 U987 ( .A(n762), .B(n761), .C(n760), .Y(n763) );
  NAND2X1 U988 ( .A(n49), .B(n763), .Y(n765) );
  NAND2X1 U989 ( .A(n779), .B(n217), .Y(n764) );
  NAND3X1 U990 ( .A(n769), .B(n765), .C(n764), .Y(n1301) );
  AOI22X1 U991 ( .A(currentPlainKey[32]), .B(n205), .C(n217), .D(n1465), .Y(
        n785) );
  NAND2X1 U992 ( .A(n197), .B(n1464), .Y(n778) );
  OAI22X1 U993 ( .A(n97), .B(n770), .C(n608), .D(n186), .Y(n774) );
  NAND2X1 U994 ( .A(n109), .B(n35), .Y(n820) );
  NAND2X1 U997 ( .A(n608), .B(n820), .Y(n802) );
  INVX2 U998 ( .A(n802), .Y(n856) );
  NAND2X1 U999 ( .A(n655), .B(n856), .Y(n771) );
  OAI22X1 U1000 ( .A(n154), .B(n820), .C(n772), .D(n771), .Y(n773) );
  OAI21X1 U1001 ( .A(n774), .B(n773), .C(n794), .Y(n777) );
  NAND2X1 U1002 ( .A(n814), .B(n1367), .Y(n776) );
  NAND3X1 U1003 ( .A(n778), .B(n777), .C(n776), .Y(n781) );
  MUX2X1 U1004 ( .B(n781), .A(n223), .S(n779), .Y(n783) );
  NAND2X1 U1005 ( .A(n785), .B(n783), .Y(n1300) );
  NAND2X1 U1006 ( .A(n814), .B(n217), .Y(n800) );
  NAND2X1 U1007 ( .A(n842), .B(n195), .Y(n792) );
  NOR2X1 U1008 ( .A(n608), .B(n181), .Y(n789) );
  INVX2 U1009 ( .A(n640), .Y(n786) );
  NAND3X1 U1011 ( .A(n856), .B(n87), .C(n786), .Y(n787) );
  OAI21X1 U1012 ( .A(n187), .B(n820), .C(n787), .Y(n788) );
  OAI21X1 U1013 ( .A(n789), .B(n788), .C(n51), .Y(n791) );
  NAND2X1 U1016 ( .A(n1367), .B(n1464), .Y(n790) );
  NAND3X1 U1017 ( .A(n792), .B(n791), .C(n790), .Y(n793) );
  NAND2X1 U1018 ( .A(n794), .B(n793), .Y(n799) );
  AND2X2 U1019 ( .A(currentPlainKey[33]), .B(n207), .Y(n795) );
  AOI21X1 U1020 ( .A(n221), .B(n1465), .C(n795), .Y(n798) );
  NAND3X1 U1021 ( .A(n800), .B(n799), .C(n798), .Y(n1299) );
  AOI22X1 U1022 ( .A(currentPlainKey[34]), .B(n205), .C(n210), .D(n1464), .Y(
        n817) );
  NAND2X1 U1023 ( .A(n197), .B(n1463), .Y(n813) );
  NAND2X1 U1024 ( .A(n8), .B(n143), .Y(n831) );
  INVX2 U1027 ( .A(n831), .Y(n902) );
  NAND2X1 U1028 ( .A(n902), .B(n1136), .Y(n805) );
  NAND2X1 U1029 ( .A(n59), .B(n175), .Y(n833) );
  INVX2 U1030 ( .A(n833), .Y(n801) );
  NAND2X1 U1031 ( .A(n628), .B(n801), .Y(n804) );
  AOI21X1 U1032 ( .A(n805), .B(n804), .C(n802), .Y(n807) );
  OAI22X1 U1033 ( .A(n97), .B(n820), .C(n581), .D(n186), .Y(n806) );
  OAI21X1 U1034 ( .A(n807), .B(n806), .C(n51), .Y(n812) );
  NAND2X1 U1035 ( .A(n842), .B(n1367), .Y(n809) );
  NAND3X1 U1036 ( .A(n813), .B(n812), .C(n809), .Y(n815) );
  MUX2X1 U1037 ( .B(n815), .A(n223), .S(n814), .Y(n816) );
  NAND2X1 U1038 ( .A(n817), .B(n816), .Y(n1298) );
  AOI22X1 U1039 ( .A(currentPlainKey[35]), .B(n205), .C(n221), .D(n1464), .Y(
        n829) );
  NAND2X1 U1040 ( .A(n1367), .B(n1463), .Y(n825) );
  NOR2X1 U1042 ( .A(n581), .B(n181), .Y(n819) );
  OAI22X1 U1043 ( .A(n137), .B(n831), .C(n613), .D(n833), .Y(n818) );
  OAI21X1 U1047 ( .A(n819), .B(n818), .C(n856), .Y(n822) );
  INVX2 U1048 ( .A(n820), .Y(n874) );
  NAND2X1 U1049 ( .A(n874), .B(n193), .Y(n821) );
  NAND3X1 U1050 ( .A(n825), .B(n822), .C(n821), .Y(n826) );
  NAND2X1 U1051 ( .A(n51), .B(n826), .Y(n828) );
  NAND2X1 U1052 ( .A(n842), .B(n217), .Y(n827) );
  NAND3X1 U1053 ( .A(n829), .B(n828), .C(n827), .Y(n1297) );
  AOI22X1 U1054 ( .A(currentPlainKey[36]), .B(n205), .C(n217), .D(n1463), .Y(
        n845) );
  NAND2X1 U1055 ( .A(n197), .B(n1462), .Y(n841) );
  OAI22X1 U1056 ( .A(n97), .B(n831), .C(n553), .D(n186), .Y(n836) );
  NAND2X1 U1060 ( .A(n8), .B(n1481), .Y(n882) );
  NAND2X1 U1061 ( .A(n553), .B(n882), .Y(n866) );
  INVX2 U1062 ( .A(n866), .Y(n917) );
  NAND2X1 U1063 ( .A(n601), .B(n917), .Y(n832) );
  OAI22X1 U1064 ( .A(n154), .B(n882), .C(n833), .D(n832), .Y(n834) );
  OAI21X1 U1065 ( .A(n836), .B(n834), .C(n856), .Y(n840) );
  NAND2X1 U1066 ( .A(n874), .B(n1367), .Y(n839) );
  NAND3X1 U1067 ( .A(n841), .B(n840), .C(n839), .Y(n843) );
  MUX2X1 U1068 ( .B(n843), .A(n223), .S(n842), .Y(n844) );
  NAND2X1 U1069 ( .A(n845), .B(n844), .Y(n1296) );
  NAND2X1 U1070 ( .A(n874), .B(n217), .Y(n861) );
  NAND2X1 U1071 ( .A(n902), .B(n195), .Y(n854) );
  NOR2X1 U1072 ( .A(n553), .B(n183), .Y(n849) );
  INVX2 U1073 ( .A(n586), .Y(n846) );
  NAND3X1 U1075 ( .A(n917), .B(n87), .C(n846), .Y(n847) );
  OAI21X1 U1076 ( .A(n185), .B(n882), .C(n847), .Y(n848) );
  OAI21X1 U1080 ( .A(n849), .B(n848), .C(n59), .Y(n853) );
  NAND2X1 U1081 ( .A(n1367), .B(n1462), .Y(n852) );
  NAND3X1 U1082 ( .A(n854), .B(n853), .C(n852), .Y(n855) );
  NAND2X1 U1083 ( .A(n856), .B(n855), .Y(n860) );
  AND2X2 U1084 ( .A(currentPlainKey[37]), .B(n207), .Y(n858) );
  AOI21X1 U1085 ( .A(n222), .B(n1463), .C(n858), .Y(n859) );
  NAND3X1 U1086 ( .A(n861), .B(n860), .C(n859), .Y(n1295) );
  AOI22X1 U1087 ( .A(currentPlainKey[38]), .B(n205), .C(n210), .D(n1462), .Y(
        n879) );
  NAND2X1 U1088 ( .A(n197), .B(n1461), .Y(n873) );
  NAND2X1 U1089 ( .A(n8), .B(n1478), .Y(n892) );
  INVX2 U1093 ( .A(n892), .Y(n965) );
  NAND2X1 U1094 ( .A(n965), .B(n1136), .Y(n868) );
  NAND2X1 U1095 ( .A(n61), .B(n175), .Y(n896) );
  INVX2 U1096 ( .A(n896), .Y(n863) );
  NAND2X1 U1097 ( .A(n574), .B(n863), .Y(n867) );
  AOI21X1 U1098 ( .A(n868), .B(n867), .C(n866), .Y(n870) );
  OAI22X1 U1099 ( .A(n180), .B(n882), .C(n524), .D(n186), .Y(n869) );
  OAI21X1 U1100 ( .A(n870), .B(n869), .C(n59), .Y(n872) );
  NAND2X1 U1101 ( .A(n902), .B(n1367), .Y(n871) );
  NAND3X1 U1102 ( .A(n873), .B(n872), .C(n871), .Y(n875) );
  MUX2X1 U1103 ( .B(n875), .A(n223), .S(n874), .Y(n876) );
  NAND2X1 U1104 ( .A(n879), .B(n876), .Y(n1294) );
  AOI22X1 U1105 ( .A(currentPlainKey[39]), .B(n205), .C(n219), .D(n1462), .Y(
        n890) );
  NAND2X1 U1106 ( .A(n1367), .B(n1461), .Y(n885) );
  NOR2X1 U1107 ( .A(n524), .B(n183), .Y(n881) );
  OAI22X1 U1108 ( .A(n187), .B(n892), .C(n558), .D(n896), .Y(n880) );
  OAI21X1 U1109 ( .A(n881), .B(n880), .C(n917), .Y(n884) );
  INVX2 U1110 ( .A(n882), .Y(n937) );
  NAND2X1 U1114 ( .A(n937), .B(n195), .Y(n883) );
  NAND3X1 U1115 ( .A(n885), .B(n884), .C(n883), .Y(n887) );
  NAND2X1 U1116 ( .A(n59), .B(n887), .Y(n889) );
  NAND2X1 U1117 ( .A(n902), .B(n217), .Y(n888) );
  NAND3X1 U1118 ( .A(n890), .B(n889), .C(n888), .Y(n1293) );
  AOI22X1 U1119 ( .A(currentPlainKey[40]), .B(n205), .C(n210), .D(n1461), .Y(
        n905) );
  NAND2X1 U1120 ( .A(n197), .B(n1460), .Y(n901) );
  OAI22X1 U1121 ( .A(n180), .B(n892), .C(n497), .D(n186), .Y(n898) );
  NAND2X1 U1122 ( .A(n8), .B(n16), .Y(n944) );
  NAND2X1 U1123 ( .A(n497), .B(n944), .Y(n927) );
  INVX2 U1124 ( .A(n927), .Y(n981) );
  NAND2X1 U1125 ( .A(n544), .B(n981), .Y(n894) );
  OAI22X1 U1129 ( .A(n154), .B(n944), .C(n896), .D(n894), .Y(n897) );
  OAI21X1 U1130 ( .A(n898), .B(n897), .C(n917), .Y(n900) );
  NAND2X1 U1131 ( .A(n937), .B(n1367), .Y(n899) );
  NAND3X1 U1132 ( .A(n901), .B(n900), .C(n899), .Y(n903) );
  MUX2X1 U1133 ( .B(n903), .A(n223), .S(n902), .Y(n904) );
  NAND2X1 U1134 ( .A(n905), .B(n904), .Y(n1292) );
  NAND2X1 U1135 ( .A(n937), .B(n217), .Y(n924) );
  NAND2X1 U1136 ( .A(n965), .B(n193), .Y(n915) );
  NOR2X1 U1137 ( .A(n497), .B(n183), .Y(n911) );
  INVX2 U1138 ( .A(n529), .Y(n906) );
  NAND3X1 U1139 ( .A(n981), .B(n87), .C(n906), .Y(n909) );
  OAI21X1 U1140 ( .A(n187), .B(n944), .C(n909), .Y(n910) );
  OAI21X1 U1141 ( .A(n911), .B(n910), .C(n61), .Y(n913) );
  NAND2X1 U1142 ( .A(n1367), .B(n1460), .Y(n912) );
  NAND3X1 U1143 ( .A(n915), .B(n913), .C(n912), .Y(n916) );
  NAND2X1 U1144 ( .A(n917), .B(n916), .Y(n923) );
  AND2X2 U1145 ( .A(currentPlainKey[41]), .B(n207), .Y(n918) );
  AOI21X1 U1146 ( .A(n222), .B(n1461), .C(n918), .Y(n920) );
  NAND3X1 U1147 ( .A(n924), .B(n923), .C(n920), .Y(n1291) );
  AOI22X1 U1148 ( .A(currentPlainKey[42]), .B(n205), .C(n210), .D(n1460), .Y(
        n940) );
  NAND2X1 U1149 ( .A(n197), .B(n1459), .Y(n936) );
  NAND2X1 U1150 ( .A(n105), .B(n925), .Y(n955) );
  INVX2 U1151 ( .A(n955), .Y(n1026) );
  NAND2X1 U1152 ( .A(n1026), .B(n1136), .Y(n929) );
  NAND2X1 U1153 ( .A(n43), .B(n87), .Y(n957) );
  INVX2 U1158 ( .A(n957), .Y(n926) );
  NAND2X1 U1159 ( .A(n517), .B(n926), .Y(n928) );
  AOI21X1 U1160 ( .A(n929), .B(n928), .C(n927), .Y(n931) );
  OAI22X1 U1161 ( .A(n97), .B(n944), .C(n470), .D(n186), .Y(n930) );
  OAI21X1 U1162 ( .A(n931), .B(n930), .C(n61), .Y(n933) );
  NAND2X1 U1163 ( .A(n965), .B(n1367), .Y(n932) );
  NAND3X1 U1164 ( .A(n936), .B(n933), .C(n932), .Y(n938) );
  MUX2X1 U1165 ( .B(n938), .A(n222), .S(n937), .Y(n939) );
  NAND2X1 U1166 ( .A(n940), .B(n939), .Y(n1290) );
  AOI22X1 U1167 ( .A(currentPlainKey[43]), .B(n205), .C(n221), .D(n1460), .Y(
        n954) );
  NAND2X1 U1168 ( .A(n1367), .B(n1459), .Y(n950) );
  NOR2X1 U1169 ( .A(n470), .B(n183), .Y(n943) );
  OAI22X1 U1170 ( .A(n187), .B(n955), .C(n502), .D(n957), .Y(n942) );
  OAI21X1 U1171 ( .A(n943), .B(n942), .C(n981), .Y(n947) );
  INVX2 U1172 ( .A(n944), .Y(n998) );
  NAND2X1 U1173 ( .A(n998), .B(n195), .Y(n945) );
  NAND3X1 U1174 ( .A(n950), .B(n947), .C(n945), .Y(n951) );
  NAND2X1 U1175 ( .A(n61), .B(n951), .Y(n953) );
  NAND2X1 U1176 ( .A(n965), .B(n217), .Y(n952) );
  NAND3X1 U1177 ( .A(n954), .B(n953), .C(n952), .Y(n1289) );
  AOI22X1 U1178 ( .A(currentPlainKey[44]), .B(n205), .C(n210), .D(n1459), .Y(
        n969) );
  NAND2X1 U1179 ( .A(n195), .B(n1458), .Y(n964) );
  OAI22X1 U1180 ( .A(n97), .B(n955), .C(n442), .D(n185), .Y(n959) );
  NAND2X1 U1181 ( .A(n105), .B(n20), .Y(n1007) );
  NAND2X1 U1188 ( .A(n442), .B(n1007), .Y(n987) );
  INVX2 U1191 ( .A(n987), .Y(n1042) );
  NAND2X1 U1192 ( .A(n490), .B(n1042), .Y(n956) );
  OAI22X1 U1193 ( .A(n154), .B(n1007), .C(n957), .D(n956), .Y(n958) );
  OAI21X1 U1194 ( .A(n959), .B(n958), .C(n981), .Y(n963) );
  NAND2X1 U1195 ( .A(n998), .B(n1367), .Y(n960) );
  NAND3X1 U1196 ( .A(n964), .B(n963), .C(n960), .Y(n966) );
  MUX2X1 U1197 ( .B(n966), .A(n222), .S(n965), .Y(n967) );
  NAND2X1 U1198 ( .A(n969), .B(n967), .Y(n1288) );
  NAND2X1 U1200 ( .A(n998), .B(n210), .Y(n985) );
  NAND2X1 U1201 ( .A(n1026), .B(n193), .Y(n979) );
  NOR2X1 U1202 ( .A(n442), .B(n183), .Y(n974) );
  INVX2 U1203 ( .A(n475), .Y(n970) );
  NAND3X1 U1204 ( .A(n1042), .B(n87), .C(n970), .Y(n971) );
  OAI21X1 U1205 ( .A(n185), .B(n1007), .C(n971), .Y(n972) );
  OAI21X1 U1206 ( .A(n974), .B(n972), .C(n43), .Y(n978) );
  NAND2X1 U1207 ( .A(n1367), .B(n1458), .Y(n977) );
  NAND3X1 U1208 ( .A(n979), .B(n978), .C(n977), .Y(n980) );
  NAND2X1 U1209 ( .A(n981), .B(n980), .Y(n984) );
  AND2X2 U1210 ( .A(currentPlainKey[45]), .B(n206), .Y(n982) );
  AOI21X1 U1211 ( .A(n221), .B(n1459), .C(n982), .Y(n983) );
  NAND3X1 U1212 ( .A(n985), .B(n984), .C(n983), .Y(n1287) );
  AOI22X1 U1213 ( .A(currentPlainKey[46]), .B(n206), .C(n210), .D(n1458), .Y(
        n1001) );
  NAND2X1 U1214 ( .A(n195), .B(n1457), .Y(n997) );
  NAND2X1 U1215 ( .A(n31), .B(n105), .Y(n1016) );
  INVX2 U1216 ( .A(n1016), .Y(n1084) );
  NAND2X1 U1217 ( .A(n1084), .B(n1136), .Y(n992) );
  NAND2X1 U1218 ( .A(n41), .B(n87), .Y(n1020) );
  INVX2 U1219 ( .A(n1020), .Y(n986) );
  NAND2X1 U1221 ( .A(n463), .B(n986), .Y(n991) );
  AOI21X1 U1222 ( .A(n992), .B(n991), .C(n987), .Y(n994) );
  OAI22X1 U1223 ( .A(n180), .B(n1007), .C(n410), .D(n185), .Y(n993) );
  OAI21X1 U1224 ( .A(n994), .B(n993), .C(n43), .Y(n996) );
  NAND2X1 U1225 ( .A(n1026), .B(n1367), .Y(n995) );
  NAND3X1 U1226 ( .A(n997), .B(n996), .C(n995), .Y(n999) );
  MUX2X1 U1227 ( .B(n999), .A(n222), .S(n998), .Y(n1000) );
  NAND2X1 U1228 ( .A(n1001), .B(n1000), .Y(n1286) );
  AOI22X1 U1229 ( .A(currentPlainKey[47]), .B(n206), .C(n219), .D(n1458), .Y(
        n1015) );
  NAND2X1 U1230 ( .A(n1367), .B(n1457), .Y(n1010) );
  NOR2X1 U1231 ( .A(n410), .B(n183), .Y(n1005) );
  OAI22X1 U1232 ( .A(n187), .B(n1016), .C(n447), .D(n1020), .Y(n1003) );
  OAI21X1 U1233 ( .A(n1005), .B(n1003), .C(n1042), .Y(n1009) );
  INVX2 U1234 ( .A(n1007), .Y(n1058) );
  NAND2X1 U1235 ( .A(n1058), .B(n193), .Y(n1008) );
  NAND3X1 U1236 ( .A(n1010), .B(n1009), .C(n1008), .Y(n1012) );
  NAND2X1 U1237 ( .A(n43), .B(n1012), .Y(n1014) );
  NAND2X1 U1238 ( .A(n1026), .B(n1363), .Y(n1013) );
  NAND3X1 U1239 ( .A(n1015), .B(n1014), .C(n1013), .Y(n1285) );
  AOI22X1 U1240 ( .A(currentPlainKey[48]), .B(n205), .C(n210), .D(n1457), .Y(
        n1029) );
  NAND2X1 U1241 ( .A(n195), .B(n1456), .Y(n1025) );
  OAI22X1 U1242 ( .A(n180), .B(n1016), .C(n379), .D(n185), .Y(n1022) );
  NAND2X1 U1243 ( .A(n105), .B(n35), .Y(n1066) );
  NAND2X1 U1244 ( .A(n379), .B(n1066), .Y(n1050) );
  INVX2 U1245 ( .A(n1050), .Y(n1098) );
  NAND2X1 U1246 ( .A(n433), .B(n1098), .Y(n1017) );
  OAI22X1 U1247 ( .A(n154), .B(n1066), .C(n1020), .D(n1017), .Y(n1021) );
  OAI21X1 U1248 ( .A(n1022), .B(n1021), .C(n1042), .Y(n1024) );
  NAND2X1 U1249 ( .A(n1058), .B(n1367), .Y(n1023) );
  NAND3X1 U1250 ( .A(n1025), .B(n1024), .C(n1023), .Y(n1027) );
  MUX2X1 U1251 ( .B(n1027), .A(n222), .S(n1026), .Y(n1028) );
  NAND2X1 U1252 ( .A(n1029), .B(n1028), .Y(n1284) );
  NAND2X1 U1253 ( .A(n1058), .B(n210), .Y(n1048) );
  NAND2X1 U1254 ( .A(n1084), .B(n193), .Y(n1040) );
  NOR2X1 U1255 ( .A(n379), .B(n183), .Y(n1036) );
  INVX2 U1256 ( .A(n415), .Y(n1030) );
  NAND3X1 U1257 ( .A(n1098), .B(n87), .C(n1030), .Y(n1032) );
  OAI21X1 U1258 ( .A(n186), .B(n1066), .C(n1032), .Y(n1035) );
  OAI21X1 U1259 ( .A(n1036), .B(n1035), .C(n41), .Y(n1039) );
  NAND2X1 U1260 ( .A(n1367), .B(n1456), .Y(n1037) );
  NAND3X1 U1261 ( .A(n1040), .B(n1039), .C(n1037), .Y(n1041) );
  NAND2X1 U1262 ( .A(n1042), .B(n1041), .Y(n1045) );
  AND2X2 U1263 ( .A(currentPlainKey[49]), .B(n207), .Y(n1043) );
  AOI21X1 U1264 ( .A(n221), .B(n1457), .C(n1043), .Y(n1044) );
  NAND3X1 U1265 ( .A(n1048), .B(n1045), .C(n1044), .Y(n1283) );
  AOI22X1 U1266 ( .A(currentPlainKey[50]), .B(n206), .C(n209), .D(n1456), .Y(
        n1061) );
  NAND2X1 U1267 ( .A(n197), .B(n1455), .Y(n1057) );
  NAND2X1 U1268 ( .A(n11), .B(n143), .Y(n1074) );
  INVX2 U1269 ( .A(n1074), .Y(n1146) );
  NAND2X1 U1270 ( .A(n1146), .B(n1136), .Y(n1052) );
  NAND2X1 U1271 ( .A(n63), .B(n87), .Y(n1076) );
  INVX2 U1272 ( .A(n1076), .Y(n1049) );
  NAND2X1 U1275 ( .A(n401), .B(n1049), .Y(n1051) );
  AOI21X1 U1276 ( .A(n1052), .B(n1051), .C(n1050), .Y(n1054) );
  OAI22X1 U1277 ( .A(n97), .B(n1066), .C(n349), .D(n185), .Y(n1053) );
  OAI21X1 U1278 ( .A(n1054), .B(n1053), .C(n41), .Y(n1056) );
  NAND2X1 U1279 ( .A(n1084), .B(n1367), .Y(n1055) );
  NAND3X1 U1280 ( .A(n1057), .B(n1056), .C(n1055), .Y(n1059) );
  MUX2X1 U1281 ( .B(n1059), .A(n222), .S(n1058), .Y(n1060) );
  NAND2X1 U1282 ( .A(n1061), .B(n1060), .Y(n1282) );
  AOI22X1 U1283 ( .A(currentPlainKey[51]), .B(n205), .C(n219), .D(n1456), .Y(
        n1073) );
  NAND2X1 U1284 ( .A(n1367), .B(n1455), .Y(n1069) );
  NOR2X1 U1285 ( .A(n349), .B(n183), .Y(n1065) );
  OAI22X1 U1286 ( .A(n187), .B(n1074), .C(n384), .D(n1076), .Y(n1064) );
  OAI21X1 U1287 ( .A(n1065), .B(n1064), .C(n1098), .Y(n1068) );
  INVX2 U1288 ( .A(n1066), .Y(n1118) );
  NAND2X1 U1289 ( .A(n1118), .B(n193), .Y(n1067) );
  NAND3X1 U1290 ( .A(n1069), .B(n1068), .C(n1067), .Y(n1070) );
  NAND2X1 U1291 ( .A(n41), .B(n1070), .Y(n1072) );
  NAND2X1 U1292 ( .A(n1084), .B(n217), .Y(n1071) );
  NAND3X1 U1293 ( .A(n1073), .B(n1072), .C(n1071), .Y(n1281) );
  AOI22X1 U1294 ( .A(currentPlainKey[52]), .B(n205), .C(n209), .D(n1455), .Y(
        n1087) );
  NAND2X1 U1295 ( .A(n195), .B(n1454), .Y(n1083) );
  OAI22X1 U1296 ( .A(n180), .B(n1074), .C(n318), .D(n185), .Y(n1080) );
  NAND2X1 U1297 ( .A(n11), .B(n1481), .Y(n1122) );
  NAND2X1 U1298 ( .A(n318), .B(n1122), .Y(n1110) );
  INVX2 U1299 ( .A(n1110), .Y(n1157) );
  NAND2X1 U1300 ( .A(n371), .B(n1157), .Y(n1075) );
  OAI22X1 U1301 ( .A(n1122), .B(n153), .C(n1076), .D(n1075), .Y(n1079) );
  OAI21X1 U1302 ( .A(n1080), .B(n1079), .C(n1098), .Y(n1082) );
  NAND2X1 U1303 ( .A(n1118), .B(n1367), .Y(n1081) );
  NAND3X1 U1304 ( .A(n1083), .B(n1082), .C(n1081), .Y(n1085) );
  MUX2X1 U1306 ( .B(n1085), .A(n222), .S(n1084), .Y(n1086) );
  NAND2X1 U1307 ( .A(n1087), .B(n1086), .Y(n1280) );
  NAND2X1 U1308 ( .A(n1118), .B(n209), .Y(n1109) );
  NAND2X1 U1309 ( .A(n1146), .B(n193), .Y(n1096) );
  NOR2X1 U1310 ( .A(n318), .B(n183), .Y(n1093) );
  INVX2 U1311 ( .A(n354), .Y(n1088) );
  NAND3X1 U1312 ( .A(n1157), .B(n175), .C(n1088), .Y(n1091) );
  OAI21X1 U1313 ( .A(n185), .B(n1122), .C(n1091), .Y(n1092) );
  OAI21X1 U1316 ( .A(n1093), .B(n1092), .C(n63), .Y(n1095) );
  NAND2X1 U1317 ( .A(n1367), .B(n1454), .Y(n1094) );
  NAND3X1 U1318 ( .A(n1096), .B(n1095), .C(n1094), .Y(n1097) );
  NAND2X1 U1319 ( .A(n1098), .B(n1097), .Y(n1102) );
  AND2X2 U1320 ( .A(currentPlainKey[53]), .B(n205), .Y(n1099) );
  AOI21X1 U1321 ( .A(n221), .B(n1455), .C(n1099), .Y(n1100) );
  NAND3X1 U1322 ( .A(n1109), .B(n1102), .C(n1100), .Y(n1279) );
  AOI22X1 U1323 ( .A(currentPlainKey[54]), .B(n207), .C(n209), .D(n1454), .Y(
        n1121) );
  NAND2X1 U1324 ( .A(n195), .B(n1453), .Y(n1117) );
  NAND2X1 U1325 ( .A(n11), .B(n1478), .Y(n1125) );
  NAND2X1 U1326 ( .A(n283), .B(n1125), .Y(n1138) );
  INVX2 U1327 ( .A(n1138), .Y(n1177) );
  NAND3X1 U1328 ( .A(n341), .B(n87), .C(n1177), .Y(n1112) );
  INVX2 U1329 ( .A(n1125), .Y(n1193) );
  NAND2X1 U1330 ( .A(n1136), .B(n1193), .Y(n1111) );
  AOI21X1 U1331 ( .A(n1112), .B(n1111), .C(n1110), .Y(n1114) );
  OAI22X1 U1332 ( .A(n283), .B(n137), .C(n97), .D(n1122), .Y(n1113) );
  OAI21X1 U1333 ( .A(n1114), .B(n1113), .C(n63), .Y(n1116) );
  NAND2X1 U1334 ( .A(n1146), .B(n1367), .Y(n1115) );
  NAND3X1 U1335 ( .A(n1117), .B(n1116), .C(n1115), .Y(n1119) );
  MUX2X1 U1336 ( .B(n1119), .A(n222), .S(n1118), .Y(n1120) );
  NAND2X1 U1337 ( .A(n1121), .B(n1120), .Y(n1278) );
  NAND2X1 U1338 ( .A(n1146), .B(n209), .Y(n1135) );
  INVX2 U1339 ( .A(n1122), .Y(n1168) );
  NAND2X1 U1340 ( .A(n1168), .B(n192), .Y(n1130) );
  NOR2X1 U1341 ( .A(n283), .B(n183), .Y(n1127) );
  INVX2 U1342 ( .A(n323), .Y(n1123) );
  NAND3X1 U1343 ( .A(n1177), .B(n175), .C(n1123), .Y(n1124) );
  OAI21X1 U1344 ( .A(n1125), .B(n137), .C(n1124), .Y(n1126) );
  OAI21X1 U1345 ( .A(n1127), .B(n1126), .C(n1157), .Y(n1129) );
  NAND2X1 U1346 ( .A(n1367), .B(n1453), .Y(n1128) );
  NAND3X1 U1347 ( .A(n1130), .B(n1129), .C(n1128), .Y(n1131) );
  NAND2X1 U1348 ( .A(n63), .B(n1131), .Y(n1134) );
  AND2X2 U1349 ( .A(currentPlainKey[55]), .B(n207), .Y(n1132) );
  AOI21X1 U1350 ( .A(n221), .B(n1454), .C(n1132), .Y(n1133) );
  NAND3X1 U1351 ( .A(n1135), .B(n1134), .C(n1133), .Y(n1277) );
  AOI22X1 U1352 ( .A(currentPlainKey[56]), .B(n206), .C(n209), .D(n1453), .Y(
        n1149) );
  NAND2X1 U1353 ( .A(n195), .B(n1452), .Y(n1145) );
  NAND2X1 U1354 ( .A(n11), .B(n16), .Y(n1173) );
  NAND3X1 U1355 ( .A(n87), .B(n1173), .C(n246), .Y(n1150) );
  INVX2 U1356 ( .A(n1150), .Y(n1263) );
  INVX2 U1357 ( .A(n1173), .Y(n1357) );
  AOI22X1 U1358 ( .A(n306), .B(n1263), .C(n1136), .D(n1357), .Y(n1139) );
  AOI22X1 U1359 ( .A(n184), .B(n1193), .C(n188), .D(n1451), .Y(n1137) );
  OAI21X1 U1360 ( .A(n1139), .B(n1138), .C(n1137), .Y(n1140) );
  NAND2X1 U1361 ( .A(n1157), .B(n1140), .Y(n1142) );
  NAND2X1 U1362 ( .A(n1168), .B(n1367), .Y(n1141) );
  NAND3X1 U1363 ( .A(n1145), .B(n1142), .C(n1141), .Y(n1147) );
  MUX2X1 U1364 ( .B(n1147), .A(n222), .S(n1146), .Y(n1148) );
  NAND2X1 U1365 ( .A(n1149), .B(n1148), .Y(n1276) );
  AOI22X1 U1366 ( .A(currentPlainKey[57]), .B(n206), .C(n219), .D(n1453), .Y(
        n1161) );
  NAND2X1 U1367 ( .A(n1367), .B(n1452), .Y(n1155) );
  NOR2X1 U1368 ( .A(n288), .B(n1150), .Y(n1152) );
  OAI22X1 U1369 ( .A(n246), .B(n97), .C(n1173), .D(n185), .Y(n1151) );
  OAI21X1 U1370 ( .A(n1152), .B(n1151), .C(n1177), .Y(n1154) );
  NAND2X1 U1371 ( .A(n1193), .B(n192), .Y(n1153) );
  NAND3X1 U1372 ( .A(n1155), .B(n1154), .C(n1153), .Y(n1156) );
  NAND2X1 U1373 ( .A(n1157), .B(n1156), .Y(n1159) );
  NAND2X1 U1374 ( .A(n1168), .B(n210), .Y(n1158) );
  NAND3X1 U1375 ( .A(n1161), .B(n1159), .C(n1158), .Y(n1275) );
  AOI22X1 U1376 ( .A(currentPlainKey[58]), .B(n205), .C(n209), .D(n1452), .Y(
        n1171) );
  NAND2X1 U1377 ( .A(n195), .B(n1451), .Y(n1167) );
  NAND2X1 U1378 ( .A(n1263), .B(n152), .Y(n1187) );
  INVX2 U1379 ( .A(n272), .Y(n1162) );
  OAI22X1 U1380 ( .A(n152), .B(n137), .C(n1173), .D(n180), .Y(n1163) );
  OAI21X1 U1381 ( .A(n1164), .B(n1163), .C(n1177), .Y(n1166) );
  NAND2X1 U1382 ( .A(n1193), .B(n1367), .Y(n1165) );
  NAND3X1 U1383 ( .A(n1167), .B(n1166), .C(n1165), .Y(n1169) );
  MUX2X1 U1384 ( .B(n1169), .A(n222), .S(n1168), .Y(n1170) );
  NAND2X1 U1385 ( .A(n1171), .B(n1170), .Y(n1274) );
  AOI22X1 U1386 ( .A(currentPlainKey[59]), .B(n205), .C(n219), .D(n1452), .Y(
        n1183) );
  OAI22X1 U1387 ( .A(n246), .B(n4), .C(n1173), .D(n1172), .Y(n1180) );
  INVX2 U1388 ( .A(n251), .Y(n1176) );
  NAND3X1 U1389 ( .A(RCV_DATA[3]), .B(n1450), .C(n1263), .Y(n1175) );
  OAI21X1 U1390 ( .A(n1187), .B(n1176), .C(n1175), .Y(n1179) );
  OAI21X1 U1391 ( .A(n1180), .B(n1179), .C(n1177), .Y(n1182) );
  NAND2X1 U1392 ( .A(n1193), .B(n210), .Y(n1181) );
  NAND3X1 U1393 ( .A(n1183), .B(n1182), .C(n1181), .Y(n1273) );
  AOI22X1 U1394 ( .A(currentPlainKey[60]), .B(n207), .C(n209), .D(n1451), .Y(
        n1196) );
  NAND2X1 U1395 ( .A(n197), .B(n1450), .Y(n1192) );
  AOI22X1 U1396 ( .A(n1497), .B(RCV_DATA[3]), .C(n1449), .D(RCV_DATA[2]), .Y(
        n1185) );
  OAI21X1 U1397 ( .A(n226), .B(n164), .C(n1185), .Y(n1189) );
  INVX2 U1398 ( .A(n1187), .Y(n1188) );
  OAI21X1 U1399 ( .A(n67), .B(n1189), .C(n1188), .Y(n1191) );
  NAND2X1 U1400 ( .A(n1367), .B(n1357), .Y(n1190) );
  NAND3X1 U1401 ( .A(n1192), .B(n1191), .C(n1190), .Y(n1194) );
  MUX2X1 U1402 ( .B(n1194), .A(n222), .S(n1193), .Y(n1195) );
  NAND2X1 U1403 ( .A(n1196), .B(n1195), .Y(n1272) );
  AOI22X1 U1404 ( .A(currentPlainKey[61]), .B(n207), .C(n219), .D(n1451), .Y(
        n1266) );
  NAND2X1 U1405 ( .A(n1450), .B(RCV_DATA[5]), .Y(n1261) );
  NAND2X1 U1406 ( .A(n211), .B(n1261), .Y(n1262) );
  NAND2X1 U1407 ( .A(n1263), .B(n1262), .Y(n1265) );
  NAND2X1 U1408 ( .A(n1357), .B(n1363), .Y(n1264) );
  NAND3X1 U1409 ( .A(n1266), .B(n1265), .C(n1264), .Y(n1271) );
  AND2X2 U1410 ( .A(n207), .B(currentPlainKey[62]), .Y(n1267) );
  AOI21X1 U1411 ( .A(n217), .B(n1450), .C(n1267), .Y(n1362) );
  NOR2X1 U1412 ( .A(n1450), .B(n1364), .Y(n1268) );
  OAI21X1 U1413 ( .A(n190), .B(n191), .C(n1268), .Y(n1359) );
  MUX2X1 U1414 ( .B(n1359), .A(n1358), .S(n1357), .Y(n1360) );
  INVX2 U1415 ( .A(n1360), .Y(n1361) );
  NAND2X1 U1416 ( .A(n1362), .B(n1361), .Y(n1270) );
  NAND2X1 U1417 ( .A(n207), .B(currentPlainKey[63]), .Y(n1373) );
  NAND2X1 U1418 ( .A(n210), .B(n1497), .Y(n1369) );
  NOR2X1 U1419 ( .A(n1449), .B(n1364), .Y(n1366) );
  INVX2 U1420 ( .A(n155), .Y(n1365) );
  OAI21X1 U1421 ( .A(n1367), .B(n1366), .C(n1365), .Y(n1368) );
  NAND2X1 U1422 ( .A(n1369), .B(n1368), .Y(n1371) );
  MUX2X1 U1423 ( .B(n1371), .A(n223), .S(n1450), .Y(n1372) );
  NAND2X1 U1424 ( .A(n1373), .B(n1372), .Y(n1269) );
  NAND2X1 U1425 ( .A(n1374), .B(n1419), .Y(n1385) );
  INVX2 U1426 ( .A(n1385), .Y(n1375) );
  NAND3X1 U1427 ( .A(n1375), .B(n242), .C(n1431), .Y(n1383) );
  INVX2 U1428 ( .A(n1383), .Y(n1381) );
  NAND2X1 U1429 ( .A(n1381), .B(keyCount[3]), .Y(n1384) );
  NAND2X1 U1430 ( .A(address[0]), .B(n1383), .Y(n1376) );
  NAND2X1 U1431 ( .A(n1384), .B(n1376), .Y(n1333) );
  NAND2X1 U1432 ( .A(address[1]), .B(n1383), .Y(n1377) );
  NAND2X1 U1433 ( .A(n1384), .B(n1377), .Y(n1334) );
  NAND2X1 U1434 ( .A(address[2]), .B(n1383), .Y(n1378) );
  NAND2X1 U1435 ( .A(n1384), .B(n1378), .Y(n1335) );
  MUX2X1 U1436 ( .B(address[3]), .A(keyCount[0]), .S(n1381), .Y(n1379) );
  NAND2X1 U1437 ( .A(n1384), .B(n1379), .Y(n1336) );
  MUX2X1 U1438 ( .B(address[4]), .A(keyCount[1]), .S(n1381), .Y(n1380) );
  NAND2X1 U1439 ( .A(n1384), .B(n1380), .Y(n1337) );
  MUX2X1 U1440 ( .B(address[5]), .A(keyCount[2]), .S(n1381), .Y(n1382) );
  NAND2X1 U1441 ( .A(n1384), .B(n1382), .Y(n1338) );
  OAI21X1 U1442 ( .A(n1503), .B(n1381), .C(n1384), .Y(n1339) );
  OAI21X1 U1443 ( .A(n1495), .B(n1381), .C(n1384), .Y(n1340) );
  OAI21X1 U1444 ( .A(n1386), .B(n1385), .C(parityError), .Y(n1389) );
  OAI21X1 U1445 ( .A(n12), .B(n13), .C(n1387), .Y(n1388) );
  NAND2X1 U1446 ( .A(n1389), .B(n1388), .Y(nextParityError) );
  NOR2X1 U1447 ( .A(keyCount[0]), .B(n1442), .Y(n1390) );
  NOR2X1 U1448 ( .A(n1390), .B(n1446), .Y(n1393) );
  INVX2 U1449 ( .A(n1448), .Y(n1391) );
  NAND2X1 U1450 ( .A(keyCount[0]), .B(n1391), .Y(n1392) );
  MUX2X1 U1451 ( .B(n1393), .A(n1392), .S(n1494), .Y(n1350) );
  NAND2X1 U1452 ( .A(n1399), .B(CLR_RBUFF), .Y(n1411) );
  INVX2 U1453 ( .A(n1411), .Y(n1404) );
  NAND2X1 U1454 ( .A(N1799), .B(n1404), .Y(n1394) );
  OAI21X1 U1455 ( .A(n1493), .B(n1395), .C(n1394), .Y(n1341) );
  NAND2X1 U1456 ( .A(N1798), .B(n1404), .Y(n1396) );
  OAI21X1 U1457 ( .A(n1492), .B(n1397), .C(n1396), .Y(n1342) );
  NAND2X1 U1458 ( .A(N1797), .B(n1404), .Y(n1398) );
  OAI21X1 U1459 ( .A(n1491), .B(n1399), .C(n1398), .Y(n1343) );
  NAND2X1 U1460 ( .A(N1796), .B(n1404), .Y(n1400) );
  OAI21X1 U1461 ( .A(n1490), .B(n1401), .C(n1400), .Y(n1344) );
  NAND2X1 U1462 ( .A(N1795), .B(n1404), .Y(n1402) );
  OAI21X1 U1463 ( .A(n1489), .B(n1403), .C(n1402), .Y(n1345) );
  NAND2X1 U1464 ( .A(N1794), .B(n1404), .Y(n1405) );
  OAI21X1 U1465 ( .A(n1488), .B(n1406), .C(n1405), .Y(n1346) );
  INVX2 U1466 ( .A(N1793), .Y(n1407) );
  OAI22X1 U1467 ( .A(n1487), .B(n1408), .C(n1411), .D(n1407), .Y(n1347) );
  INVX2 U1468 ( .A(N1792), .Y(n1410) );
  OAI22X1 U1469 ( .A(n1486), .B(n1408), .C(n1411), .D(n1410), .Y(n1348) );
  AOI21X1 U1470 ( .A(N694), .B(RBUF_FULL), .C(n1178), .Y(n1412) );
  NAND2X1 U1471 ( .A(n1412), .B(n83), .Y(n1415) );
  NAND2X1 U1472 ( .A(n1413), .B(n89), .Y(n1414) );
  NAND2X1 U1473 ( .A(n1414), .B(n1429), .Y(n1436) );
  NAND2X1 U1474 ( .A(n1415), .B(n1436), .Y(n1426) );
  INVX2 U1475 ( .A(n1426), .Y(n1418) );
  OAI21X1 U1476 ( .A(n1418), .B(n89), .C(n1416), .Y(n1354) );
  OAI21X1 U1477 ( .A(OE), .B(SBE), .C(n83), .Y(n1422) );
  OAI22X1 U1478 ( .A(RBUF_FULL), .B(n1419), .C(n131), .D(n1436), .Y(n1420) );
  AOI21X1 U1479 ( .A(n1425), .B(n1437), .C(n1420), .Y(n1421) );
  NAND3X1 U1480 ( .A(n1423), .B(n1422), .C(n1421), .Y(n1352) );
  AOI21X1 U1481 ( .A(state[1]), .B(n1426), .C(n1425), .Y(n1427) );
  NAND2X1 U1482 ( .A(n127), .B(n1427), .Y(n1351) );
  INVX2 U1483 ( .A(RBUF_FULL), .Y(n1428) );
  AOI21X1 U1484 ( .A(n1430), .B(n1429), .C(n1428), .Y(n1435) );
  NAND2X1 U1485 ( .A(n1574), .B(n1579), .Y(n1433) );
  OAI21X1 U1486 ( .A(n1433), .B(n1432), .C(n93), .Y(n1434) );
  NOR2X1 U1487 ( .A(n1435), .B(n1434), .Y(n1441) );
  INVX2 U1488 ( .A(n1160), .Y(n1437) );
  OAI22X1 U1489 ( .A(n1442), .B(n1437), .C(n139), .D(n1436), .Y(n1438) );
  NOR2X1 U1490 ( .A(n1439), .B(n1438), .Y(n1440) );
  NAND2X1 U1491 ( .A(n1441), .B(n1440), .Y(n1353) );
  NOR2X1 U1492 ( .A(keyCount[2]), .B(n1442), .Y(n1444) );
  OAI21X1 U1493 ( .A(n1444), .B(n1443), .C(keyCount[3]), .Y(n1445) );
  OAI21X1 U1494 ( .A(n1160), .B(n1448), .C(n1445), .Y(n1355) );
  NAND2X1 U1495 ( .A(n1446), .B(keyCount[0]), .Y(n1447) );
  OAI21X1 U1496 ( .A(keyCount[0]), .B(n1448), .C(n1447), .Y(n1356) );
  INVX2 U1497 ( .A(keyCount[3]), .Y(N694) );
  INVX2 U1498 ( .A(keyCount[0]), .Y(n1483) );
  INVX2 U1499 ( .A(keyCount[2]), .Y(n1484) );
  INVX2 U1500 ( .A(parityAccumulator[0]), .Y(n1486) );
  INVX2 U1501 ( .A(parityAccumulator[1]), .Y(n1487) );
  INVX2 U1502 ( .A(parityAccumulator[2]), .Y(n1488) );
  INVX2 U1503 ( .A(parityAccumulator[3]), .Y(n1489) );
  INVX2 U1504 ( .A(parityAccumulator[4]), .Y(n1490) );
  INVX2 U1505 ( .A(parityAccumulator[5]), .Y(n1491) );
  INVX2 U1506 ( .A(parityAccumulator[6]), .Y(n1492) );
  INVX2 U1507 ( .A(parityAccumulator[7]), .Y(n1493) );
  INVX2 U1508 ( .A(keyCount[1]), .Y(n1494) );
  INVX2 U1509 ( .A(address[7]), .Y(n1495) );
  INVX2 U1510 ( .A(n204), .Y(n1496) );
  INVX2 U1511 ( .A(n157), .Y(n1497) );
  INVX2 U1512 ( .A(n164), .Y(n1498) );
  INVX2 U1513 ( .A(n167), .Y(n1499) );
  INVX2 U1514 ( .A(n171), .Y(n1500) );
  INVX2 U1515 ( .A(n176), .Y(n1501) );
  INVX2 U1516 ( .A(address[6]), .Y(n1503) );
  INVX2 U1517 ( .A(n274), .Y(n1504) );
  INVX2 U1518 ( .A(n254), .Y(n1505) );
  INVX2 U1519 ( .A(n218), .Y(n1506) );
  INVX2 U1520 ( .A(n179), .Y(n1507) );
  INVX2 U1521 ( .A(address[5]), .Y(n1508) );
  INVX2 U1522 ( .A(address[4]), .Y(n1509) );
  INVX2 U1523 ( .A(currentPlainKey[63]), .Y(n1510) );
  INVX2 U1524 ( .A(currentPlainKey[62]), .Y(n1511) );
  INVX2 U1525 ( .A(currentPlainKey[61]), .Y(n1512) );
  INVX2 U1526 ( .A(currentPlainKey[60]), .Y(n1513) );
  INVX2 U1527 ( .A(currentPlainKey[59]), .Y(n1514) );
  INVX2 U1528 ( .A(currentPlainKey[58]), .Y(n1515) );
  INVX2 U1529 ( .A(currentPlainKey[57]), .Y(n1516) );
  INVX2 U1530 ( .A(currentPlainKey[56]), .Y(n1517) );
  INVX2 U1531 ( .A(currentPlainKey[55]), .Y(n1518) );
  INVX2 U1532 ( .A(currentPlainKey[54]), .Y(n1519) );
  INVX2 U1533 ( .A(currentPlainKey[53]), .Y(n1520) );
  INVX2 U1534 ( .A(currentPlainKey[52]), .Y(n1521) );
  INVX2 U1535 ( .A(currentPlainKey[51]), .Y(n1522) );
  INVX2 U1536 ( .A(currentPlainKey[50]), .Y(n1523) );
  INVX2 U1537 ( .A(currentPlainKey[49]), .Y(n1524) );
  INVX2 U1538 ( .A(currentPlainKey[48]), .Y(n1525) );
  INVX2 U1539 ( .A(currentPlainKey[47]), .Y(n1526) );
  INVX2 U1540 ( .A(currentPlainKey[46]), .Y(n1527) );
  INVX2 U1541 ( .A(currentPlainKey[45]), .Y(n1528) );
  INVX2 U1542 ( .A(currentPlainKey[44]), .Y(n1529) );
  INVX2 U1543 ( .A(currentPlainKey[43]), .Y(n1530) );
  INVX2 U1544 ( .A(currentPlainKey[42]), .Y(n1531) );
  INVX2 U1545 ( .A(currentPlainKey[41]), .Y(n1532) );
  INVX2 U1546 ( .A(currentPlainKey[40]), .Y(n1533) );
  INVX2 U1547 ( .A(currentPlainKey[39]), .Y(n1534) );
  INVX2 U1548 ( .A(currentPlainKey[38]), .Y(n1535) );
  INVX2 U1549 ( .A(currentPlainKey[37]), .Y(n1536) );
  INVX2 U1550 ( .A(currentPlainKey[36]), .Y(n1537) );
  INVX2 U1551 ( .A(currentPlainKey[35]), .Y(n1538) );
  INVX2 U1552 ( .A(currentPlainKey[34]), .Y(n1539) );
  INVX2 U1553 ( .A(currentPlainKey[33]), .Y(n1540) );
  INVX2 U1554 ( .A(currentPlainKey[32]), .Y(n1541) );
  INVX2 U1555 ( .A(currentPlainKey[31]), .Y(n1542) );
  INVX2 U1556 ( .A(currentPlainKey[30]), .Y(n1543) );
  INVX2 U1557 ( .A(currentPlainKey[29]), .Y(n1544) );
  INVX2 U1558 ( .A(currentPlainKey[28]), .Y(n1545) );
  INVX2 U1559 ( .A(currentPlainKey[27]), .Y(n1546) );
  INVX2 U1560 ( .A(currentPlainKey[26]), .Y(n1547) );
  INVX2 U1561 ( .A(currentPlainKey[25]), .Y(n1548) );
  INVX2 U1562 ( .A(currentPlainKey[24]), .Y(n1549) );
  INVX2 U1563 ( .A(currentPlainKey[23]), .Y(n1550) );
  INVX2 U1564 ( .A(currentPlainKey[22]), .Y(n1551) );
  INVX2 U1565 ( .A(currentPlainKey[21]), .Y(n1552) );
  INVX2 U1566 ( .A(currentPlainKey[20]), .Y(n1553) );
  INVX2 U1567 ( .A(currentPlainKey[19]), .Y(n1554) );
  INVX2 U1568 ( .A(currentPlainKey[18]), .Y(n1555) );
  INVX2 U1569 ( .A(currentPlainKey[17]), .Y(n1556) );
  INVX2 U1570 ( .A(currentPlainKey[16]), .Y(n1557) );
  INVX2 U1571 ( .A(currentPlainKey[15]), .Y(n1558) );
  INVX2 U1572 ( .A(currentPlainKey[14]), .Y(n1559) );
  INVX2 U1573 ( .A(currentPlainKey[13]), .Y(n1560) );
  INVX2 U1574 ( .A(currentPlainKey[12]), .Y(n1561) );
  INVX2 U1575 ( .A(currentPlainKey[11]), .Y(n1562) );
  INVX2 U1576 ( .A(currentPlainKey[10]), .Y(n1563) );
  INVX2 U1577 ( .A(currentPlainKey[9]), .Y(n1564) );
  INVX2 U1578 ( .A(currentPlainKey[8]), .Y(n1565) );
  INVX2 U1579 ( .A(currentPlainKey[7]), .Y(n1566) );
  INVX2 U1580 ( .A(currentPlainKey[6]), .Y(n1567) );
  INVX2 U1581 ( .A(currentPlainKey[5]), .Y(n1568) );
  INVX2 U1582 ( .A(currentPlainKey[4]), .Y(n1569) );
  INVX2 U1583 ( .A(currentPlainKey[0]), .Y(n1573) );
  INVX2 U1584 ( .A(SBE), .Y(n1574) );
  INVX2 U1585 ( .A(OE), .Y(n1579) );
endmodule


module uart_timer_1_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module uart_timer_1 ( CLK, RST, TIMER_TRIG, STOP_RCVING, SHIFT_STROBE );
  input CLK, RST, TIMER_TRIG;
  output STOP_RCVING, SHIFT_STROBE;
  wire   N26, N27, N28, N29, N30, N31, N32, N33, N60, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34;
  wire   [7:0] state;
  wire   [7:0] nextState;
  assign SHIFT_STROBE = N60;

  OR2X2 U21 ( .A(state[7]), .B(n50), .Y(n49) );
  OAI21X1 U38 ( .A(n20), .B(n27), .C(n35), .Y(n64) );
  NAND2X1 U39 ( .A(N33), .B(n36), .Y(n35) );
  OAI21X1 U40 ( .A(n26), .B(n20), .C(n37), .Y(n65) );
  NAND2X1 U41 ( .A(N32), .B(n36), .Y(n37) );
  OAI21X1 U42 ( .A(n25), .B(n20), .C(n38), .Y(n66) );
  NAND2X1 U43 ( .A(N31), .B(n36), .Y(n38) );
  OAI21X1 U44 ( .A(n20), .B(n24), .C(n39), .Y(n67) );
  NAND2X1 U45 ( .A(N30), .B(n36), .Y(n39) );
  OAI21X1 U46 ( .A(n23), .B(n20), .C(n40), .Y(n68) );
  NAND2X1 U47 ( .A(N29), .B(n36), .Y(n40) );
  OAI21X1 U48 ( .A(n22), .B(n20), .C(n41), .Y(n69) );
  NAND2X1 U49 ( .A(N28), .B(n36), .Y(n41) );
  OAI21X1 U50 ( .A(n20), .B(n21), .C(n42), .Y(n70) );
  NAND2X1 U51 ( .A(N27), .B(n36), .Y(n42) );
  OAI21X1 U52 ( .A(n19), .B(n20), .C(n43), .Y(n71) );
  NAND2X1 U53 ( .A(N26), .B(n36), .Y(n43) );
  NOR2X1 U54 ( .A(n44), .B(n72), .Y(n36) );
  NOR2X1 U55 ( .A(n72), .B(TIMER_TRIG), .Y(n44) );
  NOR2X1 U56 ( .A(n45), .B(n46), .Y(n72) );
  NAND3X1 U57 ( .A(nextState[6]), .B(nextState[5]), .C(n47), .Y(n46) );
  NOR2X1 U58 ( .A(n22), .B(n23), .Y(n47) );
  NAND3X1 U59 ( .A(nextState[0]), .B(n21), .C(n48), .Y(n45) );
  NOR2X1 U60 ( .A(nextState[7]), .B(nextState[4]), .Y(n48) );
  NOR2X1 U61 ( .A(state[0]), .B(n49), .Y(N60) );
  AOI21X1 U62 ( .A(n51), .B(n32), .C(n52), .Y(n50) );
  OAI21X1 U63 ( .A(n33), .B(n53), .C(n54), .Y(n52) );
  NAND3X1 U64 ( .A(state[6]), .B(state[1]), .C(n55), .Y(n54) );
  AOI21X1 U65 ( .A(n56), .B(n57), .C(state[3]), .Y(n55) );
  NAND3X1 U66 ( .A(n33), .B(n31), .C(state[4]), .Y(n57) );
  NAND3X1 U67 ( .A(state[2]), .B(n32), .C(state[5]), .Y(n56) );
  NAND2X1 U68 ( .A(state[4]), .B(n58), .Y(n53) );
  OAI21X1 U69 ( .A(state[2]), .B(n28), .C(n59), .Y(n51) );
  NAND3X1 U70 ( .A(state[2]), .B(n29), .C(n30), .Y(n59) );
  OAI22X1 U71 ( .A(state[6]), .B(n61), .C(n29), .D(n60), .Y(n58) );
  NAND3X1 U72 ( .A(n34), .B(n31), .C(state[3]), .Y(n60) );
  AOI22X1 U73 ( .A(n62), .B(state[1]), .C(n63), .D(state[5]), .Y(n61) );
  XOR2X1 U74 ( .A(n34), .B(state[3]), .Y(n63) );
  NOR2X1 U75 ( .A(state[5]), .B(state[3]), .Y(n62) );
  uart_timer_1_DW01_inc_0 add_39 ( .A(nextState), .SUM({N33, N32, N31, N30, 
        N29, N28, N27, N26}) );
  DFFSR \state_reg[3]  ( .D(nextState[3]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[5]  ( .D(nextState[5]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[5]) );
  DFFSR \state_reg[6]  ( .D(nextState[6]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[6]) );
  DFFSR \state_reg[4]  ( .D(nextState[4]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[7]  ( .D(nextState[7]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[7]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[0]) );
  DFFSR STOP_RCVING_reg ( .D(n72), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        STOP_RCVING) );
  DFFSR \nextState_reg[3]  ( .D(n68), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[3]) );
  DFFSR \nextState_reg[2]  ( .D(n69), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[2]) );
  DFFSR \nextState_reg[0]  ( .D(n71), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[0]) );
  DFFSR \nextState_reg[4]  ( .D(n67), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[4]) );
  DFFSR \nextState_reg[1]  ( .D(n70), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[1]) );
  DFFSR \nextState_reg[5]  ( .D(n66), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[5]) );
  DFFSR \nextState_reg[6]  ( .D(n65), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[6]) );
  DFFSR \nextState_reg[7]  ( .D(n64), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[7]) );
  INVX2 U20 ( .A(RST), .Y(n18) );
  INVX2 U22 ( .A(nextState[0]), .Y(n19) );
  INVX2 U23 ( .A(n44), .Y(n20) );
  INVX2 U24 ( .A(nextState[1]), .Y(n21) );
  INVX2 U25 ( .A(nextState[2]), .Y(n22) );
  INVX2 U26 ( .A(nextState[3]), .Y(n23) );
  INVX2 U27 ( .A(nextState[4]), .Y(n24) );
  INVX2 U28 ( .A(nextState[5]), .Y(n25) );
  INVX2 U29 ( .A(nextState[6]), .Y(n26) );
  INVX2 U30 ( .A(nextState[7]), .Y(n27) );
  INVX2 U31 ( .A(n58), .Y(n28) );
  INVX2 U32 ( .A(state[6]), .Y(n29) );
  INVX2 U33 ( .A(n60), .Y(n30) );
  INVX2 U34 ( .A(state[5]), .Y(n31) );
  INVX2 U35 ( .A(state[4]), .Y(n32) );
  INVX2 U36 ( .A(state[2]), .Y(n33) );
  INVX2 U37 ( .A(state[1]), .Y(n34) );
endmodule


module uart_rcv_block_1 ( CLK, RST, SERIAL_IN, KEY_ERROR, PROG_ERROR, PLAINKEY, 
        RBUF_FULL, PARITY_ERROR );
  output [63:0] PLAINKEY;
  input CLK, RST, SERIAL_IN;
  output KEY_ERROR, PROG_ERROR, RBUF_FULL, PARITY_ERROR;
  wire   START_BIT, CHK_ERROR, OE, SB_DETECT, STOP_RCVING, RBUF_LOAD, SBC_CLR,
         SBC_EN, SET_RBUF_FULL, TIMER_TRIG, CLR_RBUF, SBE, SHIFT_STROBE, n1,
         n2;
  wire   [7:0] LOAD_DATA;
  wire   [7:0] RCV_DATA;
  wire   [1:0] STOP_DATA;

  uart_edge_detector_1 U_0 ( .CLK(CLK), .RST(n1), .SERIAL_IN(SERIAL_IN), 
        .START_BIT(START_BIT) );
  uart_error_1 U_1 ( .RST(n1), .CLK(CLK), .RBUF_FULL(RBUF_FULL), .CHK_ERROR(
        CHK_ERROR), .OE(OE) );
  uart_rcu_1 U_2 ( .CLK(CLK), .RST(n1), .START_BIT(START_BIT), .STOP_RCVING(
        STOP_RCVING), .SB_DETECT(SB_DETECT), .RBUF_LOAD(RBUF_LOAD), 
        .TIMER_TRIG(TIMER_TRIG), .CHK_ERROR(CHK_ERROR), .SET_RBUF_FULL(
        SET_RBUF_FULL), .SBC_EN(SBC_EN), .SBC_CLR(SBC_CLR) );
  uart_rcv_buf_1 U_3 ( .CLK(CLK), .RST(n1), .LOAD_RBUF(RBUF_LOAD), .LOAD_DATA(
        LOAD_DATA), .RCV_DATA(RCV_DATA) );
  uart_rcv_buf_full_1 U_4 ( .CLK(CLK), .RST(n1), .CLR_RBUF(CLR_RBUF), 
        .SET_RBUF_FULL(SET_RBUF_FULL), .RBUF_FULL(RBUF_FULL) );
  uart_sb_check_1 U_5 ( .RST(n1), .CLK(CLK), .SBC_CLR(SBC_CLR), .SBC_EN(SBC_EN), .STOP_DATA(STOP_DATA), .SB_DETECT(SB_DETECT), .SBE(SBE) );
  uart_sr_10bit_1 U_6 ( .CLK(CLK), .RST(n1), .SHIFT_STROBE(SHIFT_STROBE), 
        .SERIAL_IN(SERIAL_IN), .LOAD_DATA(LOAD_DATA), .STOP_DATA(STOP_DATA) );
  keyreg_1 U_8 ( .CLK(CLK), .RST(n1), .SBE(SBE), .OE(OE), .RBUF_FULL(RBUF_FULL), .RCV_DATA(RCV_DATA), .PLAINKEY(PLAINKEY), .KEY_ERROR(KEY_ERROR), 
        .PROG_ERROR(PROG_ERROR), .CLR_RBUFF(CLR_RBUF), .PARITY_ERROR(
        PARITY_ERROR) );
  uart_timer_1 U_7 ( .CLK(CLK), .RST(n1), .TIMER_TRIG(TIMER_TRIG), 
        .STOP_RCVING(STOP_RCVING), .SHIFT_STROBE(SHIFT_STROBE) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module EDBlock_1 ( BYTE, BYTE_READY, CLK, OPCODE, RST, SERIAL_IN, DATA_IN, 
        KEY_ERROR, PARITY_ERROR, PDATA_READY, PROCESSED_DATA, PROG_ERROR, 
        RBUF_FULL, W_ENABLE, R_ENABLE, DATA, ADDR );
  input [7:0] BYTE;
  input [1:0] OPCODE;
  input [7:0] DATA_IN;
  output [7:0] PROCESSED_DATA;
  output [7:0] DATA;
  output [7:0] ADDR;
  input BYTE_READY, CLK, RST, SERIAL_IN;
  output KEY_ERROR, PARITY_ERROR, PDATA_READY, PROG_ERROR, RBUF_FULL, W_ENABLE,
         R_ENABLE;
  wire   n1, n2;
  wire   [63:0] PLAINKEY;

  KSA_1 U_0 ( .KEY(PLAINKEY), .CLK(CLK), .RST(n1), .KEY_ERROR(KEY_ERROR), 
        .BYTE_READY(BYTE_READY), .BYTE(BYTE), .OPCODE(OPCODE), .DATA_IN(
        DATA_IN), .PROCESSED_DATA(PROCESSED_DATA), .PDATA_READY(PDATA_READY), 
        .W_ENABLE(W_ENABLE), .R_ENABLE(R_ENABLE), .ADDR(ADDR), .DATA(DATA) );
  uart_rcv_block_1 U_1 ( .CLK(CLK), .RST(n1), .SERIAL_IN(SERIAL_IN), 
        .KEY_ERROR(KEY_ERROR), .PROG_ERROR(PROG_ERROR), .PLAINKEY(PLAINKEY), 
        .RBUF_FULL(RBUF_FULL), .PARITY_ERROR(PARITY_ERROR) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module RBUFFER_1 ( CLK, RST, NEXT_BYTE, DATA, OPCODE, BYTE_COUNT, EOP, B_READY, 
        R_ENABLE, PRGA_IN, PRGA_OPCODE );
  input [7:0] DATA;
  input [1:0] OPCODE;
  input [4:0] BYTE_COUNT;
  output [7:0] PRGA_IN;
  output [1:0] PRGA_OPCODE;
  input CLK, RST, NEXT_BYTE, EOP;
  output B_READY, R_ENABLE;
  wire   N39, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n97, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n86, n88, n89, n90, n91;
  wire   [2:0] state;
  wire   [2:0] nextState;
  wire   [7:0] tempData;
  wire   [1:0] tempOpcode;
  assign N39 = BYTE_COUNT[4];

  DFFPOSX1 B_READY_reg ( .D(n97), .CLK(CLK), .Q(B_READY) );
  DFFPOSX1 \tempData_reg[7]  ( .D(n71), .CLK(CLK), .Q(tempData[7]) );
  DFFPOSX1 \tempData_reg[6]  ( .D(n72), .CLK(CLK), .Q(tempData[6]) );
  DFFPOSX1 \tempData_reg[5]  ( .D(n73), .CLK(CLK), .Q(tempData[5]) );
  DFFPOSX1 \tempData_reg[4]  ( .D(n74), .CLK(CLK), .Q(tempData[4]) );
  DFFPOSX1 \tempData_reg[3]  ( .D(n75), .CLK(CLK), .Q(tempData[3]) );
  DFFPOSX1 \tempData_reg[2]  ( .D(n86), .CLK(CLK), .Q(tempData[2]) );
  DFFPOSX1 \tempData_reg[1]  ( .D(n88), .CLK(CLK), .Q(tempData[1]) );
  DFFPOSX1 \tempData_reg[0]  ( .D(n89), .CLK(CLK), .Q(tempData[0]) );
  DFFPOSX1 \tempOpcode_reg[1]  ( .D(n90), .CLK(CLK), .Q(tempOpcode[1]) );
  DFFPOSX1 \PRGA_OPCODE_reg[1]  ( .D(n87), .CLK(CLK), .Q(PRGA_OPCODE[1]) );
  DFFPOSX1 \tempOpcode_reg[0]  ( .D(n91), .CLK(CLK), .Q(tempOpcode[0]) );
  DFFPOSX1 \PRGA_OPCODE_reg[0]  ( .D(n85), .CLK(CLK), .Q(PRGA_OPCODE[0]) );
  DFFPOSX1 R_ENABLE_reg ( .D(n84), .CLK(CLK), .Q(R_ENABLE) );
  DFFPOSX1 \PRGA_IN_reg[7]  ( .D(n83), .CLK(CLK), .Q(PRGA_IN[7]) );
  DFFPOSX1 \PRGA_IN_reg[6]  ( .D(n82), .CLK(CLK), .Q(PRGA_IN[6]) );
  DFFPOSX1 \PRGA_IN_reg[5]  ( .D(n81), .CLK(CLK), .Q(PRGA_IN[5]) );
  DFFPOSX1 \PRGA_IN_reg[4]  ( .D(n80), .CLK(CLK), .Q(PRGA_IN[4]) );
  DFFPOSX1 \PRGA_IN_reg[3]  ( .D(n79), .CLK(CLK), .Q(PRGA_IN[3]) );
  DFFPOSX1 \PRGA_IN_reg[2]  ( .D(n78), .CLK(CLK), .Q(PRGA_IN[2]) );
  DFFPOSX1 \PRGA_IN_reg[1]  ( .D(n77), .CLK(CLK), .Q(PRGA_IN[1]) );
  DFFPOSX1 \PRGA_IN_reg[0]  ( .D(n76), .CLK(CLK), .Q(PRGA_IN[0]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[0]) );
  INVX2 U6 ( .A(n44), .Y(n31) );
  INVX2 U7 ( .A(RST), .Y(n4) );
  OR2X2 U8 ( .A(n42), .B(RST), .Y(n32) );
  AND2X2 U9 ( .A(n42), .B(n4), .Y(n47) );
  OAI21X1 U10 ( .A(n5), .B(n6), .C(n7), .Y(nextState[2]) );
  MUX2X1 U11 ( .B(n8), .A(n9), .S(state[0]), .Y(n7) );
  NOR2X1 U12 ( .A(state[2]), .B(n10), .Y(n9) );
  AND2X1 U13 ( .A(state[2]), .B(n11), .Y(n8) );
  OAI21X1 U14 ( .A(NEXT_BYTE), .B(n12), .C(state[1]), .Y(n11) );
  AND2X1 U15 ( .A(n13), .B(NEXT_BYTE), .Y(n5) );
  OAI21X1 U16 ( .A(state[2]), .B(n14), .C(n15), .Y(nextState[1]) );
  OAI21X1 U17 ( .A(n16), .B(n17), .C(n18), .Y(n15) );
  INVX1 U18 ( .A(n6), .Y(n17) );
  OAI21X1 U19 ( .A(state[2]), .B(n19), .C(n20), .Y(nextState[0]) );
  AOI22X1 U20 ( .A(n21), .B(n22), .C(NEXT_BYTE), .D(n23), .Y(n20) );
  OAI21X1 U21 ( .A(n13), .B(n6), .C(n24), .Y(n23) );
  INVX1 U22 ( .A(n16), .Y(n24) );
  NOR2X1 U23 ( .A(n19), .B(n12), .Y(n16) );
  NOR2X1 U24 ( .A(n25), .B(N39), .Y(n12) );
  NAND3X1 U25 ( .A(state[0]), .B(n10), .C(state[2]), .Y(n6) );
  AND2X1 U26 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n13) );
  OAI21X1 U27 ( .A(n26), .B(n18), .C(n27), .Y(n22) );
  INVX1 U28 ( .A(NEXT_BYTE), .Y(n18) );
  AOI21X1 U29 ( .A(EOP), .B(n25), .C(N39), .Y(n26) );
  NAND2X1 U30 ( .A(n28), .B(n29), .Y(n25) );
  NOR2X1 U31 ( .A(BYTE_COUNT[3]), .B(BYTE_COUNT[2]), .Y(n29) );
  NOR2X1 U32 ( .A(BYTE_COUNT[1]), .B(BYTE_COUNT[0]), .Y(n28) );
  NOR2X1 U33 ( .A(state[1]), .B(state[0]), .Y(n21) );
  INVX1 U34 ( .A(n30), .Y(n71) );
  AOI22X1 U35 ( .A(n31), .B(DATA[7]), .C(n32), .D(tempData[7]), .Y(n30) );
  INVX1 U36 ( .A(n33), .Y(n72) );
  AOI22X1 U37 ( .A(n31), .B(DATA[6]), .C(n32), .D(tempData[6]), .Y(n33) );
  INVX1 U38 ( .A(n34), .Y(n73) );
  AOI22X1 U39 ( .A(n31), .B(DATA[5]), .C(n32), .D(tempData[5]), .Y(n34) );
  INVX1 U40 ( .A(n35), .Y(n74) );
  AOI22X1 U41 ( .A(n31), .B(DATA[4]), .C(n32), .D(tempData[4]), .Y(n35) );
  INVX1 U42 ( .A(n36), .Y(n75) );
  AOI22X1 U43 ( .A(n31), .B(DATA[3]), .C(n32), .D(tempData[3]), .Y(n36) );
  INVX1 U44 ( .A(n37), .Y(n86) );
  AOI22X1 U45 ( .A(n31), .B(DATA[2]), .C(n32), .D(tempData[2]), .Y(n37) );
  INVX1 U46 ( .A(n38), .Y(n88) );
  AOI22X1 U47 ( .A(n31), .B(DATA[1]), .C(n32), .D(tempData[1]), .Y(n38) );
  INVX1 U48 ( .A(n39), .Y(n89) );
  AOI22X1 U49 ( .A(n31), .B(DATA[0]), .C(n32), .D(tempData[0]), .Y(n39) );
  INVX1 U50 ( .A(n40), .Y(n90) );
  AOI22X1 U51 ( .A(OPCODE[1]), .B(n31), .C(n32), .D(tempOpcode[1]), .Y(n40) );
  INVX1 U52 ( .A(n41), .Y(n91) );
  AOI22X1 U53 ( .A(OPCODE[0]), .B(n31), .C(n32), .D(tempOpcode[0]), .Y(n41) );
  OAI21X1 U54 ( .A(n4), .B(n43), .C(n44), .Y(n97) );
  INVX1 U55 ( .A(B_READY), .Y(n43) );
  OAI21X1 U56 ( .A(n4), .B(n45), .C(n46), .Y(n87) );
  AOI22X1 U57 ( .A(n31), .B(OPCODE[1]), .C(n47), .D(tempOpcode[1]), .Y(n46) );
  INVX1 U58 ( .A(PRGA_OPCODE[1]), .Y(n45) );
  OAI21X1 U59 ( .A(n4), .B(n48), .C(n49), .Y(n85) );
  AOI22X1 U60 ( .A(n31), .B(OPCODE[0]), .C(n47), .D(tempOpcode[0]), .Y(n49) );
  INVX1 U61 ( .A(PRGA_OPCODE[0]), .Y(n48) );
  MUX2X1 U62 ( .B(n50), .A(n51), .S(RST), .Y(n84) );
  INVX1 U63 ( .A(R_ENABLE), .Y(n51) );
  NAND3X1 U64 ( .A(n10), .B(n27), .C(state[0]), .Y(n50) );
  OAI21X1 U65 ( .A(n4), .B(n52), .C(n53), .Y(n83) );
  AOI22X1 U66 ( .A(DATA[7]), .B(n31), .C(n47), .D(tempData[7]), .Y(n53) );
  INVX1 U67 ( .A(PRGA_IN[7]), .Y(n52) );
  OAI21X1 U68 ( .A(n4), .B(n54), .C(n55), .Y(n82) );
  AOI22X1 U69 ( .A(DATA[6]), .B(n31), .C(n47), .D(tempData[6]), .Y(n55) );
  INVX1 U70 ( .A(PRGA_IN[6]), .Y(n54) );
  OAI21X1 U71 ( .A(n4), .B(n56), .C(n57), .Y(n81) );
  AOI22X1 U72 ( .A(DATA[5]), .B(n31), .C(n47), .D(tempData[5]), .Y(n57) );
  INVX1 U73 ( .A(PRGA_IN[5]), .Y(n56) );
  OAI21X1 U74 ( .A(n4), .B(n58), .C(n59), .Y(n80) );
  AOI22X1 U75 ( .A(DATA[4]), .B(n31), .C(n47), .D(tempData[4]), .Y(n59) );
  INVX1 U76 ( .A(PRGA_IN[4]), .Y(n58) );
  OAI21X1 U77 ( .A(n4), .B(n60), .C(n61), .Y(n79) );
  AOI22X1 U78 ( .A(DATA[3]), .B(n31), .C(n47), .D(tempData[3]), .Y(n61) );
  INVX1 U79 ( .A(PRGA_IN[3]), .Y(n60) );
  OAI21X1 U80 ( .A(n4), .B(n62), .C(n63), .Y(n78) );
  AOI22X1 U81 ( .A(DATA[2]), .B(n31), .C(n47), .D(tempData[2]), .Y(n63) );
  INVX1 U82 ( .A(PRGA_IN[2]), .Y(n62) );
  OAI21X1 U83 ( .A(n4), .B(n64), .C(n65), .Y(n77) );
  AOI22X1 U84 ( .A(DATA[1]), .B(n31), .C(n47), .D(tempData[1]), .Y(n65) );
  INVX1 U85 ( .A(PRGA_IN[1]), .Y(n64) );
  OAI21X1 U86 ( .A(n4), .B(n66), .C(n67), .Y(n76) );
  AOI22X1 U87 ( .A(DATA[0]), .B(n31), .C(n47), .D(tempData[0]), .Y(n67) );
  NAND2X1 U88 ( .A(n14), .B(state[2]), .Y(n42) );
  INVX1 U89 ( .A(n68), .Y(n14) );
  OAI21X1 U90 ( .A(state[1]), .B(n69), .C(n19), .Y(n68) );
  NAND2X1 U91 ( .A(state[1]), .B(n69), .Y(n19) );
  NAND3X1 U92 ( .A(n69), .B(n10), .C(n70), .Y(n44) );
  NOR2X1 U93 ( .A(RST), .B(n27), .Y(n70) );
  INVX1 U94 ( .A(state[2]), .Y(n27) );
  INVX1 U95 ( .A(state[1]), .Y(n10) );
  INVX1 U96 ( .A(state[0]), .Y(n69) );
  INVX1 U97 ( .A(PRGA_IN[0]), .Y(n66) );
endmodule


module RFIFO_1 ( CLK, RST, W_ENABLE, R_ENABLE, RCV_DATA, RCV_OPCODE, DATA, 
        OUT_OPCODE, BYTE_COUNT, EMPTY, FULL );
  input [7:0] RCV_DATA;
  input [1:0] RCV_OPCODE;
  output [7:0] DATA;
  output [1:0] OUT_OPCODE;
  output [4:0] BYTE_COUNT;
  input CLK, RST, W_ENABLE, R_ENABLE;
  output EMPTY, FULL;
  wire   state, N32, N33, N34, N43, N44, N45, N46, \opcode[0][1] ,
         \opcode[0][0] , \opcode[1][1] , \opcode[1][0] , \opcode[2][1] ,
         \opcode[2][0] , \opcode[3][1] , \opcode[3][0] , \opcode[4][1] ,
         \opcode[4][0] , \opcode[5][1] , \opcode[5][0] , \opcode[6][1] ,
         \opcode[6][0] , \opcode[7][1] , \opcode[7][0] , \opcode[8][1] ,
         \opcode[8][0] , \opcode[9][1] , \opcode[9][0] , \opcode[10][1] ,
         \opcode[10][0] , \opcode[11][1] , \opcode[11][0] , \opcode[12][1] ,
         \opcode[12][0] , \opcode[13][1] , \opcode[13][0] , \opcode[14][1] ,
         \opcode[14][0] , \opcode[15][1] , \opcode[15][0] , \opcode[16][1] ,
         \opcode[16][0] , \opcode[17][1] , \opcode[17][0] , \opcode[18][1] ,
         \opcode[18][0] , \opcode[19][1] , \opcode[19][0] , \opcode[20][1] ,
         \opcode[20][0] , \opcode[21][1] , \opcode[21][0] , \opcode[22][1] ,
         \opcode[22][0] , \opcode[23][1] , \opcode[23][0] , \opcode[24][1] ,
         \opcode[24][0] , \opcode[25][1] , \opcode[25][0] , \opcode[26][1] ,
         \opcode[26][0] , \opcode[27][1] , \opcode[27][0] , \opcode[28][1] ,
         \opcode[28][0] , \opcode[29][1] , \opcode[29][0] , \opcode[30][1] ,
         \opcode[30][0] , \opcode[31][1] , \opcode[31][0] , \memory[0][7] ,
         \memory[0][6] , \memory[0][5] , \memory[0][4] , \memory[0][3] ,
         \memory[0][2] , \memory[0][1] , \memory[0][0] , \memory[1][7] ,
         \memory[1][6] , \memory[1][5] , \memory[1][4] , \memory[1][3] ,
         \memory[1][2] , \memory[1][1] , \memory[1][0] , \memory[2][7] ,
         \memory[2][6] , \memory[2][5] , \memory[2][4] , \memory[2][3] ,
         \memory[2][2] , \memory[2][1] , \memory[2][0] , \memory[3][7] ,
         \memory[3][6] , \memory[3][5] , \memory[3][4] , \memory[3][3] ,
         \memory[3][2] , \memory[3][1] , \memory[3][0] , \memory[4][7] ,
         \memory[4][6] , \memory[4][5] , \memory[4][4] , \memory[4][3] ,
         \memory[4][2] , \memory[4][1] , \memory[4][0] , \memory[5][7] ,
         \memory[5][6] , \memory[5][5] , \memory[5][4] , \memory[5][3] ,
         \memory[5][2] , \memory[5][1] , \memory[5][0] , \memory[6][7] ,
         \memory[6][6] , \memory[6][5] , \memory[6][4] , \memory[6][3] ,
         \memory[6][2] , \memory[6][1] , \memory[6][0] , \memory[7][7] ,
         \memory[7][6] , \memory[7][5] , \memory[7][4] , \memory[7][3] ,
         \memory[7][2] , \memory[7][1] , \memory[7][0] , \memory[8][7] ,
         \memory[8][6] , \memory[8][5] , \memory[8][4] , \memory[8][3] ,
         \memory[8][2] , \memory[8][1] , \memory[8][0] , \memory[9][7] ,
         \memory[9][6] , \memory[9][5] , \memory[9][4] , \memory[9][3] ,
         \memory[9][2] , \memory[9][1] , \memory[9][0] , \memory[10][7] ,
         \memory[10][6] , \memory[10][5] , \memory[10][4] , \memory[10][3] ,
         \memory[10][2] , \memory[10][1] , \memory[10][0] , \memory[11][7] ,
         \memory[11][6] , \memory[11][5] , \memory[11][4] , \memory[11][3] ,
         \memory[11][2] , \memory[11][1] , \memory[11][0] , \memory[12][7] ,
         \memory[12][6] , \memory[12][5] , \memory[12][4] , \memory[12][3] ,
         \memory[12][2] , \memory[12][1] , \memory[12][0] , \memory[13][7] ,
         \memory[13][6] , \memory[13][5] , \memory[13][4] , \memory[13][3] ,
         \memory[13][2] , \memory[13][1] , \memory[13][0] , \memory[14][7] ,
         \memory[14][6] , \memory[14][5] , \memory[14][4] , \memory[14][3] ,
         \memory[14][2] , \memory[14][1] , \memory[14][0] , \memory[15][7] ,
         \memory[15][6] , \memory[15][5] , \memory[15][4] , \memory[15][3] ,
         \memory[15][2] , \memory[15][1] , \memory[15][0] , \memory[16][7] ,
         \memory[16][6] , \memory[16][5] , \memory[16][4] , \memory[16][3] ,
         \memory[16][2] , \memory[16][1] , \memory[16][0] , \memory[17][7] ,
         \memory[17][6] , \memory[17][5] , \memory[17][4] , \memory[17][3] ,
         \memory[17][2] , \memory[17][1] , \memory[17][0] , \memory[18][7] ,
         \memory[18][6] , \memory[18][5] , \memory[18][4] , \memory[18][3] ,
         \memory[18][2] , \memory[18][1] , \memory[18][0] , \memory[19][7] ,
         \memory[19][6] , \memory[19][5] , \memory[19][4] , \memory[19][3] ,
         \memory[19][2] , \memory[19][1] , \memory[19][0] , \memory[20][7] ,
         \memory[20][6] , \memory[20][5] , \memory[20][4] , \memory[20][3] ,
         \memory[20][2] , \memory[20][1] , \memory[20][0] , \memory[21][7] ,
         \memory[21][6] , \memory[21][5] , \memory[21][4] , \memory[21][3] ,
         \memory[21][2] , \memory[21][1] , \memory[21][0] , \memory[22][7] ,
         \memory[22][6] , \memory[22][5] , \memory[22][4] , \memory[22][3] ,
         \memory[22][2] , \memory[22][1] , \memory[22][0] , \memory[23][7] ,
         \memory[23][6] , \memory[23][5] , \memory[23][4] , \memory[23][3] ,
         \memory[23][2] , \memory[23][1] , \memory[23][0] , \memory[24][7] ,
         \memory[24][6] , \memory[24][5] , \memory[24][4] , \memory[24][3] ,
         \memory[24][2] , \memory[24][1] , \memory[24][0] , \memory[25][7] ,
         \memory[25][6] , \memory[25][5] , \memory[25][4] , \memory[25][3] ,
         \memory[25][2] , \memory[25][1] , \memory[25][0] , \memory[26][7] ,
         \memory[26][6] , \memory[26][5] , \memory[26][4] , \memory[26][3] ,
         \memory[26][2] , \memory[26][1] , \memory[26][0] , \memory[27][7] ,
         \memory[27][6] , \memory[27][5] , \memory[27][4] , \memory[27][3] ,
         \memory[27][2] , \memory[27][1] , \memory[27][0] , \memory[28][7] ,
         \memory[28][6] , \memory[28][5] , \memory[28][4] , \memory[28][3] ,
         \memory[28][2] , \memory[28][1] , \memory[28][0] , \memory[29][7] ,
         \memory[29][6] , \memory[29][5] , \memory[29][4] , \memory[29][3] ,
         \memory[29][2] , \memory[29][1] , \memory[29][0] , \memory[30][7] ,
         \memory[30][6] , \memory[30][5] , \memory[30][4] , \memory[30][3] ,
         \memory[30][2] , \memory[30][1] , \memory[30][0] , \memory[31][7] ,
         \memory[31][6] , \memory[31][5] , \memory[31][4] , \memory[31][3] ,
         \memory[31][2] , \memory[31][1] , \memory[31][0] , N48, N49, N50, N51,
         N189, N190, N191, N192, N193, N195, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, n854,
         n856, n858, n860, n862, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         \add_76_aco/carry[4] , \add_76_aco/carry[3] , \add_76_aco/carry[2] ,
         \add_76_aco/carry[1] , \sub_72/carry[4] , \sub_72/carry[3] ,
         \sub_72/carry[2] , \sub_72/carry[1] , \add_67/carry[4] ,
         \add_67/carry[3] , \add_67/carry[2] , \r83/carry[4] , \r83/carry[3] ,
         \r83/carry[2] , n1, n2, n3, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n855, n857, n859, n861,
         n863, n864, n865, n866, n867, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198;
  wire   [4:0] readptr;
  wire   [4:0] writeptr;

  DFFSR state_reg ( .D(1'b1), .CLK(CLK), .R(n85), .S(1'b1), .Q(state) );
  DFFPOSX1 FULL_reg ( .D(n1197), .CLK(CLK), .Q(FULL) );
  DFFPOSX1 \memory_reg[0][7]  ( .D(n1172), .CLK(CLK), .Q(\memory[0][7] ) );
  DFFPOSX1 \memory_reg[0][6]  ( .D(n1171), .CLK(CLK), .Q(\memory[0][6] ) );
  DFFPOSX1 \memory_reg[0][5]  ( .D(n1170), .CLK(CLK), .Q(\memory[0][5] ) );
  DFFPOSX1 \memory_reg[0][4]  ( .D(n1169), .CLK(CLK), .Q(\memory[0][4] ) );
  DFFPOSX1 \memory_reg[0][3]  ( .D(n1168), .CLK(CLK), .Q(\memory[0][3] ) );
  DFFPOSX1 \memory_reg[0][2]  ( .D(n1071), .CLK(CLK), .Q(\memory[0][2] ) );
  DFFPOSX1 \memory_reg[0][1]  ( .D(n1070), .CLK(CLK), .Q(\memory[0][1] ) );
  DFFPOSX1 \memory_reg[0][0]  ( .D(n1069), .CLK(CLK), .Q(\memory[0][0] ) );
  DFFPOSX1 \memory_reg[1][7]  ( .D(n1180), .CLK(CLK), .Q(\memory[1][7] ) );
  DFFPOSX1 \memory_reg[1][6]  ( .D(n1179), .CLK(CLK), .Q(\memory[1][6] ) );
  DFFPOSX1 \memory_reg[1][5]  ( .D(n1178), .CLK(CLK), .Q(\memory[1][5] ) );
  DFFPOSX1 \memory_reg[1][4]  ( .D(n1177), .CLK(CLK), .Q(\memory[1][4] ) );
  DFFPOSX1 \memory_reg[1][3]  ( .D(n1176), .CLK(CLK), .Q(\memory[1][3] ) );
  DFFPOSX1 \memory_reg[1][2]  ( .D(n1175), .CLK(CLK), .Q(\memory[1][2] ) );
  DFFPOSX1 \memory_reg[1][1]  ( .D(n1174), .CLK(CLK), .Q(\memory[1][1] ) );
  DFFPOSX1 \memory_reg[1][0]  ( .D(n1173), .CLK(CLK), .Q(\memory[1][0] ) );
  DFFPOSX1 \memory_reg[2][7]  ( .D(n1188), .CLK(CLK), .Q(\memory[2][7] ) );
  DFFPOSX1 \memory_reg[2][6]  ( .D(n1187), .CLK(CLK), .Q(\memory[2][6] ) );
  DFFPOSX1 \memory_reg[2][5]  ( .D(n1186), .CLK(CLK), .Q(\memory[2][5] ) );
  DFFPOSX1 \memory_reg[2][4]  ( .D(n1185), .CLK(CLK), .Q(\memory[2][4] ) );
  DFFPOSX1 \memory_reg[2][3]  ( .D(n1184), .CLK(CLK), .Q(\memory[2][3] ) );
  DFFPOSX1 \memory_reg[2][2]  ( .D(n1183), .CLK(CLK), .Q(\memory[2][2] ) );
  DFFPOSX1 \memory_reg[2][1]  ( .D(n1182), .CLK(CLK), .Q(\memory[2][1] ) );
  DFFPOSX1 \memory_reg[2][0]  ( .D(n1181), .CLK(CLK), .Q(\memory[2][0] ) );
  DFFPOSX1 \memory_reg[3][7]  ( .D(n1196), .CLK(CLK), .Q(\memory[3][7] ) );
  DFFPOSX1 \memory_reg[3][6]  ( .D(n1195), .CLK(CLK), .Q(\memory[3][6] ) );
  DFFPOSX1 \memory_reg[3][5]  ( .D(n1194), .CLK(CLK), .Q(\memory[3][5] ) );
  DFFPOSX1 \memory_reg[3][4]  ( .D(n1193), .CLK(CLK), .Q(\memory[3][4] ) );
  DFFPOSX1 \memory_reg[3][3]  ( .D(n1192), .CLK(CLK), .Q(\memory[3][3] ) );
  DFFPOSX1 \memory_reg[3][2]  ( .D(n1191), .CLK(CLK), .Q(\memory[3][2] ) );
  DFFPOSX1 \memory_reg[3][1]  ( .D(n1190), .CLK(CLK), .Q(\memory[3][1] ) );
  DFFPOSX1 \memory_reg[3][0]  ( .D(n1189), .CLK(CLK), .Q(\memory[3][0] ) );
  DFFPOSX1 \memory_reg[4][7]  ( .D(n869), .CLK(CLK), .Q(\memory[4][7] ) );
  DFFPOSX1 \memory_reg[4][6]  ( .D(n870), .CLK(CLK), .Q(\memory[4][6] ) );
  DFFPOSX1 \memory_reg[4][5]  ( .D(n871), .CLK(CLK), .Q(\memory[4][5] ) );
  DFFPOSX1 \memory_reg[4][4]  ( .D(n872), .CLK(CLK), .Q(\memory[4][4] ) );
  DFFPOSX1 \memory_reg[4][3]  ( .D(n873), .CLK(CLK), .Q(\memory[4][3] ) );
  DFFPOSX1 \memory_reg[4][2]  ( .D(n874), .CLK(CLK), .Q(\memory[4][2] ) );
  DFFPOSX1 \memory_reg[4][1]  ( .D(n875), .CLK(CLK), .Q(\memory[4][1] ) );
  DFFPOSX1 \memory_reg[4][0]  ( .D(n876), .CLK(CLK), .Q(\memory[4][0] ) );
  DFFPOSX1 \memory_reg[5][7]  ( .D(n879), .CLK(CLK), .Q(\memory[5][7] ) );
  DFFPOSX1 \memory_reg[5][6]  ( .D(n880), .CLK(CLK), .Q(\memory[5][6] ) );
  DFFPOSX1 \memory_reg[5][5]  ( .D(n881), .CLK(CLK), .Q(\memory[5][5] ) );
  DFFPOSX1 \memory_reg[5][4]  ( .D(n882), .CLK(CLK), .Q(\memory[5][4] ) );
  DFFPOSX1 \memory_reg[5][3]  ( .D(n883), .CLK(CLK), .Q(\memory[5][3] ) );
  DFFPOSX1 \memory_reg[5][2]  ( .D(n884), .CLK(CLK), .Q(\memory[5][2] ) );
  DFFPOSX1 \memory_reg[5][1]  ( .D(n885), .CLK(CLK), .Q(\memory[5][1] ) );
  DFFPOSX1 \memory_reg[5][0]  ( .D(n886), .CLK(CLK), .Q(\memory[5][0] ) );
  DFFPOSX1 \memory_reg[6][7]  ( .D(n889), .CLK(CLK), .Q(\memory[6][7] ) );
  DFFPOSX1 \memory_reg[6][6]  ( .D(n890), .CLK(CLK), .Q(\memory[6][6] ) );
  DFFPOSX1 \memory_reg[6][5]  ( .D(n891), .CLK(CLK), .Q(\memory[6][5] ) );
  DFFPOSX1 \memory_reg[6][4]  ( .D(n892), .CLK(CLK), .Q(\memory[6][4] ) );
  DFFPOSX1 \memory_reg[6][3]  ( .D(n893), .CLK(CLK), .Q(\memory[6][3] ) );
  DFFPOSX1 \memory_reg[6][2]  ( .D(n894), .CLK(CLK), .Q(\memory[6][2] ) );
  DFFPOSX1 \memory_reg[6][1]  ( .D(n895), .CLK(CLK), .Q(\memory[6][1] ) );
  DFFPOSX1 \memory_reg[6][0]  ( .D(n896), .CLK(CLK), .Q(\memory[6][0] ) );
  DFFPOSX1 \memory_reg[7][7]  ( .D(n899), .CLK(CLK), .Q(\memory[7][7] ) );
  DFFPOSX1 \memory_reg[7][6]  ( .D(n900), .CLK(CLK), .Q(\memory[7][6] ) );
  DFFPOSX1 \memory_reg[7][5]  ( .D(n901), .CLK(CLK), .Q(\memory[7][5] ) );
  DFFPOSX1 \memory_reg[7][4]  ( .D(n902), .CLK(CLK), .Q(\memory[7][4] ) );
  DFFPOSX1 \memory_reg[7][3]  ( .D(n903), .CLK(CLK), .Q(\memory[7][3] ) );
  DFFPOSX1 \memory_reg[7][2]  ( .D(n904), .CLK(CLK), .Q(\memory[7][2] ) );
  DFFPOSX1 \memory_reg[7][1]  ( .D(n905), .CLK(CLK), .Q(\memory[7][1] ) );
  DFFPOSX1 \memory_reg[7][0]  ( .D(n906), .CLK(CLK), .Q(\memory[7][0] ) );
  DFFPOSX1 \memory_reg[8][7]  ( .D(n1167), .CLK(CLK), .Q(\memory[8][7] ) );
  DFFPOSX1 \memory_reg[8][6]  ( .D(n1166), .CLK(CLK), .Q(\memory[8][6] ) );
  DFFPOSX1 \memory_reg[8][5]  ( .D(n1165), .CLK(CLK), .Q(\memory[8][5] ) );
  DFFPOSX1 \memory_reg[8][4]  ( .D(n1164), .CLK(CLK), .Q(\memory[8][4] ) );
  DFFPOSX1 \memory_reg[8][3]  ( .D(n1163), .CLK(CLK), .Q(\memory[8][3] ) );
  DFFPOSX1 \memory_reg[8][2]  ( .D(n1162), .CLK(CLK), .Q(\memory[8][2] ) );
  DFFPOSX1 \memory_reg[8][1]  ( .D(n1161), .CLK(CLK), .Q(\memory[8][1] ) );
  DFFPOSX1 \memory_reg[8][0]  ( .D(n1160), .CLK(CLK), .Q(\memory[8][0] ) );
  DFFPOSX1 \memory_reg[9][7]  ( .D(n1159), .CLK(CLK), .Q(\memory[9][7] ) );
  DFFPOSX1 \memory_reg[9][6]  ( .D(n1158), .CLK(CLK), .Q(\memory[9][6] ) );
  DFFPOSX1 \memory_reg[9][5]  ( .D(n1157), .CLK(CLK), .Q(\memory[9][5] ) );
  DFFPOSX1 \memory_reg[9][4]  ( .D(n1156), .CLK(CLK), .Q(\memory[9][4] ) );
  DFFPOSX1 \memory_reg[9][3]  ( .D(n1155), .CLK(CLK), .Q(\memory[9][3] ) );
  DFFPOSX1 \memory_reg[9][2]  ( .D(n1154), .CLK(CLK), .Q(\memory[9][2] ) );
  DFFPOSX1 \memory_reg[9][1]  ( .D(n1153), .CLK(CLK), .Q(\memory[9][1] ) );
  DFFPOSX1 \memory_reg[9][0]  ( .D(n1152), .CLK(CLK), .Q(\memory[9][0] ) );
  DFFPOSX1 \memory_reg[10][7]  ( .D(n1151), .CLK(CLK), .Q(\memory[10][7] ) );
  DFFPOSX1 \memory_reg[10][6]  ( .D(n1150), .CLK(CLK), .Q(\memory[10][6] ) );
  DFFPOSX1 \memory_reg[10][5]  ( .D(n1149), .CLK(CLK), .Q(\memory[10][5] ) );
  DFFPOSX1 \memory_reg[10][4]  ( .D(n1148), .CLK(CLK), .Q(\memory[10][4] ) );
  DFFPOSX1 \memory_reg[10][3]  ( .D(n1147), .CLK(CLK), .Q(\memory[10][3] ) );
  DFFPOSX1 \memory_reg[10][2]  ( .D(n1146), .CLK(CLK), .Q(\memory[10][2] ) );
  DFFPOSX1 \memory_reg[10][1]  ( .D(n1145), .CLK(CLK), .Q(\memory[10][1] ) );
  DFFPOSX1 \memory_reg[10][0]  ( .D(n1144), .CLK(CLK), .Q(\memory[10][0] ) );
  DFFPOSX1 \memory_reg[11][7]  ( .D(n1143), .CLK(CLK), .Q(\memory[11][7] ) );
  DFFPOSX1 \memory_reg[11][6]  ( .D(n1142), .CLK(CLK), .Q(\memory[11][6] ) );
  DFFPOSX1 \memory_reg[11][5]  ( .D(n1141), .CLK(CLK), .Q(\memory[11][5] ) );
  DFFPOSX1 \memory_reg[11][4]  ( .D(n1140), .CLK(CLK), .Q(\memory[11][4] ) );
  DFFPOSX1 \memory_reg[11][3]  ( .D(n1139), .CLK(CLK), .Q(\memory[11][3] ) );
  DFFPOSX1 \memory_reg[11][2]  ( .D(n1138), .CLK(CLK), .Q(\memory[11][2] ) );
  DFFPOSX1 \memory_reg[11][1]  ( .D(n1137), .CLK(CLK), .Q(\memory[11][1] ) );
  DFFPOSX1 \memory_reg[11][0]  ( .D(n1136), .CLK(CLK), .Q(\memory[11][0] ) );
  DFFPOSX1 \memory_reg[12][7]  ( .D(n1027), .CLK(CLK), .Q(\memory[12][7] ) );
  DFFPOSX1 \memory_reg[12][6]  ( .D(n1028), .CLK(CLK), .Q(\memory[12][6] ) );
  DFFPOSX1 \memory_reg[12][5]  ( .D(n1029), .CLK(CLK), .Q(\memory[12][5] ) );
  DFFPOSX1 \memory_reg[12][4]  ( .D(n1064), .CLK(CLK), .Q(\memory[12][4] ) );
  DFFPOSX1 \memory_reg[12][3]  ( .D(n1065), .CLK(CLK), .Q(\memory[12][3] ) );
  DFFPOSX1 \memory_reg[12][2]  ( .D(n1066), .CLK(CLK), .Q(\memory[12][2] ) );
  DFFPOSX1 \memory_reg[12][1]  ( .D(n1067), .CLK(CLK), .Q(\memory[12][1] ) );
  DFFPOSX1 \memory_reg[12][0]  ( .D(n1068), .CLK(CLK), .Q(\memory[12][0] ) );
  DFFPOSX1 \memory_reg[13][7]  ( .D(n1019), .CLK(CLK), .Q(\memory[13][7] ) );
  DFFPOSX1 \memory_reg[13][6]  ( .D(n1020), .CLK(CLK), .Q(\memory[13][6] ) );
  DFFPOSX1 \memory_reg[13][5]  ( .D(n1021), .CLK(CLK), .Q(\memory[13][5] ) );
  DFFPOSX1 \memory_reg[13][4]  ( .D(n1022), .CLK(CLK), .Q(\memory[13][4] ) );
  DFFPOSX1 \memory_reg[13][3]  ( .D(n1023), .CLK(CLK), .Q(\memory[13][3] ) );
  DFFPOSX1 \memory_reg[13][2]  ( .D(n1024), .CLK(CLK), .Q(\memory[13][2] ) );
  DFFPOSX1 \memory_reg[13][1]  ( .D(n1025), .CLK(CLK), .Q(\memory[13][1] ) );
  DFFPOSX1 \memory_reg[13][0]  ( .D(n1026), .CLK(CLK), .Q(\memory[13][0] ) );
  DFFPOSX1 \memory_reg[14][7]  ( .D(n1011), .CLK(CLK), .Q(\memory[14][7] ) );
  DFFPOSX1 \memory_reg[14][6]  ( .D(n1012), .CLK(CLK), .Q(\memory[14][6] ) );
  DFFPOSX1 \memory_reg[14][5]  ( .D(n1013), .CLK(CLK), .Q(\memory[14][5] ) );
  DFFPOSX1 \memory_reg[14][4]  ( .D(n1014), .CLK(CLK), .Q(\memory[14][4] ) );
  DFFPOSX1 \memory_reg[14][3]  ( .D(n1015), .CLK(CLK), .Q(\memory[14][3] ) );
  DFFPOSX1 \memory_reg[14][2]  ( .D(n1016), .CLK(CLK), .Q(\memory[14][2] ) );
  DFFPOSX1 \memory_reg[14][1]  ( .D(n1017), .CLK(CLK), .Q(\memory[14][1] ) );
  DFFPOSX1 \memory_reg[14][0]  ( .D(n1018), .CLK(CLK), .Q(\memory[14][0] ) );
  DFFPOSX1 \memory_reg[15][7]  ( .D(n1003), .CLK(CLK), .Q(\memory[15][7] ) );
  DFFPOSX1 \memory_reg[15][6]  ( .D(n1004), .CLK(CLK), .Q(\memory[15][6] ) );
  DFFPOSX1 \memory_reg[15][5]  ( .D(n1005), .CLK(CLK), .Q(\memory[15][5] ) );
  DFFPOSX1 \memory_reg[15][4]  ( .D(n1006), .CLK(CLK), .Q(\memory[15][4] ) );
  DFFPOSX1 \memory_reg[15][3]  ( .D(n1007), .CLK(CLK), .Q(\memory[15][3] ) );
  DFFPOSX1 \memory_reg[15][2]  ( .D(n1008), .CLK(CLK), .Q(\memory[15][2] ) );
  DFFPOSX1 \memory_reg[15][1]  ( .D(n1009), .CLK(CLK), .Q(\memory[15][1] ) );
  DFFPOSX1 \memory_reg[15][0]  ( .D(n1010), .CLK(CLK), .Q(\memory[15][0] ) );
  DFFPOSX1 \memory_reg[16][7]  ( .D(n1135), .CLK(CLK), .Q(\memory[16][7] ) );
  DFFPOSX1 \memory_reg[16][6]  ( .D(n1134), .CLK(CLK), .Q(\memory[16][6] ) );
  DFFPOSX1 \memory_reg[16][5]  ( .D(n1133), .CLK(CLK), .Q(\memory[16][5] ) );
  DFFPOSX1 \memory_reg[16][4]  ( .D(n1132), .CLK(CLK), .Q(\memory[16][4] ) );
  DFFPOSX1 \memory_reg[16][3]  ( .D(n1131), .CLK(CLK), .Q(\memory[16][3] ) );
  DFFPOSX1 \memory_reg[16][2]  ( .D(n1130), .CLK(CLK), .Q(\memory[16][2] ) );
  DFFPOSX1 \memory_reg[16][1]  ( .D(n1129), .CLK(CLK), .Q(\memory[16][1] ) );
  DFFPOSX1 \memory_reg[16][0]  ( .D(n1128), .CLK(CLK), .Q(\memory[16][0] ) );
  DFFPOSX1 \memory_reg[17][7]  ( .D(n1127), .CLK(CLK), .Q(\memory[17][7] ) );
  DFFPOSX1 \memory_reg[17][6]  ( .D(n1126), .CLK(CLK), .Q(\memory[17][6] ) );
  DFFPOSX1 \memory_reg[17][5]  ( .D(n1125), .CLK(CLK), .Q(\memory[17][5] ) );
  DFFPOSX1 \memory_reg[17][4]  ( .D(n1124), .CLK(CLK), .Q(\memory[17][4] ) );
  DFFPOSX1 \memory_reg[17][3]  ( .D(n1123), .CLK(CLK), .Q(\memory[17][3] ) );
  DFFPOSX1 \memory_reg[17][2]  ( .D(n1122), .CLK(CLK), .Q(\memory[17][2] ) );
  DFFPOSX1 \memory_reg[17][1]  ( .D(n1121), .CLK(CLK), .Q(\memory[17][1] ) );
  DFFPOSX1 \memory_reg[17][0]  ( .D(n1120), .CLK(CLK), .Q(\memory[17][0] ) );
  DFFPOSX1 \memory_reg[18][7]  ( .D(n1119), .CLK(CLK), .Q(\memory[18][7] ) );
  DFFPOSX1 \memory_reg[18][6]  ( .D(n1118), .CLK(CLK), .Q(\memory[18][6] ) );
  DFFPOSX1 \memory_reg[18][5]  ( .D(n1117), .CLK(CLK), .Q(\memory[18][5] ) );
  DFFPOSX1 \memory_reg[18][4]  ( .D(n1116), .CLK(CLK), .Q(\memory[18][4] ) );
  DFFPOSX1 \memory_reg[18][3]  ( .D(n1115), .CLK(CLK), .Q(\memory[18][3] ) );
  DFFPOSX1 \memory_reg[18][2]  ( .D(n1114), .CLK(CLK), .Q(\memory[18][2] ) );
  DFFPOSX1 \memory_reg[18][1]  ( .D(n1113), .CLK(CLK), .Q(\memory[18][1] ) );
  DFFPOSX1 \memory_reg[18][0]  ( .D(n1112), .CLK(CLK), .Q(\memory[18][0] ) );
  DFFPOSX1 \memory_reg[19][7]  ( .D(n1111), .CLK(CLK), .Q(\memory[19][7] ) );
  DFFPOSX1 \memory_reg[19][6]  ( .D(n1110), .CLK(CLK), .Q(\memory[19][6] ) );
  DFFPOSX1 \memory_reg[19][5]  ( .D(n1109), .CLK(CLK), .Q(\memory[19][5] ) );
  DFFPOSX1 \memory_reg[19][4]  ( .D(n1108), .CLK(CLK), .Q(\memory[19][4] ) );
  DFFPOSX1 \memory_reg[19][3]  ( .D(n1107), .CLK(CLK), .Q(\memory[19][3] ) );
  DFFPOSX1 \memory_reg[19][2]  ( .D(n1106), .CLK(CLK), .Q(\memory[19][2] ) );
  DFFPOSX1 \memory_reg[19][1]  ( .D(n1105), .CLK(CLK), .Q(\memory[19][1] ) );
  DFFPOSX1 \memory_reg[19][0]  ( .D(n1104), .CLK(CLK), .Q(\memory[19][0] ) );
  DFFPOSX1 \memory_reg[20][7]  ( .D(n995), .CLK(CLK), .Q(\memory[20][7] ) );
  DFFPOSX1 \memory_reg[20][6]  ( .D(n996), .CLK(CLK), .Q(\memory[20][6] ) );
  DFFPOSX1 \memory_reg[20][5]  ( .D(n997), .CLK(CLK), .Q(\memory[20][5] ) );
  DFFPOSX1 \memory_reg[20][4]  ( .D(n998), .CLK(CLK), .Q(\memory[20][4] ) );
  DFFPOSX1 \memory_reg[20][3]  ( .D(n999), .CLK(CLK), .Q(\memory[20][3] ) );
  DFFPOSX1 \memory_reg[20][2]  ( .D(n1000), .CLK(CLK), .Q(\memory[20][2] ) );
  DFFPOSX1 \memory_reg[20][1]  ( .D(n1001), .CLK(CLK), .Q(\memory[20][1] ) );
  DFFPOSX1 \memory_reg[20][0]  ( .D(n1002), .CLK(CLK), .Q(\memory[20][0] ) );
  DFFPOSX1 \memory_reg[21][7]  ( .D(n987), .CLK(CLK), .Q(\memory[21][7] ) );
  DFFPOSX1 \memory_reg[21][6]  ( .D(n988), .CLK(CLK), .Q(\memory[21][6] ) );
  DFFPOSX1 \memory_reg[21][5]  ( .D(n989), .CLK(CLK), .Q(\memory[21][5] ) );
  DFFPOSX1 \memory_reg[21][4]  ( .D(n990), .CLK(CLK), .Q(\memory[21][4] ) );
  DFFPOSX1 \memory_reg[21][3]  ( .D(n991), .CLK(CLK), .Q(\memory[21][3] ) );
  DFFPOSX1 \memory_reg[21][2]  ( .D(n992), .CLK(CLK), .Q(\memory[21][2] ) );
  DFFPOSX1 \memory_reg[21][1]  ( .D(n993), .CLK(CLK), .Q(\memory[21][1] ) );
  DFFPOSX1 \memory_reg[21][0]  ( .D(n994), .CLK(CLK), .Q(\memory[21][0] ) );
  DFFPOSX1 \memory_reg[22][7]  ( .D(n979), .CLK(CLK), .Q(\memory[22][7] ) );
  DFFPOSX1 \memory_reg[22][6]  ( .D(n980), .CLK(CLK), .Q(\memory[22][6] ) );
  DFFPOSX1 \memory_reg[22][5]  ( .D(n981), .CLK(CLK), .Q(\memory[22][5] ) );
  DFFPOSX1 \memory_reg[22][4]  ( .D(n982), .CLK(CLK), .Q(\memory[22][4] ) );
  DFFPOSX1 \memory_reg[22][3]  ( .D(n983), .CLK(CLK), .Q(\memory[22][3] ) );
  DFFPOSX1 \memory_reg[22][2]  ( .D(n984), .CLK(CLK), .Q(\memory[22][2] ) );
  DFFPOSX1 \memory_reg[22][1]  ( .D(n985), .CLK(CLK), .Q(\memory[22][1] ) );
  DFFPOSX1 \memory_reg[22][0]  ( .D(n986), .CLK(CLK), .Q(\memory[22][0] ) );
  DFFPOSX1 \memory_reg[23][7]  ( .D(n971), .CLK(CLK), .Q(\memory[23][7] ) );
  DFFPOSX1 \memory_reg[23][6]  ( .D(n972), .CLK(CLK), .Q(\memory[23][6] ) );
  DFFPOSX1 \memory_reg[23][5]  ( .D(n973), .CLK(CLK), .Q(\memory[23][5] ) );
  DFFPOSX1 \memory_reg[23][4]  ( .D(n974), .CLK(CLK), .Q(\memory[23][4] ) );
  DFFPOSX1 \memory_reg[23][3]  ( .D(n975), .CLK(CLK), .Q(\memory[23][3] ) );
  DFFPOSX1 \memory_reg[23][2]  ( .D(n976), .CLK(CLK), .Q(\memory[23][2] ) );
  DFFPOSX1 \memory_reg[23][1]  ( .D(n977), .CLK(CLK), .Q(\memory[23][1] ) );
  DFFPOSX1 \memory_reg[23][0]  ( .D(n978), .CLK(CLK), .Q(\memory[23][0] ) );
  DFFPOSX1 \memory_reg[24][7]  ( .D(n963), .CLK(CLK), .Q(\memory[24][7] ) );
  DFFPOSX1 \memory_reg[24][6]  ( .D(n964), .CLK(CLK), .Q(\memory[24][6] ) );
  DFFPOSX1 \memory_reg[24][5]  ( .D(n965), .CLK(CLK), .Q(\memory[24][5] ) );
  DFFPOSX1 \memory_reg[24][4]  ( .D(n966), .CLK(CLK), .Q(\memory[24][4] ) );
  DFFPOSX1 \memory_reg[24][3]  ( .D(n967), .CLK(CLK), .Q(\memory[24][3] ) );
  DFFPOSX1 \memory_reg[24][2]  ( .D(n968), .CLK(CLK), .Q(\memory[24][2] ) );
  DFFPOSX1 \memory_reg[24][1]  ( .D(n969), .CLK(CLK), .Q(\memory[24][1] ) );
  DFFPOSX1 \memory_reg[24][0]  ( .D(n970), .CLK(CLK), .Q(\memory[24][0] ) );
  DFFPOSX1 \memory_reg[25][7]  ( .D(n955), .CLK(CLK), .Q(\memory[25][7] ) );
  DFFPOSX1 \memory_reg[25][6]  ( .D(n956), .CLK(CLK), .Q(\memory[25][6] ) );
  DFFPOSX1 \memory_reg[25][5]  ( .D(n957), .CLK(CLK), .Q(\memory[25][5] ) );
  DFFPOSX1 \memory_reg[25][4]  ( .D(n958), .CLK(CLK), .Q(\memory[25][4] ) );
  DFFPOSX1 \memory_reg[25][3]  ( .D(n959), .CLK(CLK), .Q(\memory[25][3] ) );
  DFFPOSX1 \memory_reg[25][2]  ( .D(n960), .CLK(CLK), .Q(\memory[25][2] ) );
  DFFPOSX1 \memory_reg[25][1]  ( .D(n961), .CLK(CLK), .Q(\memory[25][1] ) );
  DFFPOSX1 \memory_reg[25][0]  ( .D(n962), .CLK(CLK), .Q(\memory[25][0] ) );
  DFFPOSX1 \memory_reg[26][7]  ( .D(n947), .CLK(CLK), .Q(\memory[26][7] ) );
  DFFPOSX1 \memory_reg[26][6]  ( .D(n948), .CLK(CLK), .Q(\memory[26][6] ) );
  DFFPOSX1 \memory_reg[26][5]  ( .D(n949), .CLK(CLK), .Q(\memory[26][5] ) );
  DFFPOSX1 \memory_reg[26][4]  ( .D(n950), .CLK(CLK), .Q(\memory[26][4] ) );
  DFFPOSX1 \memory_reg[26][3]  ( .D(n951), .CLK(CLK), .Q(\memory[26][3] ) );
  DFFPOSX1 \memory_reg[26][2]  ( .D(n952), .CLK(CLK), .Q(\memory[26][2] ) );
  DFFPOSX1 \memory_reg[26][1]  ( .D(n953), .CLK(CLK), .Q(\memory[26][1] ) );
  DFFPOSX1 \memory_reg[26][0]  ( .D(n954), .CLK(CLK), .Q(\memory[26][0] ) );
  DFFPOSX1 \memory_reg[27][7]  ( .D(n939), .CLK(CLK), .Q(\memory[27][7] ) );
  DFFPOSX1 \memory_reg[27][6]  ( .D(n940), .CLK(CLK), .Q(\memory[27][6] ) );
  DFFPOSX1 \memory_reg[27][5]  ( .D(n941), .CLK(CLK), .Q(\memory[27][5] ) );
  DFFPOSX1 \memory_reg[27][4]  ( .D(n942), .CLK(CLK), .Q(\memory[27][4] ) );
  DFFPOSX1 \memory_reg[27][3]  ( .D(n943), .CLK(CLK), .Q(\memory[27][3] ) );
  DFFPOSX1 \memory_reg[27][2]  ( .D(n944), .CLK(CLK), .Q(\memory[27][2] ) );
  DFFPOSX1 \memory_reg[27][1]  ( .D(n945), .CLK(CLK), .Q(\memory[27][1] ) );
  DFFPOSX1 \memory_reg[27][0]  ( .D(n946), .CLK(CLK), .Q(\memory[27][0] ) );
  DFFPOSX1 \memory_reg[28][7]  ( .D(n1103), .CLK(CLK), .Q(\memory[28][7] ) );
  DFFPOSX1 \memory_reg[28][6]  ( .D(n1102), .CLK(CLK), .Q(\memory[28][6] ) );
  DFFPOSX1 \memory_reg[28][5]  ( .D(n1101), .CLK(CLK), .Q(\memory[28][5] ) );
  DFFPOSX1 \memory_reg[28][4]  ( .D(n1100), .CLK(CLK), .Q(\memory[28][4] ) );
  DFFPOSX1 \memory_reg[28][3]  ( .D(n1099), .CLK(CLK), .Q(\memory[28][3] ) );
  DFFPOSX1 \memory_reg[28][2]  ( .D(n1098), .CLK(CLK), .Q(\memory[28][2] ) );
  DFFPOSX1 \memory_reg[28][1]  ( .D(n1097), .CLK(CLK), .Q(\memory[28][1] ) );
  DFFPOSX1 \memory_reg[28][0]  ( .D(n1096), .CLK(CLK), .Q(\memory[28][0] ) );
  DFFPOSX1 \memory_reg[29][7]  ( .D(n1095), .CLK(CLK), .Q(\memory[29][7] ) );
  DFFPOSX1 \memory_reg[29][6]  ( .D(n1094), .CLK(CLK), .Q(\memory[29][6] ) );
  DFFPOSX1 \memory_reg[29][5]  ( .D(n1093), .CLK(CLK), .Q(\memory[29][5] ) );
  DFFPOSX1 \memory_reg[29][4]  ( .D(n1092), .CLK(CLK), .Q(\memory[29][4] ) );
  DFFPOSX1 \memory_reg[29][3]  ( .D(n1091), .CLK(CLK), .Q(\memory[29][3] ) );
  DFFPOSX1 \memory_reg[29][2]  ( .D(n1090), .CLK(CLK), .Q(\memory[29][2] ) );
  DFFPOSX1 \memory_reg[29][1]  ( .D(n1089), .CLK(CLK), .Q(\memory[29][1] ) );
  DFFPOSX1 \memory_reg[29][0]  ( .D(n1088), .CLK(CLK), .Q(\memory[29][0] ) );
  DFFPOSX1 \memory_reg[30][7]  ( .D(n1087), .CLK(CLK), .Q(\memory[30][7] ) );
  DFFPOSX1 \memory_reg[30][6]  ( .D(n1086), .CLK(CLK), .Q(\memory[30][6] ) );
  DFFPOSX1 \memory_reg[30][5]  ( .D(n1085), .CLK(CLK), .Q(\memory[30][5] ) );
  DFFPOSX1 \memory_reg[30][4]  ( .D(n1084), .CLK(CLK), .Q(\memory[30][4] ) );
  DFFPOSX1 \memory_reg[30][3]  ( .D(n1083), .CLK(CLK), .Q(\memory[30][3] ) );
  DFFPOSX1 \memory_reg[30][2]  ( .D(n1082), .CLK(CLK), .Q(\memory[30][2] ) );
  DFFPOSX1 \memory_reg[30][1]  ( .D(n1081), .CLK(CLK), .Q(\memory[30][1] ) );
  DFFPOSX1 \memory_reg[30][0]  ( .D(n1080), .CLK(CLK), .Q(\memory[30][0] ) );
  DFFPOSX1 \memory_reg[31][7]  ( .D(n1079), .CLK(CLK), .Q(\memory[31][7] ) );
  DFFPOSX1 \memory_reg[31][6]  ( .D(n1078), .CLK(CLK), .Q(\memory[31][6] ) );
  DFFPOSX1 \memory_reg[31][5]  ( .D(n1077), .CLK(CLK), .Q(\memory[31][5] ) );
  DFFPOSX1 \memory_reg[31][4]  ( .D(n1076), .CLK(CLK), .Q(\memory[31][4] ) );
  DFFPOSX1 \memory_reg[31][3]  ( .D(n1075), .CLK(CLK), .Q(\memory[31][3] ) );
  DFFPOSX1 \memory_reg[31][2]  ( .D(n1074), .CLK(CLK), .Q(\memory[31][2] ) );
  DFFPOSX1 \memory_reg[31][1]  ( .D(n1073), .CLK(CLK), .Q(\memory[31][1] ) );
  DFFPOSX1 \memory_reg[31][0]  ( .D(n1072), .CLK(CLK), .Q(\memory[31][0] ) );
  DFFPOSX1 \opcode_reg[0][1]  ( .D(n932), .CLK(CLK), .Q(\opcode[0][1] ) );
  DFFPOSX1 \opcode_reg[0][0]  ( .D(n931), .CLK(CLK), .Q(\opcode[0][0] ) );
  DFFPOSX1 \opcode_reg[1][1]  ( .D(n934), .CLK(CLK), .Q(\opcode[1][1] ) );
  DFFPOSX1 \opcode_reg[1][0]  ( .D(n933), .CLK(CLK), .Q(\opcode[1][0] ) );
  DFFPOSX1 \opcode_reg[2][1]  ( .D(n936), .CLK(CLK), .Q(\opcode[2][1] ) );
  DFFPOSX1 \opcode_reg[2][0]  ( .D(n935), .CLK(CLK), .Q(\opcode[2][0] ) );
  DFFPOSX1 \opcode_reg[3][1]  ( .D(n938), .CLK(CLK), .Q(\opcode[3][1] ) );
  DFFPOSX1 \opcode_reg[3][0]  ( .D(n937), .CLK(CLK), .Q(\opcode[3][0] ) );
  DFFPOSX1 \opcode_reg[4][1]  ( .D(n877), .CLK(CLK), .Q(\opcode[4][1] ) );
  DFFPOSX1 \opcode_reg[4][0]  ( .D(n878), .CLK(CLK), .Q(\opcode[4][0] ) );
  DFFPOSX1 \opcode_reg[5][1]  ( .D(n887), .CLK(CLK), .Q(\opcode[5][1] ) );
  DFFPOSX1 \opcode_reg[5][0]  ( .D(n888), .CLK(CLK), .Q(\opcode[5][0] ) );
  DFFPOSX1 \opcode_reg[6][1]  ( .D(n897), .CLK(CLK), .Q(\opcode[6][1] ) );
  DFFPOSX1 \opcode_reg[6][0]  ( .D(n898), .CLK(CLK), .Q(\opcode[6][0] ) );
  DFFPOSX1 \opcode_reg[7][1]  ( .D(n907), .CLK(CLK), .Q(\opcode[7][1] ) );
  DFFPOSX1 \opcode_reg[7][0]  ( .D(n908), .CLK(CLK), .Q(\opcode[7][0] ) );
  DFFPOSX1 \opcode_reg[8][1]  ( .D(n1063), .CLK(CLK), .Q(\opcode[8][1] ) );
  DFFPOSX1 \opcode_reg[8][0]  ( .D(n1062), .CLK(CLK), .Q(\opcode[8][0] ) );
  DFFPOSX1 \opcode_reg[9][1]  ( .D(n1061), .CLK(CLK), .Q(\opcode[9][1] ) );
  DFFPOSX1 \opcode_reg[9][0]  ( .D(n1060), .CLK(CLK), .Q(\opcode[9][0] ) );
  DFFPOSX1 \opcode_reg[10][1]  ( .D(n1059), .CLK(CLK), .Q(\opcode[10][1] ) );
  DFFPOSX1 \opcode_reg[10][0]  ( .D(n1058), .CLK(CLK), .Q(\opcode[10][0] ) );
  DFFPOSX1 \opcode_reg[11][1]  ( .D(n1057), .CLK(CLK), .Q(\opcode[11][1] ) );
  DFFPOSX1 \opcode_reg[11][0]  ( .D(n1056), .CLK(CLK), .Q(\opcode[11][0] ) );
  DFFPOSX1 \opcode_reg[12][1]  ( .D(n929), .CLK(CLK), .Q(\opcode[12][1] ) );
  DFFPOSX1 \opcode_reg[12][0]  ( .D(n930), .CLK(CLK), .Q(\opcode[12][0] ) );
  DFFPOSX1 \opcode_reg[13][1]  ( .D(n927), .CLK(CLK), .Q(\opcode[13][1] ) );
  DFFPOSX1 \opcode_reg[13][0]  ( .D(n928), .CLK(CLK), .Q(\opcode[13][0] ) );
  DFFPOSX1 \opcode_reg[14][1]  ( .D(n925), .CLK(CLK), .Q(\opcode[14][1] ) );
  DFFPOSX1 \opcode_reg[14][0]  ( .D(n926), .CLK(CLK), .Q(\opcode[14][0] ) );
  DFFPOSX1 \opcode_reg[15][1]  ( .D(n923), .CLK(CLK), .Q(\opcode[15][1] ) );
  DFFPOSX1 \opcode_reg[15][0]  ( .D(n924), .CLK(CLK), .Q(\opcode[15][0] ) );
  DFFPOSX1 \opcode_reg[16][1]  ( .D(n1055), .CLK(CLK), .Q(\opcode[16][1] ) );
  DFFPOSX1 \opcode_reg[16][0]  ( .D(n1054), .CLK(CLK), .Q(\opcode[16][0] ) );
  DFFPOSX1 \opcode_reg[17][1]  ( .D(n1053), .CLK(CLK), .Q(\opcode[17][1] ) );
  DFFPOSX1 \opcode_reg[17][0]  ( .D(n1052), .CLK(CLK), .Q(\opcode[17][0] ) );
  DFFPOSX1 \opcode_reg[18][1]  ( .D(n1051), .CLK(CLK), .Q(\opcode[18][1] ) );
  DFFPOSX1 \opcode_reg[18][0]  ( .D(n1050), .CLK(CLK), .Q(\opcode[18][0] ) );
  DFFPOSX1 \opcode_reg[19][1]  ( .D(n1049), .CLK(CLK), .Q(\opcode[19][1] ) );
  DFFPOSX1 \opcode_reg[19][0]  ( .D(n1048), .CLK(CLK), .Q(\opcode[19][0] ) );
  DFFPOSX1 \opcode_reg[20][1]  ( .D(n921), .CLK(CLK), .Q(\opcode[20][1] ) );
  DFFPOSX1 \opcode_reg[20][0]  ( .D(n922), .CLK(CLK), .Q(\opcode[20][0] ) );
  DFFPOSX1 \opcode_reg[21][1]  ( .D(n919), .CLK(CLK), .Q(\opcode[21][1] ) );
  DFFPOSX1 \opcode_reg[21][0]  ( .D(n920), .CLK(CLK), .Q(\opcode[21][0] ) );
  DFFPOSX1 \opcode_reg[22][1]  ( .D(n917), .CLK(CLK), .Q(\opcode[22][1] ) );
  DFFPOSX1 \opcode_reg[22][0]  ( .D(n918), .CLK(CLK), .Q(\opcode[22][0] ) );
  DFFPOSX1 \opcode_reg[23][1]  ( .D(n915), .CLK(CLK), .Q(\opcode[23][1] ) );
  DFFPOSX1 \opcode_reg[23][0]  ( .D(n916), .CLK(CLK), .Q(\opcode[23][0] ) );
  DFFPOSX1 \opcode_reg[24][1]  ( .D(n913), .CLK(CLK), .Q(\opcode[24][1] ) );
  DFFPOSX1 \opcode_reg[24][0]  ( .D(n914), .CLK(CLK), .Q(\opcode[24][0] ) );
  DFFPOSX1 \opcode_reg[25][1]  ( .D(n911), .CLK(CLK), .Q(\opcode[25][1] ) );
  DFFPOSX1 \opcode_reg[25][0]  ( .D(n912), .CLK(CLK), .Q(\opcode[25][0] ) );
  DFFPOSX1 \opcode_reg[26][1]  ( .D(n909), .CLK(CLK), .Q(\opcode[26][1] ) );
  DFFPOSX1 \opcode_reg[26][0]  ( .D(n910), .CLK(CLK), .Q(\opcode[26][0] ) );
  DFFPOSX1 \opcode_reg[27][1]  ( .D(n866), .CLK(CLK), .Q(\opcode[27][1] ) );
  DFFPOSX1 \opcode_reg[27][0]  ( .D(n867), .CLK(CLK), .Q(\opcode[27][0] ) );
  DFFPOSX1 \opcode_reg[28][1]  ( .D(n1047), .CLK(CLK), .Q(\opcode[28][1] ) );
  DFFPOSX1 \opcode_reg[28][0]  ( .D(n1046), .CLK(CLK), .Q(\opcode[28][0] ) );
  DFFPOSX1 \opcode_reg[29][1]  ( .D(n1045), .CLK(CLK), .Q(\opcode[29][1] ) );
  DFFPOSX1 \opcode_reg[29][0]  ( .D(n1044), .CLK(CLK), .Q(\opcode[29][0] ) );
  DFFPOSX1 \opcode_reg[30][1]  ( .D(n1043), .CLK(CLK), .Q(\opcode[30][1] ) );
  DFFPOSX1 \opcode_reg[30][0]  ( .D(n1042), .CLK(CLK), .Q(\opcode[30][0] ) );
  DFFPOSX1 \opcode_reg[31][1]  ( .D(n1041), .CLK(CLK), .Q(\opcode[31][1] ) );
  DFFPOSX1 \opcode_reg[31][0]  ( .D(n1040), .CLK(CLK), .Q(\opcode[31][0] ) );
  DFFPOSX1 \DATA_reg[7]  ( .D(n1039), .CLK(CLK), .Q(DATA[7]) );
  DFFPOSX1 \DATA_reg[6]  ( .D(n1038), .CLK(CLK), .Q(DATA[6]) );
  DFFPOSX1 \DATA_reg[5]  ( .D(n1037), .CLK(CLK), .Q(DATA[5]) );
  DFFPOSX1 \DATA_reg[4]  ( .D(n1036), .CLK(CLK), .Q(DATA[4]) );
  DFFPOSX1 \DATA_reg[3]  ( .D(n1035), .CLK(CLK), .Q(DATA[3]) );
  DFFPOSX1 \DATA_reg[2]  ( .D(n1034), .CLK(CLK), .Q(DATA[2]) );
  DFFPOSX1 \DATA_reg[1]  ( .D(n1033), .CLK(CLK), .Q(DATA[1]) );
  DFFPOSX1 \DATA_reg[0]  ( .D(n1032), .CLK(CLK), .Q(DATA[0]) );
  DFFPOSX1 \OUT_OPCODE_reg[1]  ( .D(n1031), .CLK(CLK), .Q(OUT_OPCODE[1]) );
  DFFPOSX1 \OUT_OPCODE_reg[0]  ( .D(n1030), .CLK(CLK), .Q(OUT_OPCODE[0]) );
  DFFPOSX1 EMPTY_reg ( .D(n1198), .CLK(CLK), .Q(EMPTY) );
  FAX1 \sub_72/U2_1  ( .A(n67), .B(n514), .C(\sub_72/carry[1] ), .YC(
        \sub_72/carry[2] ), .YS(N190) );
  FAX1 \sub_72/U2_2  ( .A(n65), .B(n851), .C(\sub_72/carry[2] ), .YC(
        \sub_72/carry[3] ), .YS(N191) );
  FAX1 \sub_72/U2_3  ( .A(n71), .B(n821), .C(\sub_72/carry[3] ), .YC(
        \sub_72/carry[4] ), .YS(N192) );
  FAX1 \sub_72/U2_4  ( .A(writeptr[4]), .B(n842), .C(\sub_72/carry[4] ), .YS(
        N193) );
  HAX1 \add_67/U1_1_1  ( .A(n67), .B(n69), .YC(\add_67/carry[2] ), .YS(N48) );
  HAX1 \add_67/U1_1_2  ( .A(n65), .B(\add_67/carry[2] ), .YC(\add_67/carry[3] ), .YS(N49) );
  HAX1 \add_67/U1_1_3  ( .A(n71), .B(\add_67/carry[3] ), .YC(\add_67/carry[4] ), .YS(N50) );
  HAX1 \r83/U1_1_1  ( .A(writeptr[1]), .B(writeptr[0]), .YC(\r83/carry[2] ), 
        .YS(N32) );
  HAX1 \r83/U1_1_2  ( .A(writeptr[2]), .B(\r83/carry[2] ), .YC(\r83/carry[3] ), 
        .YS(N33) );
  HAX1 \r83/U1_1_3  ( .A(writeptr[3]), .B(\r83/carry[3] ), .YC(\r83/carry[4] ), 
        .YS(N34) );
  DFFSR \BYTE_COUNT_reg[0]  ( .D(N338), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        BYTE_COUNT[0]) );
  DFFSR \BYTE_COUNT_reg[1]  ( .D(N339), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        BYTE_COUNT[1]) );
  DFFSR \BYTE_COUNT_reg[2]  ( .D(N340), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        BYTE_COUNT[2]) );
  DFFSR \readptr_reg[0]  ( .D(N343), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        readptr[0]) );
  DFFSR \BYTE_COUNT_reg[3]  ( .D(N341), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        BYTE_COUNT[3]) );
  DFFSR \readptr_reg[1]  ( .D(N344), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        readptr[1]) );
  DFFSR \BYTE_COUNT_reg[4]  ( .D(N342), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        BYTE_COUNT[4]) );
  DFFSR \readptr_reg[2]  ( .D(N345), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        readptr[2]) );
  DFFSR \readptr_reg[3]  ( .D(N346), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        readptr[3]) );
  DFFSR \writeptr_reg[4]  ( .D(n862), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        writeptr[4]) );
  DFFSR \writeptr_reg[3]  ( .D(n860), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        writeptr[3]) );
  DFFSR \writeptr_reg[2]  ( .D(n854), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        writeptr[2]) );
  DFFSR \writeptr_reg[1]  ( .D(n856), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        writeptr[1]) );
  DFFSR \writeptr_reg[0]  ( .D(n858), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        writeptr[0]) );
  DFFSR \readptr_reg[4]  ( .D(N347), .CLK(CLK), .R(n85), .S(1'b1), .Q(
        readptr[4]) );
  BUFX2 U3 ( .A(n351), .Y(n63) );
  BUFX2 U4 ( .A(n277), .Y(n20) );
  BUFX2 U5 ( .A(n449), .Y(n62) );
  INVX2 U6 ( .A(n34), .Y(n61) );
  INVX2 U7 ( .A(n33), .Y(n45) );
  BUFX2 U8 ( .A(n116), .Y(n46) );
  INVX4 U9 ( .A(n26), .Y(n121) );
  INVX2 U10 ( .A(n27), .Y(n47) );
  INVX2 U11 ( .A(n28), .Y(n48) );
  INVX2 U12 ( .A(n29), .Y(n60) );
  INVX2 U13 ( .A(n30), .Y(n59) );
  INVX2 U14 ( .A(n31), .Y(n58) );
  INVX2 U15 ( .A(n32), .Y(n57) );
  INVX2 U16 ( .A(n35), .Y(n53) );
  INVX2 U17 ( .A(n36), .Y(n54) );
  INVX2 U18 ( .A(n40), .Y(n55) );
  INVX2 U19 ( .A(n41), .Y(n56) );
  INVX2 U20 ( .A(n39), .Y(n52) );
  INVX2 U21 ( .A(n37), .Y(n51) );
  INVX2 U22 ( .A(n2), .Y(n50) );
  INVX2 U23 ( .A(n38), .Y(n49) );
  AND2X2 U24 ( .A(n493), .B(n70), .Y(n1) );
  OR2X2 U25 ( .A(n19), .B(n134), .Y(n2) );
  AND2X2 U26 ( .A(n493), .B(n71), .Y(n3) );
  INVX2 U42 ( .A(n146), .Y(n309) );
  NAND2X1 U43 ( .A(n63), .B(n3), .Y(n174) );
  NAND2X1 U44 ( .A(n63), .B(n1), .Y(n209) );
  BUFX2 U45 ( .A(n277), .Y(n19) );
  INVX2 U46 ( .A(n135), .Y(n126) );
  INVX2 U47 ( .A(writeptr[0]), .Y(n68) );
  INVX2 U48 ( .A(writeptr[1]), .Y(n66) );
  OR2X2 U49 ( .A(n145), .B(n174), .Y(n21) );
  INVX4 U50 ( .A(n21), .Y(n458) );
  OR2X2 U51 ( .A(n134), .B(n174), .Y(n22) );
  INVX4 U52 ( .A(n22), .Y(n106) );
  OR2X2 U53 ( .A(n184), .B(n174), .Y(n23) );
  INVX4 U54 ( .A(n23), .Y(n101) );
  OR2X2 U55 ( .A(n140), .B(n174), .Y(n24) );
  INVX4 U56 ( .A(n24), .Y(n111) );
  OR2X2 U57 ( .A(n235), .B(n174), .Y(n25) );
  INVX4 U58 ( .A(n25), .Y(n432) );
  OR2X2 U59 ( .A(n151), .B(n209), .Y(n26) );
  OR2X2 U60 ( .A(n209), .B(n226), .Y(n27) );
  OR2X2 U61 ( .A(n209), .B(n235), .Y(n28) );
  OR2X2 U62 ( .A(n209), .B(n175), .Y(n29) );
  OR2X2 U63 ( .A(n209), .B(n184), .Y(n30) );
  OR2X2 U64 ( .A(n209), .B(n134), .Y(n31) );
  OR2X2 U65 ( .A(n209), .B(n140), .Y(n32) );
  OR2X2 U66 ( .A(n174), .B(n175), .Y(n33) );
  OR2X2 U67 ( .A(n174), .B(n226), .Y(n34) );
  INVX2 U68 ( .A(RCV_OPCODE[0]), .Y(n76) );
  OR2X2 U69 ( .A(n20), .B(n145), .Y(n35) );
  OR2X2 U70 ( .A(n20), .B(n151), .Y(n36) );
  INVX2 U71 ( .A(n500), .Y(n96) );
  XNOR2X1 U72 ( .A(readptr[0]), .B(n69), .Y(n516) );
  OR2X2 U73 ( .A(n19), .B(n184), .Y(n37) );
  OR2X2 U74 ( .A(n19), .B(n140), .Y(n38) );
  OR2X2 U75 ( .A(n20), .B(n175), .Y(n39) );
  OR2X2 U76 ( .A(n20), .B(n226), .Y(n40) );
  OR2X2 U77 ( .A(n20), .B(n235), .Y(n41) );
  INVX2 U78 ( .A(RST), .Y(n85) );
  INVX2 U79 ( .A(n508), .Y(n156) );
  INVX2 U80 ( .A(n68), .Y(n69) );
  INVX2 U81 ( .A(n66), .Y(n67) );
  INVX2 U82 ( .A(n70), .Y(n71) );
  INVX2 U83 ( .A(n64), .Y(n65) );
  INVX2 U84 ( .A(RCV_DATA[7]), .Y(n77) );
  INVX2 U85 ( .A(RCV_DATA[1]), .Y(n83) );
  INVX2 U86 ( .A(RCV_DATA[3]), .Y(n81) );
  INVX2 U87 ( .A(RCV_DATA[5]), .Y(n79) );
  INVX2 U88 ( .A(RCV_DATA[0]), .Y(n84) );
  INVX2 U89 ( .A(RCV_DATA[2]), .Y(n82) );
  INVX2 U90 ( .A(RCV_DATA[4]), .Y(n80) );
  INVX2 U91 ( .A(RCV_DATA[6]), .Y(n78) );
  XNOR2X1 U92 ( .A(readptr[4]), .B(n42), .Y(n513) );
  XNOR2X1 U93 ( .A(\r83/carry[4] ), .B(writeptr[4]), .Y(n42) );
  INVX2 U94 ( .A(writeptr[2]), .Y(n64) );
  INVX2 U95 ( .A(writeptr[3]), .Y(n70) );
  BUFX2 U96 ( .A(state), .Y(n72) );
  INVX2 U97 ( .A(RCV_OPCODE[0]), .Y(n93) );
  INVX2 U98 ( .A(n507), .Y(n353) );
  INVX1 U99 ( .A(n63), .Y(n43) );
  INVX2 U100 ( .A(n43), .Y(n44) );
  AND2X2 U101 ( .A(n475), .B(n63), .Y(n244) );
  INVX1 U102 ( .A(RCV_OPCODE[1]), .Y(n73) );
  INVX1 U103 ( .A(RCV_OPCODE[1]), .Y(n74) );
  AND2X2 U104 ( .A(RCV_OPCODE[1]), .B(RCV_OPCODE[0]), .Y(n480) );
  INVX1 U105 ( .A(RCV_OPCODE[1]), .Y(n75) );
  AND2X2 U106 ( .A(n480), .B(n353), .Y(n356) );
  AND2X2 U107 ( .A(n815), .B(n817), .Y(n534) );
  AND2X2 U108 ( .A(n813), .B(n817), .Y(n533) );
  AND2X2 U109 ( .A(n815), .B(n818), .Y(n536) );
  AND2X2 U110 ( .A(n813), .B(n818), .Y(n535) );
  AND2X2 U111 ( .A(n829), .B(n817), .Y(n547) );
  AND2X2 U112 ( .A(n817), .B(n828), .Y(n546) );
  AND2X2 U113 ( .A(n818), .B(n829), .Y(n549) );
  AND2X2 U114 ( .A(n818), .B(n828), .Y(n548) );
  AND2X2 U115 ( .A(n840), .B(n818), .Y(n562) );
  AND2X2 U116 ( .A(n839), .B(n818), .Y(n561) );
  AND2X2 U117 ( .A(n840), .B(n817), .Y(n564) );
  AND2X2 U118 ( .A(n839), .B(n817), .Y(n563) );
  AND2X2 U119 ( .A(n850), .B(n817), .Y(n575) );
  AND2X2 U120 ( .A(n849), .B(n817), .Y(n574) );
  AND2X2 U121 ( .A(n850), .B(n818), .Y(n577) );
  AND2X2 U122 ( .A(n849), .B(n818), .Y(n576) );
  OR2X1 U123 ( .A(n820), .B(n69), .Y(\sub_72/carry[1] ) );
  XNOR2X1 U124 ( .A(n69), .B(n820), .Y(N189) );
  XOR2X1 U125 ( .A(readptr[4]), .B(\add_76_aco/carry[4] ), .Y(N337) );
  AND2X1 U126 ( .A(readptr[3]), .B(\add_76_aco/carry[3] ), .Y(
        \add_76_aco/carry[4] ) );
  XOR2X1 U127 ( .A(\add_76_aco/carry[3] ), .B(readptr[3]), .Y(N336) );
  AND2X1 U128 ( .A(readptr[2]), .B(\add_76_aco/carry[2] ), .Y(
        \add_76_aco/carry[3] ) );
  XOR2X1 U129 ( .A(\add_76_aco/carry[2] ), .B(readptr[2]), .Y(N335) );
  AND2X1 U130 ( .A(readptr[1]), .B(\add_76_aco/carry[1] ), .Y(
        \add_76_aco/carry[2] ) );
  XOR2X1 U131 ( .A(\add_76_aco/carry[1] ), .B(readptr[1]), .Y(N334) );
  AND2X1 U132 ( .A(readptr[0]), .B(N195), .Y(\add_76_aco/carry[1] ) );
  XOR2X1 U133 ( .A(N195), .B(readptr[0]), .Y(N333) );
  NOR2X1 U134 ( .A(n67), .B(n69), .Y(n87) );
  AOI21X1 U135 ( .A(n69), .B(n67), .C(n87), .Y(n86) );
  NAND2X1 U136 ( .A(n87), .B(n64), .Y(n88) );
  OAI21X1 U137 ( .A(n87), .B(n64), .C(n88), .Y(N44) );
  XNOR2X1 U138 ( .A(n71), .B(n88), .Y(N45) );
  NOR2X1 U139 ( .A(n71), .B(n88), .Y(n89) );
  XOR2X1 U140 ( .A(writeptr[4]), .B(n89), .Y(N46) );
  INVX2 U141 ( .A(n86), .Y(N43) );
  XOR2X1 U142 ( .A(\add_67/carry[4] ), .B(writeptr[4]), .Y(N51) );
  MUX2X1 U143 ( .B(n74), .A(n91), .S(n92), .Y(n866) );
  MUX2X1 U144 ( .B(n76), .A(n94), .S(n92), .Y(n867) );
  AOI21X1 U145 ( .A(n95), .B(n96), .C(n45), .Y(n92) );
  MUX2X1 U146 ( .B(n73), .A(n97), .S(n98), .Y(n909) );
  MUX2X1 U147 ( .B(n76), .A(n99), .S(n98), .Y(n910) );
  AOI21X1 U148 ( .A(n96), .B(n100), .C(n101), .Y(n98) );
  MUX2X1 U149 ( .B(n73), .A(n102), .S(n103), .Y(n911) );
  MUX2X1 U150 ( .B(n76), .A(n104), .S(n103), .Y(n912) );
  AOI21X1 U151 ( .A(n96), .B(n105), .C(n106), .Y(n103) );
  MUX2X1 U152 ( .B(n73), .A(n107), .S(n108), .Y(n913) );
  MUX2X1 U153 ( .B(n76), .A(n109), .S(n108), .Y(n914) );
  AOI21X1 U154 ( .A(n96), .B(n110), .C(n111), .Y(n108) );
  MUX2X1 U155 ( .B(n73), .A(n112), .S(n113), .Y(n915) );
  INVX1 U156 ( .A(\opcode[23][1] ), .Y(n112) );
  MUX2X1 U157 ( .B(n76), .A(n114), .S(n113), .Y(n916) );
  AOI21X1 U158 ( .A(n96), .B(n115), .C(n46), .Y(n113) );
  INVX1 U159 ( .A(\opcode[23][0] ), .Y(n114) );
  MUX2X1 U160 ( .B(n73), .A(n117), .S(n118), .Y(n917) );
  INVX1 U161 ( .A(\opcode[22][1] ), .Y(n117) );
  MUX2X1 U162 ( .B(n76), .A(n119), .S(n118), .Y(n918) );
  AOI21X1 U163 ( .A(n96), .B(n120), .C(n121), .Y(n118) );
  INVX1 U164 ( .A(\opcode[22][0] ), .Y(n119) );
  MUX2X1 U165 ( .B(n73), .A(n122), .S(n123), .Y(n919) );
  INVX1 U166 ( .A(\opcode[21][1] ), .Y(n122) );
  MUX2X1 U167 ( .B(n76), .A(n124), .S(n123), .Y(n920) );
  AOI21X1 U168 ( .A(n125), .B(n126), .C(n47), .Y(n123) );
  INVX1 U169 ( .A(\opcode[21][0] ), .Y(n124) );
  MUX2X1 U170 ( .B(n73), .A(n127), .S(n128), .Y(n921) );
  INVX1 U171 ( .A(\opcode[20][1] ), .Y(n127) );
  MUX2X1 U172 ( .B(n76), .A(n129), .S(n128), .Y(n922) );
  AOI21X1 U173 ( .A(n130), .B(n126), .C(n48), .Y(n128) );
  INVX1 U174 ( .A(\opcode[20][0] ), .Y(n129) );
  INVX1 U175 ( .A(n131), .Y(n923) );
  MUX2X1 U176 ( .B(\opcode[15][1] ), .A(RCV_OPCODE[1]), .S(n132), .Y(n131) );
  INVX1 U177 ( .A(n133), .Y(n924) );
  MUX2X1 U178 ( .B(\opcode[15][0] ), .A(RCV_OPCODE[0]), .S(n132), .Y(n133) );
  OAI21X1 U179 ( .A(n134), .B(n135), .C(n136), .Y(n132) );
  INVX1 U180 ( .A(n137), .Y(n925) );
  MUX2X1 U181 ( .B(\opcode[14][1] ), .A(RCV_OPCODE[1]), .S(n138), .Y(n137) );
  INVX1 U182 ( .A(n139), .Y(n926) );
  MUX2X1 U183 ( .B(\opcode[14][0] ), .A(RCV_OPCODE[0]), .S(n138), .Y(n139) );
  OAI21X1 U184 ( .A(n140), .B(n135), .C(n141), .Y(n138) );
  MUX2X1 U185 ( .B(n142), .A(n75), .S(n143), .Y(n927) );
  INVX1 U186 ( .A(\opcode[13][1] ), .Y(n142) );
  MUX2X1 U187 ( .B(n144), .A(n76), .S(n143), .Y(n928) );
  OAI21X1 U188 ( .A(n145), .B(n146), .C(n147), .Y(n143) );
  INVX1 U189 ( .A(\opcode[13][0] ), .Y(n144) );
  MUX2X1 U190 ( .B(n148), .A(n75), .S(n149), .Y(n929) );
  INVX1 U191 ( .A(\opcode[12][1] ), .Y(n148) );
  MUX2X1 U192 ( .B(n150), .A(n76), .S(n149), .Y(n930) );
  OAI21X1 U193 ( .A(n151), .B(n146), .C(n152), .Y(n149) );
  INVX1 U194 ( .A(\opcode[12][0] ), .Y(n150) );
  MUX2X1 U195 ( .B(n76), .A(n153), .S(n154), .Y(n931) );
  MUX2X1 U196 ( .B(n73), .A(n155), .S(n154), .Y(n932) );
  AOI21X1 U197 ( .A(n110), .B(n156), .C(n49), .Y(n154) );
  MUX2X1 U198 ( .B(n76), .A(n157), .S(n158), .Y(n933) );
  MUX2X1 U199 ( .B(n73), .A(n159), .S(n158), .Y(n934) );
  AOI21X1 U200 ( .A(n105), .B(n156), .C(n50), .Y(n158) );
  MUX2X1 U201 ( .B(n76), .A(n160), .S(n161), .Y(n935) );
  MUX2X1 U202 ( .B(n73), .A(n162), .S(n161), .Y(n936) );
  AOI21X1 U203 ( .A(n100), .B(n156), .C(n51), .Y(n161) );
  MUX2X1 U204 ( .B(n76), .A(n163), .S(n164), .Y(n937) );
  MUX2X1 U205 ( .B(n73), .A(n165), .S(n164), .Y(n938) );
  AOI21X1 U206 ( .A(n95), .B(n156), .C(n52), .Y(n164) );
  MUX2X1 U207 ( .B(n166), .A(n77), .S(n45), .Y(n939) );
  MUX2X1 U208 ( .B(n167), .A(n78), .S(n45), .Y(n940) );
  MUX2X1 U209 ( .B(n168), .A(n79), .S(n45), .Y(n941) );
  MUX2X1 U210 ( .B(n169), .A(n80), .S(n45), .Y(n942) );
  MUX2X1 U211 ( .B(n170), .A(n81), .S(n45), .Y(n943) );
  MUX2X1 U212 ( .B(n171), .A(n82), .S(n45), .Y(n944) );
  MUX2X1 U213 ( .B(n172), .A(n83), .S(n45), .Y(n945) );
  MUX2X1 U214 ( .B(n173), .A(n84), .S(n45), .Y(n946) );
  MUX2X1 U215 ( .B(n176), .A(n77), .S(n101), .Y(n947) );
  MUX2X1 U216 ( .B(n177), .A(n78), .S(n101), .Y(n948) );
  MUX2X1 U217 ( .B(n178), .A(n79), .S(n101), .Y(n949) );
  MUX2X1 U218 ( .B(n179), .A(n80), .S(n101), .Y(n950) );
  MUX2X1 U219 ( .B(n180), .A(n81), .S(n101), .Y(n951) );
  MUX2X1 U220 ( .B(n181), .A(n82), .S(n101), .Y(n952) );
  MUX2X1 U221 ( .B(n182), .A(n83), .S(n101), .Y(n953) );
  MUX2X1 U222 ( .B(n183), .A(n84), .S(n101), .Y(n954) );
  MUX2X1 U223 ( .B(n185), .A(n77), .S(n106), .Y(n955) );
  MUX2X1 U224 ( .B(n186), .A(n78), .S(n106), .Y(n956) );
  MUX2X1 U225 ( .B(n187), .A(n79), .S(n106), .Y(n957) );
  MUX2X1 U226 ( .B(n188), .A(n80), .S(n106), .Y(n958) );
  MUX2X1 U227 ( .B(n189), .A(n81), .S(n106), .Y(n959) );
  MUX2X1 U228 ( .B(n190), .A(n82), .S(n106), .Y(n960) );
  MUX2X1 U229 ( .B(n191), .A(n83), .S(n106), .Y(n961) );
  MUX2X1 U230 ( .B(n192), .A(n84), .S(n106), .Y(n962) );
  MUX2X1 U231 ( .B(n193), .A(n77), .S(n111), .Y(n963) );
  MUX2X1 U232 ( .B(n194), .A(n78), .S(n111), .Y(n964) );
  MUX2X1 U233 ( .B(n195), .A(n79), .S(n111), .Y(n965) );
  MUX2X1 U234 ( .B(n196), .A(n80), .S(n111), .Y(n966) );
  MUX2X1 U235 ( .B(n197), .A(n81), .S(n111), .Y(n967) );
  MUX2X1 U236 ( .B(n198), .A(n82), .S(n111), .Y(n968) );
  MUX2X1 U237 ( .B(n199), .A(n83), .S(n111), .Y(n969) );
  MUX2X1 U238 ( .B(n200), .A(n84), .S(n111), .Y(n970) );
  MUX2X1 U239 ( .B(n201), .A(n77), .S(n46), .Y(n971) );
  INVX1 U240 ( .A(\memory[23][7] ), .Y(n201) );
  MUX2X1 U241 ( .B(n202), .A(n78), .S(n46), .Y(n972) );
  INVX1 U242 ( .A(\memory[23][6] ), .Y(n202) );
  MUX2X1 U243 ( .B(n203), .A(n79), .S(n46), .Y(n973) );
  INVX1 U244 ( .A(\memory[23][5] ), .Y(n203) );
  MUX2X1 U245 ( .B(n204), .A(n80), .S(n46), .Y(n974) );
  INVX1 U246 ( .A(\memory[23][4] ), .Y(n204) );
  MUX2X1 U247 ( .B(n205), .A(n81), .S(n46), .Y(n975) );
  INVX1 U248 ( .A(\memory[23][3] ), .Y(n205) );
  MUX2X1 U249 ( .B(n206), .A(n82), .S(n46), .Y(n976) );
  INVX1 U250 ( .A(\memory[23][2] ), .Y(n206) );
  MUX2X1 U251 ( .B(n207), .A(n83), .S(n46), .Y(n977) );
  INVX1 U252 ( .A(\memory[23][1] ), .Y(n207) );
  MUX2X1 U253 ( .B(n208), .A(n84), .S(n46), .Y(n978) );
  NOR2X1 U254 ( .A(n145), .B(n209), .Y(n116) );
  INVX1 U255 ( .A(\memory[23][0] ), .Y(n208) );
  MUX2X1 U256 ( .B(n210), .A(n77), .S(n121), .Y(n979) );
  INVX1 U257 ( .A(\memory[22][7] ), .Y(n210) );
  MUX2X1 U258 ( .B(n211), .A(n78), .S(n121), .Y(n980) );
  INVX1 U259 ( .A(\memory[22][6] ), .Y(n211) );
  MUX2X1 U260 ( .B(n212), .A(n79), .S(n121), .Y(n981) );
  INVX1 U261 ( .A(\memory[22][5] ), .Y(n212) );
  MUX2X1 U262 ( .B(n213), .A(n80), .S(n121), .Y(n982) );
  INVX1 U263 ( .A(\memory[22][4] ), .Y(n213) );
  MUX2X1 U264 ( .B(n214), .A(n81), .S(n121), .Y(n983) );
  INVX1 U265 ( .A(\memory[22][3] ), .Y(n214) );
  MUX2X1 U266 ( .B(n215), .A(n82), .S(n121), .Y(n984) );
  INVX1 U267 ( .A(\memory[22][2] ), .Y(n215) );
  MUX2X1 U268 ( .B(n216), .A(n83), .S(n121), .Y(n985) );
  INVX1 U269 ( .A(\memory[22][1] ), .Y(n216) );
  MUX2X1 U270 ( .B(n217), .A(n84), .S(n121), .Y(n986) );
  INVX1 U271 ( .A(\memory[22][0] ), .Y(n217) );
  MUX2X1 U272 ( .B(n218), .A(n77), .S(n47), .Y(n987) );
  INVX1 U273 ( .A(\memory[21][7] ), .Y(n218) );
  MUX2X1 U274 ( .B(n219), .A(n78), .S(n47), .Y(n988) );
  INVX1 U275 ( .A(\memory[21][6] ), .Y(n219) );
  MUX2X1 U276 ( .B(n220), .A(n79), .S(n47), .Y(n989) );
  INVX1 U277 ( .A(\memory[21][5] ), .Y(n220) );
  MUX2X1 U278 ( .B(n221), .A(n80), .S(n47), .Y(n990) );
  INVX1 U279 ( .A(\memory[21][4] ), .Y(n221) );
  MUX2X1 U280 ( .B(n222), .A(n81), .S(n47), .Y(n991) );
  INVX1 U281 ( .A(\memory[21][3] ), .Y(n222) );
  MUX2X1 U282 ( .B(n223), .A(n82), .S(n47), .Y(n992) );
  INVX1 U283 ( .A(\memory[21][2] ), .Y(n223) );
  MUX2X1 U284 ( .B(n224), .A(n83), .S(n47), .Y(n993) );
  INVX1 U285 ( .A(\memory[21][1] ), .Y(n224) );
  MUX2X1 U286 ( .B(n225), .A(n84), .S(n47), .Y(n994) );
  INVX1 U287 ( .A(\memory[21][0] ), .Y(n225) );
  MUX2X1 U288 ( .B(n227), .A(n77), .S(n48), .Y(n995) );
  INVX1 U289 ( .A(\memory[20][7] ), .Y(n227) );
  MUX2X1 U290 ( .B(n228), .A(n78), .S(n48), .Y(n996) );
  INVX1 U291 ( .A(\memory[20][6] ), .Y(n228) );
  MUX2X1 U292 ( .B(n229), .A(n79), .S(n48), .Y(n997) );
  INVX1 U293 ( .A(\memory[20][5] ), .Y(n229) );
  MUX2X1 U294 ( .B(n230), .A(n80), .S(n48), .Y(n998) );
  INVX1 U295 ( .A(\memory[20][4] ), .Y(n230) );
  MUX2X1 U296 ( .B(n231), .A(n81), .S(n48), .Y(n999) );
  INVX1 U297 ( .A(\memory[20][3] ), .Y(n231) );
  MUX2X1 U298 ( .B(n232), .A(n82), .S(n48), .Y(n1000) );
  INVX1 U299 ( .A(\memory[20][2] ), .Y(n232) );
  MUX2X1 U300 ( .B(n233), .A(n83), .S(n48), .Y(n1001) );
  INVX1 U301 ( .A(\memory[20][1] ), .Y(n233) );
  MUX2X1 U302 ( .B(n234), .A(n84), .S(n48), .Y(n1002) );
  INVX1 U303 ( .A(\memory[20][0] ), .Y(n234) );
  MUX2X1 U304 ( .B(n77), .A(n236), .S(n136), .Y(n1003) );
  INVX1 U305 ( .A(\memory[15][7] ), .Y(n236) );
  MUX2X1 U306 ( .B(n78), .A(n237), .S(n136), .Y(n1004) );
  INVX1 U307 ( .A(\memory[15][6] ), .Y(n237) );
  MUX2X1 U308 ( .B(n79), .A(n238), .S(n136), .Y(n1005) );
  INVX1 U309 ( .A(\memory[15][5] ), .Y(n238) );
  MUX2X1 U310 ( .B(n80), .A(n239), .S(n136), .Y(n1006) );
  INVX1 U311 ( .A(\memory[15][4] ), .Y(n239) );
  MUX2X1 U312 ( .B(n81), .A(n240), .S(n136), .Y(n1007) );
  INVX1 U313 ( .A(\memory[15][3] ), .Y(n240) );
  MUX2X1 U314 ( .B(n82), .A(n241), .S(n136), .Y(n1008) );
  INVX1 U315 ( .A(\memory[15][2] ), .Y(n241) );
  MUX2X1 U316 ( .B(n83), .A(n242), .S(n136), .Y(n1009) );
  INVX1 U317 ( .A(\memory[15][1] ), .Y(n242) );
  MUX2X1 U318 ( .B(n84), .A(n243), .S(n136), .Y(n1010) );
  NAND2X1 U319 ( .A(n244), .B(n125), .Y(n136) );
  INVX1 U320 ( .A(\memory[15][0] ), .Y(n243) );
  MUX2X1 U321 ( .B(n77), .A(n245), .S(n141), .Y(n1011) );
  INVX1 U322 ( .A(\memory[14][7] ), .Y(n245) );
  MUX2X1 U323 ( .B(n78), .A(n246), .S(n141), .Y(n1012) );
  INVX1 U324 ( .A(\memory[14][6] ), .Y(n246) );
  MUX2X1 U325 ( .B(n79), .A(n247), .S(n141), .Y(n1013) );
  INVX1 U326 ( .A(\memory[14][5] ), .Y(n247) );
  MUX2X1 U327 ( .B(n80), .A(n248), .S(n141), .Y(n1014) );
  INVX1 U328 ( .A(\memory[14][4] ), .Y(n248) );
  MUX2X1 U329 ( .B(n81), .A(n249), .S(n141), .Y(n1015) );
  INVX1 U330 ( .A(\memory[14][3] ), .Y(n249) );
  MUX2X1 U331 ( .B(n82), .A(n250), .S(n141), .Y(n1016) );
  INVX1 U332 ( .A(\memory[14][2] ), .Y(n250) );
  MUX2X1 U333 ( .B(n83), .A(n251), .S(n141), .Y(n1017) );
  INVX1 U334 ( .A(\memory[14][1] ), .Y(n251) );
  MUX2X1 U335 ( .B(n84), .A(n252), .S(n141), .Y(n1018) );
  NAND2X1 U336 ( .A(n244), .B(n130), .Y(n141) );
  INVX1 U337 ( .A(\memory[14][0] ), .Y(n252) );
  MUX2X1 U338 ( .B(n77), .A(n253), .S(n147), .Y(n1019) );
  INVX1 U339 ( .A(\memory[13][7] ), .Y(n253) );
  MUX2X1 U340 ( .B(n78), .A(n254), .S(n147), .Y(n1020) );
  INVX1 U341 ( .A(\memory[13][6] ), .Y(n254) );
  MUX2X1 U342 ( .B(n79), .A(n255), .S(n147), .Y(n1021) );
  INVX1 U343 ( .A(\memory[13][5] ), .Y(n255) );
  MUX2X1 U344 ( .B(n80), .A(n256), .S(n147), .Y(n1022) );
  INVX1 U345 ( .A(\memory[13][4] ), .Y(n256) );
  MUX2X1 U346 ( .B(n81), .A(n257), .S(n147), .Y(n1023) );
  INVX1 U347 ( .A(\memory[13][3] ), .Y(n257) );
  MUX2X1 U348 ( .B(n82), .A(n258), .S(n147), .Y(n1024) );
  INVX1 U349 ( .A(\memory[13][2] ), .Y(n258) );
  MUX2X1 U350 ( .B(n83), .A(n259), .S(n147), .Y(n1025) );
  INVX1 U351 ( .A(\memory[13][1] ), .Y(n259) );
  MUX2X1 U352 ( .B(n84), .A(n260), .S(n147), .Y(n1026) );
  NAND2X1 U353 ( .A(n244), .B(n95), .Y(n147) );
  INVX1 U354 ( .A(\memory[13][0] ), .Y(n260) );
  MUX2X1 U355 ( .B(n77), .A(n261), .S(n152), .Y(n1027) );
  INVX1 U356 ( .A(\memory[12][7] ), .Y(n261) );
  MUX2X1 U357 ( .B(n78), .A(n262), .S(n152), .Y(n1028) );
  INVX1 U358 ( .A(\memory[12][6] ), .Y(n262) );
  MUX2X1 U359 ( .B(n79), .A(n263), .S(n152), .Y(n1029) );
  INVX1 U360 ( .A(\memory[12][5] ), .Y(n263) );
  MUX2X1 U361 ( .B(n80), .A(n264), .S(n152), .Y(n1064) );
  INVX1 U362 ( .A(\memory[12][4] ), .Y(n264) );
  MUX2X1 U363 ( .B(n81), .A(n265), .S(n152), .Y(n1065) );
  INVX1 U364 ( .A(\memory[12][3] ), .Y(n265) );
  MUX2X1 U365 ( .B(n82), .A(n266), .S(n152), .Y(n1066) );
  INVX1 U366 ( .A(\memory[12][2] ), .Y(n266) );
  MUX2X1 U367 ( .B(n83), .A(n267), .S(n152), .Y(n1067) );
  INVX1 U368 ( .A(\memory[12][1] ), .Y(n267) );
  MUX2X1 U369 ( .B(n84), .A(n268), .S(n152), .Y(n1068) );
  NAND2X1 U370 ( .A(n244), .B(n100), .Y(n152) );
  INVX1 U371 ( .A(\memory[12][0] ), .Y(n268) );
  MUX2X1 U372 ( .B(n269), .A(n84), .S(n49), .Y(n1069) );
  MUX2X1 U373 ( .B(n270), .A(n83), .S(n49), .Y(n1070) );
  MUX2X1 U374 ( .B(n271), .A(n82), .S(n49), .Y(n1071) );
  MUX2X1 U375 ( .B(n272), .A(n81), .S(n49), .Y(n1168) );
  MUX2X1 U376 ( .B(n273), .A(n80), .S(n49), .Y(n1169) );
  MUX2X1 U377 ( .B(n274), .A(n79), .S(n49), .Y(n1170) );
  MUX2X1 U378 ( .B(n275), .A(n78), .S(n49), .Y(n1171) );
  MUX2X1 U379 ( .B(n276), .A(n77), .S(n49), .Y(n1172) );
  MUX2X1 U380 ( .B(n278), .A(n84), .S(n50), .Y(n1173) );
  MUX2X1 U381 ( .B(n279), .A(n83), .S(n50), .Y(n1174) );
  MUX2X1 U382 ( .B(n280), .A(n82), .S(n50), .Y(n1175) );
  MUX2X1 U383 ( .B(n281), .A(n81), .S(n50), .Y(n1176) );
  MUX2X1 U384 ( .B(n282), .A(n80), .S(n50), .Y(n1177) );
  MUX2X1 U385 ( .B(n283), .A(n79), .S(n50), .Y(n1178) );
  MUX2X1 U386 ( .B(n284), .A(n78), .S(n50), .Y(n1179) );
  MUX2X1 U387 ( .B(n285), .A(n77), .S(n50), .Y(n1180) );
  MUX2X1 U388 ( .B(n286), .A(n84), .S(n51), .Y(n1181) );
  MUX2X1 U389 ( .B(n287), .A(n83), .S(n51), .Y(n1182) );
  MUX2X1 U390 ( .B(n288), .A(n82), .S(n51), .Y(n1183) );
  MUX2X1 U391 ( .B(n289), .A(n81), .S(n51), .Y(n1184) );
  MUX2X1 U392 ( .B(n290), .A(n80), .S(n51), .Y(n1185) );
  MUX2X1 U393 ( .B(n291), .A(n79), .S(n51), .Y(n1186) );
  MUX2X1 U394 ( .B(n292), .A(n78), .S(n51), .Y(n1187) );
  MUX2X1 U395 ( .B(n293), .A(n77), .S(n51), .Y(n1188) );
  MUX2X1 U396 ( .B(n294), .A(n84), .S(n52), .Y(n1189) );
  MUX2X1 U397 ( .B(n295), .A(n83), .S(n52), .Y(n1190) );
  MUX2X1 U398 ( .B(n296), .A(n82), .S(n52), .Y(n1191) );
  MUX2X1 U399 ( .B(n297), .A(n81), .S(n52), .Y(n1192) );
  MUX2X1 U400 ( .B(n298), .A(n80), .S(n52), .Y(n1193) );
  MUX2X1 U401 ( .B(n299), .A(n79), .S(n52), .Y(n1194) );
  MUX2X1 U402 ( .B(n300), .A(n78), .S(n52), .Y(n1195) );
  MUX2X1 U403 ( .B(n301), .A(n77), .S(n52), .Y(n1196) );
  MUX2X1 U404 ( .B(n302), .A(n303), .S(RST), .Y(n1197) );
  INVX1 U405 ( .A(FULL), .Y(n303) );
  MUX2X1 U406 ( .B(n304), .A(n305), .S(RST), .Y(n1198) );
  INVX1 U407 ( .A(EMPTY), .Y(n305) );
  MUX2X1 U408 ( .B(n76), .A(n306), .S(n307), .Y(n908) );
  INVX1 U409 ( .A(\opcode[7][0] ), .Y(n306) );
  MUX2X1 U410 ( .B(n73), .A(n308), .S(n307), .Y(n907) );
  AOI21X1 U411 ( .A(n115), .B(n309), .C(n53), .Y(n307) );
  INVX1 U412 ( .A(\opcode[7][1] ), .Y(n308) );
  MUX2X1 U413 ( .B(n310), .A(n84), .S(n53), .Y(n906) );
  INVX1 U414 ( .A(\memory[7][0] ), .Y(n310) );
  MUX2X1 U415 ( .B(n311), .A(n83), .S(n53), .Y(n905) );
  INVX1 U416 ( .A(\memory[7][1] ), .Y(n311) );
  MUX2X1 U417 ( .B(n312), .A(n82), .S(n53), .Y(n904) );
  INVX1 U418 ( .A(\memory[7][2] ), .Y(n312) );
  MUX2X1 U419 ( .B(n313), .A(n81), .S(n53), .Y(n903) );
  INVX1 U420 ( .A(\memory[7][3] ), .Y(n313) );
  MUX2X1 U421 ( .B(n314), .A(n80), .S(n53), .Y(n902) );
  INVX1 U422 ( .A(\memory[7][4] ), .Y(n314) );
  MUX2X1 U423 ( .B(n315), .A(n79), .S(n53), .Y(n901) );
  INVX1 U424 ( .A(\memory[7][5] ), .Y(n315) );
  MUX2X1 U425 ( .B(n316), .A(n78), .S(n53), .Y(n900) );
  INVX1 U426 ( .A(\memory[7][6] ), .Y(n316) );
  MUX2X1 U427 ( .B(n317), .A(n77), .S(n53), .Y(n899) );
  INVX1 U428 ( .A(\memory[7][7] ), .Y(n317) );
  MUX2X1 U429 ( .B(n76), .A(n318), .S(n319), .Y(n898) );
  INVX1 U430 ( .A(\opcode[6][0] ), .Y(n318) );
  MUX2X1 U431 ( .B(n74), .A(n320), .S(n319), .Y(n897) );
  AOI21X1 U432 ( .A(n120), .B(n309), .C(n54), .Y(n319) );
  INVX1 U433 ( .A(\opcode[6][1] ), .Y(n320) );
  MUX2X1 U434 ( .B(n321), .A(n84), .S(n54), .Y(n896) );
  INVX1 U435 ( .A(\memory[6][0] ), .Y(n321) );
  MUX2X1 U436 ( .B(n322), .A(n83), .S(n54), .Y(n895) );
  INVX1 U437 ( .A(\memory[6][1] ), .Y(n322) );
  MUX2X1 U438 ( .B(n323), .A(n82), .S(n54), .Y(n894) );
  INVX1 U439 ( .A(\memory[6][2] ), .Y(n323) );
  MUX2X1 U440 ( .B(n324), .A(n81), .S(n54), .Y(n893) );
  INVX1 U441 ( .A(\memory[6][3] ), .Y(n324) );
  MUX2X1 U442 ( .B(n325), .A(n80), .S(n54), .Y(n892) );
  INVX1 U443 ( .A(\memory[6][4] ), .Y(n325) );
  MUX2X1 U444 ( .B(n326), .A(n79), .S(n54), .Y(n891) );
  INVX1 U445 ( .A(\memory[6][5] ), .Y(n326) );
  MUX2X1 U446 ( .B(n327), .A(n78), .S(n54), .Y(n890) );
  INVX1 U447 ( .A(\memory[6][6] ), .Y(n327) );
  MUX2X1 U448 ( .B(n328), .A(n77), .S(n54), .Y(n889) );
  INVX1 U449 ( .A(\memory[6][7] ), .Y(n328) );
  MUX2X1 U450 ( .B(n93), .A(n329), .S(n330), .Y(n888) );
  INVX1 U451 ( .A(\opcode[5][0] ), .Y(n329) );
  MUX2X1 U452 ( .B(n74), .A(n331), .S(n330), .Y(n887) );
  AOI21X1 U453 ( .A(n125), .B(n156), .C(n55), .Y(n330) );
  INVX1 U454 ( .A(\opcode[5][1] ), .Y(n331) );
  MUX2X1 U455 ( .B(n332), .A(n84), .S(n55), .Y(n886) );
  INVX1 U456 ( .A(\memory[5][0] ), .Y(n332) );
  MUX2X1 U457 ( .B(n333), .A(n83), .S(n55), .Y(n885) );
  INVX1 U458 ( .A(\memory[5][1] ), .Y(n333) );
  MUX2X1 U459 ( .B(n334), .A(n82), .S(n55), .Y(n884) );
  INVX1 U460 ( .A(\memory[5][2] ), .Y(n334) );
  MUX2X1 U461 ( .B(n335), .A(n81), .S(n55), .Y(n883) );
  INVX1 U462 ( .A(\memory[5][3] ), .Y(n335) );
  MUX2X1 U463 ( .B(n336), .A(n80), .S(n55), .Y(n882) );
  INVX1 U464 ( .A(\memory[5][4] ), .Y(n336) );
  MUX2X1 U465 ( .B(n337), .A(n79), .S(n55), .Y(n881) );
  INVX1 U466 ( .A(\memory[5][5] ), .Y(n337) );
  MUX2X1 U467 ( .B(n338), .A(n78), .S(n55), .Y(n880) );
  INVX1 U468 ( .A(\memory[5][6] ), .Y(n338) );
  MUX2X1 U469 ( .B(n339), .A(n77), .S(n55), .Y(n879) );
  INVX1 U470 ( .A(\memory[5][7] ), .Y(n339) );
  MUX2X1 U471 ( .B(n76), .A(n340), .S(n341), .Y(n878) );
  INVX1 U472 ( .A(\opcode[4][0] ), .Y(n340) );
  MUX2X1 U473 ( .B(n74), .A(n342), .S(n341), .Y(n877) );
  AOI21X1 U474 ( .A(n130), .B(n156), .C(n56), .Y(n341) );
  INVX1 U475 ( .A(\opcode[4][1] ), .Y(n342) );
  MUX2X1 U476 ( .B(n343), .A(n84), .S(n56), .Y(n876) );
  INVX1 U477 ( .A(\memory[4][0] ), .Y(n343) );
  MUX2X1 U478 ( .B(n344), .A(n83), .S(n56), .Y(n875) );
  INVX1 U479 ( .A(\memory[4][1] ), .Y(n344) );
  MUX2X1 U480 ( .B(n345), .A(n82), .S(n56), .Y(n874) );
  INVX1 U481 ( .A(\memory[4][2] ), .Y(n345) );
  MUX2X1 U482 ( .B(n346), .A(n81), .S(n56), .Y(n873) );
  INVX1 U483 ( .A(\memory[4][3] ), .Y(n346) );
  MUX2X1 U484 ( .B(n347), .A(n80), .S(n56), .Y(n872) );
  INVX1 U485 ( .A(\memory[4][4] ), .Y(n347) );
  MUX2X1 U486 ( .B(n348), .A(n79), .S(n56), .Y(n871) );
  INVX1 U487 ( .A(\memory[4][5] ), .Y(n348) );
  MUX2X1 U488 ( .B(n349), .A(n78), .S(n56), .Y(n870) );
  INVX1 U489 ( .A(\memory[4][6] ), .Y(n349) );
  MUX2X1 U490 ( .B(n350), .A(n77), .S(n56), .Y(n869) );
  NAND3X1 U491 ( .A(n63), .B(n70), .C(n352), .Y(n277) );
  INVX1 U492 ( .A(\memory[4][7] ), .Y(n350) );
  OAI21X1 U493 ( .A(n353), .B(n354), .C(n355), .Y(n862) );
  AOI22X1 U494 ( .A(N51), .B(n44), .C(N46), .D(n356), .Y(n355) );
  OAI21X1 U495 ( .A(n353), .B(n70), .C(n357), .Y(n860) );
  AOI22X1 U496 ( .A(N50), .B(n44), .C(N45), .D(n356), .Y(n357) );
  OAI21X1 U497 ( .A(n353), .B(n358), .C(n359), .Y(n858) );
  AOI22X1 U498 ( .A(n358), .B(n44), .C(n358), .D(n356), .Y(n359) );
  OAI21X1 U499 ( .A(n353), .B(n360), .C(n361), .Y(n856) );
  AOI22X1 U500 ( .A(N48), .B(n44), .C(N43), .D(n356), .Y(n361) );
  OAI21X1 U501 ( .A(n353), .B(n64), .C(n362), .Y(n854) );
  AOI22X1 U502 ( .A(N49), .B(n44), .C(N44), .D(n356), .Y(n362) );
  MUX2X1 U503 ( .B(n77), .A(n363), .S(n364), .Y(n1167) );
  MUX2X1 U504 ( .B(n78), .A(n365), .S(n364), .Y(n1166) );
  MUX2X1 U505 ( .B(n79), .A(n366), .S(n364), .Y(n1165) );
  MUX2X1 U506 ( .B(n80), .A(n367), .S(n364), .Y(n1164) );
  MUX2X1 U507 ( .B(n81), .A(n368), .S(n364), .Y(n1163) );
  MUX2X1 U508 ( .B(n82), .A(n369), .S(n364), .Y(n1162) );
  MUX2X1 U509 ( .B(n83), .A(n370), .S(n364), .Y(n1161) );
  MUX2X1 U510 ( .B(n84), .A(n371), .S(n364), .Y(n1160) );
  MUX2X1 U511 ( .B(n77), .A(n372), .S(n373), .Y(n1159) );
  MUX2X1 U512 ( .B(n78), .A(n374), .S(n373), .Y(n1158) );
  MUX2X1 U513 ( .B(n79), .A(n375), .S(n373), .Y(n1157) );
  MUX2X1 U514 ( .B(n80), .A(n376), .S(n373), .Y(n1156) );
  MUX2X1 U515 ( .B(n81), .A(n377), .S(n373), .Y(n1155) );
  MUX2X1 U516 ( .B(n82), .A(n378), .S(n373), .Y(n1154) );
  MUX2X1 U517 ( .B(n83), .A(n379), .S(n373), .Y(n1153) );
  MUX2X1 U518 ( .B(n84), .A(n380), .S(n373), .Y(n1152) );
  MUX2X1 U519 ( .B(n77), .A(n381), .S(n382), .Y(n1151) );
  MUX2X1 U520 ( .B(n78), .A(n383), .S(n382), .Y(n1150) );
  MUX2X1 U521 ( .B(n79), .A(n384), .S(n382), .Y(n1149) );
  MUX2X1 U522 ( .B(n80), .A(n385), .S(n382), .Y(n1148) );
  MUX2X1 U523 ( .B(n81), .A(n386), .S(n382), .Y(n1147) );
  MUX2X1 U524 ( .B(n82), .A(n387), .S(n382), .Y(n1146) );
  MUX2X1 U525 ( .B(n83), .A(n388), .S(n382), .Y(n1145) );
  MUX2X1 U526 ( .B(n84), .A(n389), .S(n382), .Y(n1144) );
  MUX2X1 U527 ( .B(n390), .A(n77), .S(n391), .Y(n1143) );
  MUX2X1 U528 ( .B(n392), .A(n78), .S(n391), .Y(n1142) );
  MUX2X1 U529 ( .B(n393), .A(n79), .S(n391), .Y(n1141) );
  MUX2X1 U530 ( .B(n394), .A(n80), .S(n391), .Y(n1140) );
  MUX2X1 U531 ( .B(n395), .A(n81), .S(n391), .Y(n1139) );
  MUX2X1 U532 ( .B(n396), .A(n82), .S(n391), .Y(n1138) );
  MUX2X1 U533 ( .B(n397), .A(n83), .S(n391), .Y(n1137) );
  MUX2X1 U534 ( .B(n398), .A(n84), .S(n391), .Y(n1136) );
  AND2X1 U535 ( .A(n244), .B(n105), .Y(n391) );
  MUX2X1 U536 ( .B(n399), .A(n77), .S(n57), .Y(n1135) );
  MUX2X1 U537 ( .B(n400), .A(n78), .S(n57), .Y(n1134) );
  MUX2X1 U538 ( .B(n401), .A(n79), .S(n57), .Y(n1133) );
  MUX2X1 U539 ( .B(n402), .A(n80), .S(n57), .Y(n1132) );
  MUX2X1 U540 ( .B(n403), .A(n81), .S(n57), .Y(n1131) );
  MUX2X1 U541 ( .B(n404), .A(n82), .S(n57), .Y(n1130) );
  MUX2X1 U542 ( .B(n405), .A(n83), .S(n57), .Y(n1129) );
  MUX2X1 U543 ( .B(n406), .A(n84), .S(n57), .Y(n1128) );
  MUX2X1 U544 ( .B(n407), .A(n77), .S(n58), .Y(n1127) );
  MUX2X1 U545 ( .B(n408), .A(n78), .S(n58), .Y(n1126) );
  MUX2X1 U546 ( .B(n409), .A(n79), .S(n58), .Y(n1125) );
  MUX2X1 U547 ( .B(n410), .A(n80), .S(n58), .Y(n1124) );
  MUX2X1 U548 ( .B(n411), .A(n81), .S(n58), .Y(n1123) );
  MUX2X1 U549 ( .B(n412), .A(n82), .S(n58), .Y(n1122) );
  MUX2X1 U550 ( .B(n413), .A(n83), .S(n58), .Y(n1121) );
  MUX2X1 U551 ( .B(n414), .A(n84), .S(n58), .Y(n1120) );
  MUX2X1 U552 ( .B(n415), .A(n77), .S(n59), .Y(n1119) );
  MUX2X1 U553 ( .B(n416), .A(n78), .S(n59), .Y(n1118) );
  MUX2X1 U554 ( .B(n417), .A(n79), .S(n59), .Y(n1117) );
  MUX2X1 U555 ( .B(n418), .A(n80), .S(n59), .Y(n1116) );
  MUX2X1 U556 ( .B(n419), .A(n81), .S(n59), .Y(n1115) );
  MUX2X1 U557 ( .B(n420), .A(n82), .S(n59), .Y(n1114) );
  MUX2X1 U558 ( .B(n421), .A(n83), .S(n59), .Y(n1113) );
  MUX2X1 U559 ( .B(n422), .A(n84), .S(n59), .Y(n1112) );
  MUX2X1 U560 ( .B(n423), .A(n77), .S(n60), .Y(n1111) );
  MUX2X1 U561 ( .B(n424), .A(n78), .S(n60), .Y(n1110) );
  MUX2X1 U562 ( .B(n425), .A(n79), .S(n60), .Y(n1109) );
  MUX2X1 U563 ( .B(n426), .A(n80), .S(n60), .Y(n1108) );
  MUX2X1 U564 ( .B(n427), .A(n81), .S(n60), .Y(n1107) );
  MUX2X1 U565 ( .B(n428), .A(n82), .S(n60), .Y(n1106) );
  MUX2X1 U566 ( .B(n429), .A(n83), .S(n60), .Y(n1105) );
  MUX2X1 U567 ( .B(n430), .A(n84), .S(n60), .Y(n1104) );
  INVX1 U568 ( .A(n431), .Y(n1103) );
  MUX2X1 U569 ( .B(\memory[28][7] ), .A(RCV_DATA[7]), .S(n432), .Y(n431) );
  INVX1 U570 ( .A(n433), .Y(n1102) );
  MUX2X1 U571 ( .B(\memory[28][6] ), .A(RCV_DATA[6]), .S(n432), .Y(n433) );
  INVX1 U572 ( .A(n434), .Y(n1101) );
  MUX2X1 U573 ( .B(\memory[28][5] ), .A(RCV_DATA[5]), .S(n432), .Y(n434) );
  INVX1 U574 ( .A(n435), .Y(n1100) );
  MUX2X1 U575 ( .B(\memory[28][4] ), .A(RCV_DATA[4]), .S(n432), .Y(n435) );
  INVX1 U576 ( .A(n436), .Y(n1099) );
  MUX2X1 U577 ( .B(\memory[28][3] ), .A(RCV_DATA[3]), .S(n432), .Y(n436) );
  INVX1 U578 ( .A(n437), .Y(n1098) );
  MUX2X1 U579 ( .B(\memory[28][2] ), .A(RCV_DATA[2]), .S(n432), .Y(n437) );
  INVX1 U580 ( .A(n438), .Y(n1097) );
  MUX2X1 U581 ( .B(\memory[28][1] ), .A(RCV_DATA[1]), .S(n432), .Y(n438) );
  INVX1 U582 ( .A(n439), .Y(n1096) );
  MUX2X1 U583 ( .B(\memory[28][0] ), .A(RCV_DATA[0]), .S(n432), .Y(n439) );
  INVX1 U584 ( .A(n440), .Y(n1095) );
  MUX2X1 U585 ( .B(\memory[29][7] ), .A(RCV_DATA[7]), .S(n61), .Y(n440) );
  INVX1 U586 ( .A(n441), .Y(n1094) );
  MUX2X1 U587 ( .B(\memory[29][6] ), .A(RCV_DATA[6]), .S(n61), .Y(n441) );
  INVX1 U588 ( .A(n442), .Y(n1093) );
  MUX2X1 U589 ( .B(\memory[29][5] ), .A(RCV_DATA[5]), .S(n61), .Y(n442) );
  INVX1 U590 ( .A(n443), .Y(n1092) );
  MUX2X1 U591 ( .B(\memory[29][4] ), .A(RCV_DATA[4]), .S(n61), .Y(n443) );
  INVX1 U592 ( .A(n444), .Y(n1091) );
  MUX2X1 U593 ( .B(\memory[29][3] ), .A(RCV_DATA[3]), .S(n61), .Y(n444) );
  INVX1 U594 ( .A(n445), .Y(n1090) );
  MUX2X1 U595 ( .B(\memory[29][2] ), .A(RCV_DATA[2]), .S(n61), .Y(n445) );
  INVX1 U596 ( .A(n446), .Y(n1089) );
  MUX2X1 U597 ( .B(\memory[29][1] ), .A(RCV_DATA[1]), .S(n61), .Y(n446) );
  INVX1 U598 ( .A(n447), .Y(n1088) );
  MUX2X1 U599 ( .B(\memory[29][0] ), .A(RCV_DATA[0]), .S(n61), .Y(n447) );
  INVX1 U600 ( .A(n448), .Y(n1087) );
  MUX2X1 U601 ( .B(\memory[30][7] ), .A(RCV_DATA[7]), .S(n62), .Y(n448) );
  INVX1 U602 ( .A(n450), .Y(n1086) );
  MUX2X1 U603 ( .B(\memory[30][6] ), .A(RCV_DATA[6]), .S(n62), .Y(n450) );
  INVX1 U604 ( .A(n451), .Y(n1085) );
  MUX2X1 U605 ( .B(\memory[30][5] ), .A(RCV_DATA[5]), .S(n62), .Y(n451) );
  INVX1 U606 ( .A(n452), .Y(n1084) );
  MUX2X1 U607 ( .B(\memory[30][4] ), .A(RCV_DATA[4]), .S(n62), .Y(n452) );
  INVX1 U608 ( .A(n453), .Y(n1083) );
  MUX2X1 U609 ( .B(\memory[30][3] ), .A(RCV_DATA[3]), .S(n62), .Y(n453) );
  INVX1 U610 ( .A(n454), .Y(n1082) );
  MUX2X1 U611 ( .B(\memory[30][2] ), .A(RCV_DATA[2]), .S(n62), .Y(n454) );
  INVX1 U612 ( .A(n455), .Y(n1081) );
  MUX2X1 U613 ( .B(\memory[30][1] ), .A(RCV_DATA[1]), .S(n62), .Y(n455) );
  INVX1 U614 ( .A(n456), .Y(n1080) );
  MUX2X1 U615 ( .B(\memory[30][0] ), .A(RCV_DATA[0]), .S(n62), .Y(n456) );
  INVX1 U616 ( .A(n457), .Y(n1079) );
  MUX2X1 U617 ( .B(\memory[31][7] ), .A(RCV_DATA[7]), .S(n458), .Y(n457) );
  INVX1 U618 ( .A(n459), .Y(n1078) );
  MUX2X1 U619 ( .B(\memory[31][6] ), .A(RCV_DATA[6]), .S(n458), .Y(n459) );
  INVX1 U620 ( .A(n460), .Y(n1077) );
  MUX2X1 U621 ( .B(\memory[31][5] ), .A(RCV_DATA[5]), .S(n458), .Y(n460) );
  INVX1 U622 ( .A(n461), .Y(n1076) );
  MUX2X1 U623 ( .B(\memory[31][4] ), .A(RCV_DATA[4]), .S(n458), .Y(n461) );
  INVX1 U624 ( .A(n462), .Y(n1075) );
  MUX2X1 U625 ( .B(\memory[31][3] ), .A(RCV_DATA[3]), .S(n458), .Y(n462) );
  INVX1 U626 ( .A(n463), .Y(n1074) );
  MUX2X1 U627 ( .B(\memory[31][2] ), .A(RCV_DATA[2]), .S(n458), .Y(n463) );
  INVX1 U628 ( .A(n464), .Y(n1073) );
  MUX2X1 U629 ( .B(\memory[31][1] ), .A(RCV_DATA[1]), .S(n458), .Y(n464) );
  INVX1 U630 ( .A(n465), .Y(n1072) );
  MUX2X1 U631 ( .B(\memory[31][0] ), .A(RCV_DATA[0]), .S(n458), .Y(n465) );
  MUX2X1 U632 ( .B(n466), .A(n75), .S(n467), .Y(n1063) );
  MUX2X1 U633 ( .B(n468), .A(n76), .S(n467), .Y(n1062) );
  OAI21X1 U634 ( .A(n184), .B(n146), .C(n364), .Y(n467) );
  NAND2X1 U635 ( .A(n244), .B(n120), .Y(n364) );
  MUX2X1 U636 ( .B(n469), .A(n75), .S(n470), .Y(n1061) );
  MUX2X1 U637 ( .B(n471), .A(n76), .S(n470), .Y(n1060) );
  OAI21X1 U638 ( .A(n175), .B(n146), .C(n373), .Y(n470) );
  NAND2X1 U639 ( .A(n244), .B(n115), .Y(n373) );
  MUX2X1 U640 ( .B(n472), .A(n75), .S(n473), .Y(n1059) );
  MUX2X1 U641 ( .B(n474), .A(n76), .S(n473), .Y(n1058) );
  OAI21X1 U642 ( .A(n235), .B(n146), .C(n382), .Y(n473) );
  NAND2X1 U643 ( .A(n244), .B(n110), .Y(n382) );
  NAND2X1 U644 ( .A(n475), .B(n356), .Y(n146) );
  MUX2X1 U645 ( .B(n74), .A(n476), .S(n477), .Y(n1057) );
  MUX2X1 U646 ( .B(n76), .A(n478), .S(n477), .Y(n1056) );
  NAND3X1 U647 ( .A(n475), .B(n353), .C(n479), .Y(n477) );
  MUX2X1 U648 ( .B(n175), .A(n226), .S(n480), .Y(n479) );
  AND2X1 U649 ( .A(n352), .B(n71), .Y(n475) );
  MUX2X1 U650 ( .B(n74), .A(n481), .S(n482), .Y(n1055) );
  MUX2X1 U651 ( .B(n76), .A(n483), .S(n482), .Y(n1054) );
  AOI21X1 U652 ( .A(n110), .B(n126), .C(n57), .Y(n482) );
  INVX1 U653 ( .A(n184), .Y(n110) );
  MUX2X1 U654 ( .B(n74), .A(n484), .S(n485), .Y(n1053) );
  MUX2X1 U655 ( .B(n76), .A(n486), .S(n485), .Y(n1052) );
  AOI21X1 U656 ( .A(n105), .B(n126), .C(n58), .Y(n485) );
  INVX1 U657 ( .A(n175), .Y(n105) );
  MUX2X1 U658 ( .B(n74), .A(n487), .S(n488), .Y(n1051) );
  MUX2X1 U659 ( .B(n76), .A(n489), .S(n488), .Y(n1050) );
  AOI21X1 U660 ( .A(n100), .B(n126), .C(n59), .Y(n488) );
  NAND3X1 U661 ( .A(n358), .B(n64), .C(n67), .Y(n184) );
  INVX1 U662 ( .A(n235), .Y(n100) );
  MUX2X1 U663 ( .B(n74), .A(n490), .S(n491), .Y(n1049) );
  MUX2X1 U664 ( .B(n76), .A(n492), .S(n491), .Y(n1048) );
  AOI21X1 U665 ( .A(n95), .B(n126), .C(n60), .Y(n491) );
  NAND3X1 U666 ( .A(n69), .B(n64), .C(n67), .Y(n175) );
  NAND3X1 U667 ( .A(n493), .B(n70), .C(n356), .Y(n135) );
  INVX1 U668 ( .A(n226), .Y(n95) );
  MUX2X1 U669 ( .B(n74), .A(n494), .S(n495), .Y(n1047) );
  INVX1 U670 ( .A(\opcode[28][1] ), .Y(n494) );
  MUX2X1 U671 ( .B(n76), .A(n496), .S(n495), .Y(n1046) );
  AOI21X1 U672 ( .A(n96), .B(n130), .C(n432), .Y(n495) );
  NAND3X1 U673 ( .A(n358), .B(n360), .C(n65), .Y(n235) );
  INVX1 U674 ( .A(n151), .Y(n130) );
  INVX1 U675 ( .A(\opcode[28][0] ), .Y(n496) );
  MUX2X1 U676 ( .B(n74), .A(n497), .S(n498), .Y(n1045) );
  INVX1 U677 ( .A(\opcode[29][1] ), .Y(n497) );
  MUX2X1 U678 ( .B(n76), .A(n499), .S(n498), .Y(n1044) );
  AOI21X1 U679 ( .A(n96), .B(n125), .C(n61), .Y(n498) );
  NAND3X1 U680 ( .A(n69), .B(n360), .C(n65), .Y(n226) );
  INVX1 U681 ( .A(n145), .Y(n125) );
  NAND3X1 U682 ( .A(n356), .B(n493), .C(n71), .Y(n500) );
  INVX1 U683 ( .A(\opcode[29][0] ), .Y(n499) );
  MUX2X1 U684 ( .B(n74), .A(n501), .S(n502), .Y(n1043) );
  INVX1 U685 ( .A(\opcode[30][1] ), .Y(n501) );
  MUX2X1 U686 ( .B(n76), .A(n503), .S(n502), .Y(n1042) );
  AOI21X1 U687 ( .A(n120), .B(n156), .C(n62), .Y(n502) );
  NOR2X1 U688 ( .A(n151), .B(n174), .Y(n449) );
  NAND3X1 U689 ( .A(n65), .B(n358), .C(n67), .Y(n151) );
  INVX1 U690 ( .A(n140), .Y(n120) );
  NAND3X1 U691 ( .A(n360), .B(n64), .C(n358), .Y(n140) );
  INVX1 U692 ( .A(n69), .Y(n358) );
  INVX1 U693 ( .A(\opcode[30][0] ), .Y(n503) );
  MUX2X1 U694 ( .B(n75), .A(n504), .S(n505), .Y(n1041) );
  INVX1 U695 ( .A(\opcode[31][1] ), .Y(n504) );
  MUX2X1 U696 ( .B(n93), .A(n506), .S(n505), .Y(n1040) );
  AOI21X1 U697 ( .A(n115), .B(n156), .C(n458), .Y(n505) );
  NOR2X1 U698 ( .A(n507), .B(n480), .Y(n351) );
  NOR2X1 U699 ( .A(n354), .B(RST), .Y(n493) );
  INVX1 U700 ( .A(writeptr[4]), .Y(n354) );
  NAND3X1 U701 ( .A(n65), .B(n69), .C(n67), .Y(n145) );
  NAND3X1 U702 ( .A(n356), .B(n70), .C(n352), .Y(n508) );
  NOR2X1 U703 ( .A(writeptr[4]), .B(RST), .Y(n352) );
  NAND2X1 U704 ( .A(W_ENABLE), .B(n302), .Y(n507) );
  NAND3X1 U705 ( .A(n509), .B(n510), .C(n511), .Y(n302) );
  NOR2X1 U706 ( .A(n512), .B(n513), .Y(n511) );
  XOR2X1 U707 ( .A(readptr[3]), .B(N34), .Y(n512) );
  XOR2X1 U708 ( .A(n514), .B(N32), .Y(n510) );
  NOR2X1 U709 ( .A(n515), .B(n516), .Y(n509) );
  XOR2X1 U710 ( .A(readptr[2]), .B(N33), .Y(n515) );
  INVX1 U711 ( .A(n134), .Y(n115) );
  NAND3X1 U712 ( .A(n360), .B(n64), .C(n69), .Y(n134) );
  INVX1 U713 ( .A(n67), .Y(n360) );
  INVX1 U714 ( .A(\opcode[31][0] ), .Y(n506) );
  INVX1 U715 ( .A(n517), .Y(n1039) );
  MUX2X1 U716 ( .B(n518), .A(DATA[7]), .S(n519), .Y(n517) );
  NAND2X1 U717 ( .A(n520), .B(n521), .Y(n518) );
  NOR2X1 U718 ( .A(n522), .B(n523), .Y(n521) );
  NAND3X1 U719 ( .A(n524), .B(n525), .C(n526), .Y(n523) );
  NOR2X1 U720 ( .A(n527), .B(n528), .Y(n526) );
  OAI22X1 U721 ( .A(n399), .B(n529), .C(n407), .D(n530), .Y(n528) );
  INVX1 U722 ( .A(\memory[17][7] ), .Y(n407) );
  INVX1 U723 ( .A(\memory[16][7] ), .Y(n399) );
  OAI22X1 U724 ( .A(n415), .B(n531), .C(n423), .D(n532), .Y(n527) );
  INVX1 U725 ( .A(\memory[19][7] ), .Y(n423) );
  INVX1 U726 ( .A(\memory[18][7] ), .Y(n415) );
  AOI22X1 U727 ( .A(n533), .B(\memory[23][7] ), .C(n534), .D(\memory[22][7] ), 
        .Y(n525) );
  AOI22X1 U728 ( .A(n535), .B(\memory[21][7] ), .C(n536), .D(\memory[20][7] ), 
        .Y(n524) );
  NAND3X1 U729 ( .A(n537), .B(n538), .C(n539), .Y(n522) );
  NOR2X1 U730 ( .A(n540), .B(n541), .Y(n539) );
  OAI22X1 U731 ( .A(n193), .B(n542), .C(n185), .D(n543), .Y(n541) );
  INVX1 U732 ( .A(\memory[25][7] ), .Y(n185) );
  INVX1 U733 ( .A(\memory[24][7] ), .Y(n193) );
  OAI22X1 U734 ( .A(n176), .B(n544), .C(n166), .D(n545), .Y(n540) );
  INVX1 U735 ( .A(\memory[27][7] ), .Y(n166) );
  INVX1 U736 ( .A(\memory[26][7] ), .Y(n176) );
  AOI22X1 U737 ( .A(n546), .B(\memory[31][7] ), .C(n547), .D(\memory[30][7] ), 
        .Y(n538) );
  AOI22X1 U738 ( .A(n548), .B(\memory[29][7] ), .C(n549), .D(\memory[28][7] ), 
        .Y(n537) );
  NOR2X1 U739 ( .A(n550), .B(n551), .Y(n520) );
  NAND3X1 U740 ( .A(n552), .B(n553), .C(n554), .Y(n551) );
  NOR2X1 U741 ( .A(n555), .B(n556), .Y(n554) );
  OAI22X1 U742 ( .A(n301), .B(n557), .C(n293), .D(n558), .Y(n556) );
  INVX1 U743 ( .A(\memory[2][7] ), .Y(n293) );
  INVX1 U744 ( .A(\memory[3][7] ), .Y(n301) );
  OAI22X1 U745 ( .A(n285), .B(n559), .C(n276), .D(n560), .Y(n555) );
  INVX1 U746 ( .A(\memory[0][7] ), .Y(n276) );
  INVX1 U747 ( .A(\memory[1][7] ), .Y(n285) );
  AOI22X1 U748 ( .A(n561), .B(\memory[4][7] ), .C(n562), .D(\memory[5][7] ), 
        .Y(n553) );
  AOI22X1 U749 ( .A(n563), .B(\memory[6][7] ), .C(n564), .D(\memory[7][7] ), 
        .Y(n552) );
  NAND3X1 U750 ( .A(n565), .B(n566), .C(n567), .Y(n550) );
  NOR2X1 U751 ( .A(n568), .B(n569), .Y(n567) );
  OAI22X1 U752 ( .A(n363), .B(n570), .C(n372), .D(n571), .Y(n569) );
  INVX1 U753 ( .A(\memory[9][7] ), .Y(n372) );
  INVX1 U754 ( .A(\memory[8][7] ), .Y(n363) );
  OAI22X1 U755 ( .A(n381), .B(n572), .C(n390), .D(n573), .Y(n568) );
  INVX1 U756 ( .A(\memory[11][7] ), .Y(n390) );
  INVX1 U757 ( .A(\memory[10][7] ), .Y(n381) );
  AOI22X1 U758 ( .A(n574), .B(\memory[15][7] ), .C(n575), .D(\memory[14][7] ), 
        .Y(n566) );
  AOI22X1 U759 ( .A(n576), .B(\memory[13][7] ), .C(n577), .D(\memory[12][7] ), 
        .Y(n565) );
  INVX1 U760 ( .A(n578), .Y(n1038) );
  MUX2X1 U761 ( .B(n579), .A(DATA[6]), .S(n519), .Y(n578) );
  NAND2X1 U762 ( .A(n580), .B(n581), .Y(n579) );
  NOR2X1 U763 ( .A(n582), .B(n583), .Y(n581) );
  NAND3X1 U764 ( .A(n584), .B(n585), .C(n586), .Y(n583) );
  NOR2X1 U765 ( .A(n587), .B(n588), .Y(n586) );
  OAI22X1 U766 ( .A(n400), .B(n529), .C(n408), .D(n530), .Y(n588) );
  INVX1 U767 ( .A(\memory[17][6] ), .Y(n408) );
  INVX1 U768 ( .A(\memory[16][6] ), .Y(n400) );
  OAI22X1 U769 ( .A(n416), .B(n531), .C(n424), .D(n532), .Y(n587) );
  INVX1 U770 ( .A(\memory[19][6] ), .Y(n424) );
  INVX1 U771 ( .A(\memory[18][6] ), .Y(n416) );
  AOI22X1 U772 ( .A(n533), .B(\memory[23][6] ), .C(n534), .D(\memory[22][6] ), 
        .Y(n585) );
  AOI22X1 U773 ( .A(n535), .B(\memory[21][6] ), .C(n536), .D(\memory[20][6] ), 
        .Y(n584) );
  NAND3X1 U774 ( .A(n589), .B(n590), .C(n591), .Y(n582) );
  NOR2X1 U775 ( .A(n592), .B(n593), .Y(n591) );
  OAI22X1 U776 ( .A(n194), .B(n542), .C(n186), .D(n543), .Y(n593) );
  INVX1 U777 ( .A(\memory[25][6] ), .Y(n186) );
  INVX1 U778 ( .A(\memory[24][6] ), .Y(n194) );
  OAI22X1 U779 ( .A(n177), .B(n544), .C(n167), .D(n545), .Y(n592) );
  INVX1 U780 ( .A(\memory[27][6] ), .Y(n167) );
  INVX1 U781 ( .A(\memory[26][6] ), .Y(n177) );
  AOI22X1 U782 ( .A(n546), .B(\memory[31][6] ), .C(n547), .D(\memory[30][6] ), 
        .Y(n590) );
  AOI22X1 U783 ( .A(n548), .B(\memory[29][6] ), .C(n549), .D(\memory[28][6] ), 
        .Y(n589) );
  NOR2X1 U784 ( .A(n594), .B(n595), .Y(n580) );
  NAND3X1 U785 ( .A(n596), .B(n597), .C(n598), .Y(n595) );
  NOR2X1 U786 ( .A(n599), .B(n600), .Y(n598) );
  OAI22X1 U787 ( .A(n300), .B(n557), .C(n292), .D(n558), .Y(n600) );
  INVX1 U788 ( .A(\memory[2][6] ), .Y(n292) );
  INVX1 U789 ( .A(\memory[3][6] ), .Y(n300) );
  OAI22X1 U790 ( .A(n284), .B(n559), .C(n275), .D(n560), .Y(n599) );
  INVX1 U791 ( .A(\memory[0][6] ), .Y(n275) );
  INVX1 U792 ( .A(\memory[1][6] ), .Y(n284) );
  AOI22X1 U793 ( .A(n561), .B(\memory[4][6] ), .C(n562), .D(\memory[5][6] ), 
        .Y(n597) );
  AOI22X1 U794 ( .A(n563), .B(\memory[6][6] ), .C(n564), .D(\memory[7][6] ), 
        .Y(n596) );
  NAND3X1 U795 ( .A(n601), .B(n602), .C(n603), .Y(n594) );
  NOR2X1 U796 ( .A(n604), .B(n605), .Y(n603) );
  OAI22X1 U797 ( .A(n365), .B(n570), .C(n374), .D(n571), .Y(n605) );
  INVX1 U798 ( .A(\memory[9][6] ), .Y(n374) );
  INVX1 U799 ( .A(\memory[8][6] ), .Y(n365) );
  OAI22X1 U800 ( .A(n383), .B(n572), .C(n392), .D(n573), .Y(n604) );
  INVX1 U801 ( .A(\memory[11][6] ), .Y(n392) );
  INVX1 U802 ( .A(\memory[10][6] ), .Y(n383) );
  AOI22X1 U803 ( .A(n574), .B(\memory[15][6] ), .C(n575), .D(\memory[14][6] ), 
        .Y(n602) );
  AOI22X1 U804 ( .A(n576), .B(\memory[13][6] ), .C(n577), .D(\memory[12][6] ), 
        .Y(n601) );
  INVX1 U805 ( .A(n606), .Y(n1037) );
  MUX2X1 U806 ( .B(n607), .A(DATA[5]), .S(n519), .Y(n606) );
  NAND2X1 U807 ( .A(n608), .B(n609), .Y(n607) );
  NOR2X1 U808 ( .A(n610), .B(n611), .Y(n609) );
  NAND3X1 U809 ( .A(n612), .B(n613), .C(n614), .Y(n611) );
  NOR2X1 U810 ( .A(n615), .B(n616), .Y(n614) );
  OAI22X1 U811 ( .A(n401), .B(n529), .C(n409), .D(n530), .Y(n616) );
  INVX1 U812 ( .A(\memory[17][5] ), .Y(n409) );
  INVX1 U813 ( .A(\memory[16][5] ), .Y(n401) );
  OAI22X1 U814 ( .A(n417), .B(n531), .C(n425), .D(n532), .Y(n615) );
  INVX1 U815 ( .A(\memory[19][5] ), .Y(n425) );
  INVX1 U816 ( .A(\memory[18][5] ), .Y(n417) );
  AOI22X1 U817 ( .A(n533), .B(\memory[23][5] ), .C(n534), .D(\memory[22][5] ), 
        .Y(n613) );
  AOI22X1 U818 ( .A(n535), .B(\memory[21][5] ), .C(n536), .D(\memory[20][5] ), 
        .Y(n612) );
  NAND3X1 U819 ( .A(n617), .B(n618), .C(n619), .Y(n610) );
  NOR2X1 U820 ( .A(n620), .B(n621), .Y(n619) );
  OAI22X1 U821 ( .A(n195), .B(n542), .C(n187), .D(n543), .Y(n621) );
  INVX1 U822 ( .A(\memory[25][5] ), .Y(n187) );
  INVX1 U823 ( .A(\memory[24][5] ), .Y(n195) );
  OAI22X1 U824 ( .A(n178), .B(n544), .C(n168), .D(n545), .Y(n620) );
  INVX1 U825 ( .A(\memory[27][5] ), .Y(n168) );
  INVX1 U826 ( .A(\memory[26][5] ), .Y(n178) );
  AOI22X1 U827 ( .A(n546), .B(\memory[31][5] ), .C(n547), .D(\memory[30][5] ), 
        .Y(n618) );
  AOI22X1 U828 ( .A(n548), .B(\memory[29][5] ), .C(n549), .D(\memory[28][5] ), 
        .Y(n617) );
  NOR2X1 U829 ( .A(n622), .B(n623), .Y(n608) );
  NAND3X1 U830 ( .A(n624), .B(n625), .C(n626), .Y(n623) );
  NOR2X1 U831 ( .A(n627), .B(n628), .Y(n626) );
  OAI22X1 U832 ( .A(n299), .B(n557), .C(n291), .D(n558), .Y(n628) );
  INVX1 U833 ( .A(\memory[2][5] ), .Y(n291) );
  INVX1 U834 ( .A(\memory[3][5] ), .Y(n299) );
  OAI22X1 U835 ( .A(n283), .B(n559), .C(n274), .D(n560), .Y(n627) );
  INVX1 U836 ( .A(\memory[0][5] ), .Y(n274) );
  INVX1 U837 ( .A(\memory[1][5] ), .Y(n283) );
  AOI22X1 U838 ( .A(n561), .B(\memory[4][5] ), .C(n562), .D(\memory[5][5] ), 
        .Y(n625) );
  AOI22X1 U839 ( .A(n563), .B(\memory[6][5] ), .C(n564), .D(\memory[7][5] ), 
        .Y(n624) );
  NAND3X1 U840 ( .A(n629), .B(n630), .C(n631), .Y(n622) );
  NOR2X1 U841 ( .A(n632), .B(n633), .Y(n631) );
  OAI22X1 U842 ( .A(n366), .B(n570), .C(n375), .D(n571), .Y(n633) );
  INVX1 U843 ( .A(\memory[9][5] ), .Y(n375) );
  INVX1 U844 ( .A(\memory[8][5] ), .Y(n366) );
  OAI22X1 U845 ( .A(n384), .B(n572), .C(n393), .D(n573), .Y(n632) );
  INVX1 U846 ( .A(\memory[11][5] ), .Y(n393) );
  INVX1 U847 ( .A(\memory[10][5] ), .Y(n384) );
  AOI22X1 U848 ( .A(n574), .B(\memory[15][5] ), .C(n575), .D(\memory[14][5] ), 
        .Y(n630) );
  AOI22X1 U849 ( .A(n576), .B(\memory[13][5] ), .C(n577), .D(\memory[12][5] ), 
        .Y(n629) );
  INVX1 U850 ( .A(n634), .Y(n1036) );
  MUX2X1 U851 ( .B(n635), .A(DATA[4]), .S(n519), .Y(n634) );
  NAND2X1 U852 ( .A(n636), .B(n637), .Y(n635) );
  NOR2X1 U853 ( .A(n638), .B(n639), .Y(n637) );
  NAND3X1 U854 ( .A(n640), .B(n641), .C(n642), .Y(n639) );
  NOR2X1 U855 ( .A(n643), .B(n644), .Y(n642) );
  OAI22X1 U856 ( .A(n402), .B(n529), .C(n410), .D(n530), .Y(n644) );
  INVX1 U857 ( .A(\memory[17][4] ), .Y(n410) );
  INVX1 U858 ( .A(\memory[16][4] ), .Y(n402) );
  OAI22X1 U859 ( .A(n418), .B(n531), .C(n426), .D(n532), .Y(n643) );
  INVX1 U860 ( .A(\memory[19][4] ), .Y(n426) );
  INVX1 U861 ( .A(\memory[18][4] ), .Y(n418) );
  AOI22X1 U862 ( .A(n533), .B(\memory[23][4] ), .C(n534), .D(\memory[22][4] ), 
        .Y(n641) );
  AOI22X1 U863 ( .A(n535), .B(\memory[21][4] ), .C(n536), .D(\memory[20][4] ), 
        .Y(n640) );
  NAND3X1 U864 ( .A(n645), .B(n646), .C(n647), .Y(n638) );
  NOR2X1 U865 ( .A(n648), .B(n649), .Y(n647) );
  OAI22X1 U866 ( .A(n196), .B(n542), .C(n188), .D(n543), .Y(n649) );
  INVX1 U867 ( .A(\memory[25][4] ), .Y(n188) );
  INVX1 U868 ( .A(\memory[24][4] ), .Y(n196) );
  OAI22X1 U869 ( .A(n179), .B(n544), .C(n169), .D(n545), .Y(n648) );
  INVX1 U870 ( .A(\memory[27][4] ), .Y(n169) );
  INVX1 U871 ( .A(\memory[26][4] ), .Y(n179) );
  AOI22X1 U872 ( .A(n546), .B(\memory[31][4] ), .C(n547), .D(\memory[30][4] ), 
        .Y(n646) );
  AOI22X1 U873 ( .A(n548), .B(\memory[29][4] ), .C(n549), .D(\memory[28][4] ), 
        .Y(n645) );
  NOR2X1 U874 ( .A(n650), .B(n651), .Y(n636) );
  NAND3X1 U875 ( .A(n652), .B(n653), .C(n654), .Y(n651) );
  NOR2X1 U876 ( .A(n655), .B(n656), .Y(n654) );
  OAI22X1 U877 ( .A(n298), .B(n557), .C(n290), .D(n558), .Y(n656) );
  INVX1 U878 ( .A(\memory[2][4] ), .Y(n290) );
  INVX1 U879 ( .A(\memory[3][4] ), .Y(n298) );
  OAI22X1 U880 ( .A(n282), .B(n559), .C(n273), .D(n560), .Y(n655) );
  INVX1 U881 ( .A(\memory[0][4] ), .Y(n273) );
  INVX1 U882 ( .A(\memory[1][4] ), .Y(n282) );
  AOI22X1 U883 ( .A(n561), .B(\memory[4][4] ), .C(n562), .D(\memory[5][4] ), 
        .Y(n653) );
  AOI22X1 U884 ( .A(n563), .B(\memory[6][4] ), .C(n564), .D(\memory[7][4] ), 
        .Y(n652) );
  NAND3X1 U885 ( .A(n657), .B(n658), .C(n659), .Y(n650) );
  NOR2X1 U886 ( .A(n660), .B(n661), .Y(n659) );
  OAI22X1 U887 ( .A(n367), .B(n570), .C(n376), .D(n571), .Y(n661) );
  INVX1 U888 ( .A(\memory[9][4] ), .Y(n376) );
  INVX1 U889 ( .A(\memory[8][4] ), .Y(n367) );
  OAI22X1 U890 ( .A(n385), .B(n572), .C(n394), .D(n573), .Y(n660) );
  INVX1 U891 ( .A(\memory[11][4] ), .Y(n394) );
  INVX1 U892 ( .A(\memory[10][4] ), .Y(n385) );
  AOI22X1 U893 ( .A(n574), .B(\memory[15][4] ), .C(n575), .D(\memory[14][4] ), 
        .Y(n658) );
  AOI22X1 U894 ( .A(n576), .B(\memory[13][4] ), .C(n577), .D(\memory[12][4] ), 
        .Y(n657) );
  INVX1 U895 ( .A(n662), .Y(n1035) );
  MUX2X1 U896 ( .B(n663), .A(DATA[3]), .S(n519), .Y(n662) );
  NAND2X1 U897 ( .A(n664), .B(n665), .Y(n663) );
  NOR2X1 U898 ( .A(n666), .B(n667), .Y(n665) );
  NAND3X1 U899 ( .A(n668), .B(n669), .C(n670), .Y(n667) );
  NOR2X1 U900 ( .A(n671), .B(n672), .Y(n670) );
  OAI22X1 U901 ( .A(n403), .B(n529), .C(n411), .D(n530), .Y(n672) );
  INVX1 U902 ( .A(\memory[17][3] ), .Y(n411) );
  INVX1 U903 ( .A(\memory[16][3] ), .Y(n403) );
  OAI22X1 U904 ( .A(n419), .B(n531), .C(n427), .D(n532), .Y(n671) );
  INVX1 U905 ( .A(\memory[19][3] ), .Y(n427) );
  INVX1 U906 ( .A(\memory[18][3] ), .Y(n419) );
  AOI22X1 U907 ( .A(n533), .B(\memory[23][3] ), .C(n534), .D(\memory[22][3] ), 
        .Y(n669) );
  AOI22X1 U908 ( .A(n535), .B(\memory[21][3] ), .C(n536), .D(\memory[20][3] ), 
        .Y(n668) );
  NAND3X1 U909 ( .A(n673), .B(n674), .C(n675), .Y(n666) );
  NOR2X1 U910 ( .A(n676), .B(n677), .Y(n675) );
  OAI22X1 U911 ( .A(n197), .B(n542), .C(n189), .D(n543), .Y(n677) );
  INVX1 U912 ( .A(\memory[25][3] ), .Y(n189) );
  INVX1 U913 ( .A(\memory[24][3] ), .Y(n197) );
  OAI22X1 U914 ( .A(n180), .B(n544), .C(n170), .D(n545), .Y(n676) );
  INVX1 U915 ( .A(\memory[27][3] ), .Y(n170) );
  INVX1 U916 ( .A(\memory[26][3] ), .Y(n180) );
  AOI22X1 U917 ( .A(n546), .B(\memory[31][3] ), .C(n547), .D(\memory[30][3] ), 
        .Y(n674) );
  AOI22X1 U918 ( .A(n548), .B(\memory[29][3] ), .C(n549), .D(\memory[28][3] ), 
        .Y(n673) );
  NOR2X1 U919 ( .A(n678), .B(n679), .Y(n664) );
  NAND3X1 U920 ( .A(n680), .B(n681), .C(n682), .Y(n679) );
  NOR2X1 U921 ( .A(n683), .B(n684), .Y(n682) );
  OAI22X1 U922 ( .A(n297), .B(n557), .C(n289), .D(n558), .Y(n684) );
  INVX1 U923 ( .A(\memory[2][3] ), .Y(n289) );
  INVX1 U924 ( .A(\memory[3][3] ), .Y(n297) );
  OAI22X1 U925 ( .A(n281), .B(n559), .C(n272), .D(n560), .Y(n683) );
  INVX1 U926 ( .A(\memory[0][3] ), .Y(n272) );
  INVX1 U927 ( .A(\memory[1][3] ), .Y(n281) );
  AOI22X1 U928 ( .A(n561), .B(\memory[4][3] ), .C(n562), .D(\memory[5][3] ), 
        .Y(n681) );
  AOI22X1 U929 ( .A(n563), .B(\memory[6][3] ), .C(n564), .D(\memory[7][3] ), 
        .Y(n680) );
  NAND3X1 U930 ( .A(n685), .B(n686), .C(n687), .Y(n678) );
  NOR2X1 U931 ( .A(n688), .B(n689), .Y(n687) );
  OAI22X1 U932 ( .A(n368), .B(n570), .C(n377), .D(n571), .Y(n689) );
  INVX1 U933 ( .A(\memory[9][3] ), .Y(n377) );
  INVX1 U934 ( .A(\memory[8][3] ), .Y(n368) );
  OAI22X1 U935 ( .A(n386), .B(n572), .C(n395), .D(n573), .Y(n688) );
  INVX1 U936 ( .A(\memory[11][3] ), .Y(n395) );
  INVX1 U937 ( .A(\memory[10][3] ), .Y(n386) );
  AOI22X1 U938 ( .A(n574), .B(\memory[15][3] ), .C(n575), .D(\memory[14][3] ), 
        .Y(n686) );
  AOI22X1 U939 ( .A(n576), .B(\memory[13][3] ), .C(n577), .D(\memory[12][3] ), 
        .Y(n685) );
  INVX1 U940 ( .A(n690), .Y(n1034) );
  MUX2X1 U941 ( .B(n691), .A(DATA[2]), .S(n519), .Y(n690) );
  NAND2X1 U942 ( .A(n692), .B(n693), .Y(n691) );
  NOR2X1 U943 ( .A(n694), .B(n695), .Y(n693) );
  NAND3X1 U944 ( .A(n696), .B(n697), .C(n698), .Y(n695) );
  NOR2X1 U945 ( .A(n699), .B(n700), .Y(n698) );
  OAI22X1 U946 ( .A(n404), .B(n529), .C(n412), .D(n530), .Y(n700) );
  INVX1 U947 ( .A(\memory[17][2] ), .Y(n412) );
  INVX1 U948 ( .A(\memory[16][2] ), .Y(n404) );
  OAI22X1 U949 ( .A(n420), .B(n531), .C(n428), .D(n532), .Y(n699) );
  INVX1 U950 ( .A(\memory[19][2] ), .Y(n428) );
  INVX1 U951 ( .A(\memory[18][2] ), .Y(n420) );
  AOI22X1 U952 ( .A(n533), .B(\memory[23][2] ), .C(n534), .D(\memory[22][2] ), 
        .Y(n697) );
  AOI22X1 U953 ( .A(n535), .B(\memory[21][2] ), .C(n536), .D(\memory[20][2] ), 
        .Y(n696) );
  NAND3X1 U954 ( .A(n701), .B(n702), .C(n703), .Y(n694) );
  NOR2X1 U955 ( .A(n704), .B(n705), .Y(n703) );
  OAI22X1 U956 ( .A(n198), .B(n542), .C(n190), .D(n543), .Y(n705) );
  INVX1 U957 ( .A(\memory[25][2] ), .Y(n190) );
  INVX1 U958 ( .A(\memory[24][2] ), .Y(n198) );
  OAI22X1 U959 ( .A(n181), .B(n544), .C(n171), .D(n545), .Y(n704) );
  INVX1 U960 ( .A(\memory[27][2] ), .Y(n171) );
  INVX1 U961 ( .A(\memory[26][2] ), .Y(n181) );
  AOI22X1 U962 ( .A(n546), .B(\memory[31][2] ), .C(n547), .D(\memory[30][2] ), 
        .Y(n702) );
  AOI22X1 U963 ( .A(n548), .B(\memory[29][2] ), .C(n549), .D(\memory[28][2] ), 
        .Y(n701) );
  NOR2X1 U964 ( .A(n706), .B(n707), .Y(n692) );
  NAND3X1 U965 ( .A(n708), .B(n709), .C(n710), .Y(n707) );
  NOR2X1 U966 ( .A(n711), .B(n712), .Y(n710) );
  OAI22X1 U967 ( .A(n296), .B(n557), .C(n288), .D(n558), .Y(n712) );
  INVX1 U968 ( .A(\memory[2][2] ), .Y(n288) );
  INVX1 U969 ( .A(\memory[3][2] ), .Y(n296) );
  OAI22X1 U970 ( .A(n280), .B(n559), .C(n271), .D(n560), .Y(n711) );
  INVX1 U971 ( .A(\memory[0][2] ), .Y(n271) );
  INVX1 U972 ( .A(\memory[1][2] ), .Y(n280) );
  AOI22X1 U973 ( .A(n561), .B(\memory[4][2] ), .C(n562), .D(\memory[5][2] ), 
        .Y(n709) );
  AOI22X1 U974 ( .A(n563), .B(\memory[6][2] ), .C(n564), .D(\memory[7][2] ), 
        .Y(n708) );
  NAND3X1 U975 ( .A(n713), .B(n714), .C(n715), .Y(n706) );
  NOR2X1 U976 ( .A(n716), .B(n717), .Y(n715) );
  OAI22X1 U977 ( .A(n369), .B(n570), .C(n378), .D(n571), .Y(n717) );
  INVX1 U978 ( .A(\memory[9][2] ), .Y(n378) );
  INVX1 U979 ( .A(\memory[8][2] ), .Y(n369) );
  OAI22X1 U980 ( .A(n387), .B(n572), .C(n396), .D(n573), .Y(n716) );
  INVX1 U981 ( .A(\memory[11][2] ), .Y(n396) );
  INVX1 U982 ( .A(\memory[10][2] ), .Y(n387) );
  AOI22X1 U983 ( .A(n574), .B(\memory[15][2] ), .C(n575), .D(\memory[14][2] ), 
        .Y(n714) );
  AOI22X1 U984 ( .A(n576), .B(\memory[13][2] ), .C(n577), .D(\memory[12][2] ), 
        .Y(n713) );
  INVX1 U985 ( .A(n718), .Y(n1033) );
  MUX2X1 U986 ( .B(n719), .A(DATA[1]), .S(n519), .Y(n718) );
  NAND2X1 U987 ( .A(n720), .B(n721), .Y(n719) );
  NOR2X1 U988 ( .A(n722), .B(n723), .Y(n721) );
  NAND3X1 U989 ( .A(n724), .B(n725), .C(n726), .Y(n723) );
  NOR2X1 U990 ( .A(n727), .B(n728), .Y(n726) );
  OAI22X1 U991 ( .A(n405), .B(n529), .C(n413), .D(n530), .Y(n728) );
  INVX1 U992 ( .A(\memory[17][1] ), .Y(n413) );
  INVX1 U993 ( .A(\memory[16][1] ), .Y(n405) );
  OAI22X1 U994 ( .A(n421), .B(n531), .C(n429), .D(n532), .Y(n727) );
  INVX1 U995 ( .A(\memory[19][1] ), .Y(n429) );
  INVX1 U996 ( .A(\memory[18][1] ), .Y(n421) );
  AOI22X1 U997 ( .A(n533), .B(\memory[23][1] ), .C(n534), .D(\memory[22][1] ), 
        .Y(n725) );
  AOI22X1 U998 ( .A(n535), .B(\memory[21][1] ), .C(n536), .D(\memory[20][1] ), 
        .Y(n724) );
  NAND3X1 U999 ( .A(n729), .B(n730), .C(n731), .Y(n722) );
  NOR2X1 U1000 ( .A(n732), .B(n733), .Y(n731) );
  OAI22X1 U1001 ( .A(n199), .B(n542), .C(n191), .D(n543), .Y(n733) );
  INVX1 U1002 ( .A(\memory[25][1] ), .Y(n191) );
  INVX1 U1003 ( .A(\memory[24][1] ), .Y(n199) );
  OAI22X1 U1004 ( .A(n182), .B(n544), .C(n172), .D(n545), .Y(n732) );
  INVX1 U1005 ( .A(\memory[27][1] ), .Y(n172) );
  INVX1 U1006 ( .A(\memory[26][1] ), .Y(n182) );
  AOI22X1 U1007 ( .A(n546), .B(\memory[31][1] ), .C(n547), .D(\memory[30][1] ), 
        .Y(n730) );
  AOI22X1 U1008 ( .A(n548), .B(\memory[29][1] ), .C(n549), .D(\memory[28][1] ), 
        .Y(n729) );
  NOR2X1 U1009 ( .A(n734), .B(n735), .Y(n720) );
  NAND3X1 U1010 ( .A(n736), .B(n737), .C(n738), .Y(n735) );
  NOR2X1 U1011 ( .A(n739), .B(n740), .Y(n738) );
  OAI22X1 U1012 ( .A(n295), .B(n557), .C(n287), .D(n558), .Y(n740) );
  INVX1 U1013 ( .A(\memory[2][1] ), .Y(n287) );
  INVX1 U1014 ( .A(\memory[3][1] ), .Y(n295) );
  OAI22X1 U1015 ( .A(n279), .B(n559), .C(n270), .D(n560), .Y(n739) );
  INVX1 U1016 ( .A(\memory[0][1] ), .Y(n270) );
  INVX1 U1017 ( .A(\memory[1][1] ), .Y(n279) );
  AOI22X1 U1018 ( .A(n561), .B(\memory[4][1] ), .C(n562), .D(\memory[5][1] ), 
        .Y(n737) );
  AOI22X1 U1019 ( .A(n563), .B(\memory[6][1] ), .C(n564), .D(\memory[7][1] ), 
        .Y(n736) );
  NAND3X1 U1020 ( .A(n741), .B(n742), .C(n743), .Y(n734) );
  NOR2X1 U1021 ( .A(n744), .B(n745), .Y(n743) );
  OAI22X1 U1022 ( .A(n370), .B(n570), .C(n379), .D(n571), .Y(n745) );
  INVX1 U1023 ( .A(\memory[9][1] ), .Y(n379) );
  INVX1 U1024 ( .A(\memory[8][1] ), .Y(n370) );
  OAI22X1 U1025 ( .A(n388), .B(n572), .C(n397), .D(n573), .Y(n744) );
  INVX1 U1026 ( .A(\memory[11][1] ), .Y(n397) );
  INVX1 U1027 ( .A(\memory[10][1] ), .Y(n388) );
  AOI22X1 U1028 ( .A(n574), .B(\memory[15][1] ), .C(n575), .D(\memory[14][1] ), 
        .Y(n742) );
  AOI22X1 U1029 ( .A(n576), .B(\memory[13][1] ), .C(n577), .D(\memory[12][1] ), 
        .Y(n741) );
  INVX1 U1030 ( .A(n746), .Y(n1032) );
  MUX2X1 U1031 ( .B(n747), .A(DATA[0]), .S(n519), .Y(n746) );
  NAND2X1 U1032 ( .A(n748), .B(n749), .Y(n747) );
  NOR2X1 U1033 ( .A(n750), .B(n751), .Y(n749) );
  NAND3X1 U1034 ( .A(n752), .B(n753), .C(n754), .Y(n751) );
  NOR2X1 U1035 ( .A(n755), .B(n756), .Y(n754) );
  OAI22X1 U1036 ( .A(n406), .B(n529), .C(n414), .D(n530), .Y(n756) );
  INVX1 U1037 ( .A(\memory[17][0] ), .Y(n414) );
  INVX1 U1038 ( .A(\memory[16][0] ), .Y(n406) );
  OAI22X1 U1039 ( .A(n422), .B(n531), .C(n430), .D(n532), .Y(n755) );
  INVX1 U1040 ( .A(\memory[19][0] ), .Y(n430) );
  INVX1 U1041 ( .A(\memory[18][0] ), .Y(n422) );
  AOI22X1 U1042 ( .A(n533), .B(\memory[23][0] ), .C(n534), .D(\memory[22][0] ), 
        .Y(n753) );
  AOI22X1 U1043 ( .A(n535), .B(\memory[21][0] ), .C(n536), .D(\memory[20][0] ), 
        .Y(n752) );
  NAND3X1 U1044 ( .A(n757), .B(n758), .C(n759), .Y(n750) );
  NOR2X1 U1045 ( .A(n760), .B(n761), .Y(n759) );
  OAI22X1 U1046 ( .A(n200), .B(n542), .C(n192), .D(n543), .Y(n761) );
  INVX1 U1047 ( .A(\memory[25][0] ), .Y(n192) );
  INVX1 U1048 ( .A(\memory[24][0] ), .Y(n200) );
  OAI22X1 U1049 ( .A(n183), .B(n544), .C(n173), .D(n545), .Y(n760) );
  INVX1 U1050 ( .A(\memory[27][0] ), .Y(n173) );
  INVX1 U1051 ( .A(\memory[26][0] ), .Y(n183) );
  AOI22X1 U1052 ( .A(n546), .B(\memory[31][0] ), .C(n547), .D(\memory[30][0] ), 
        .Y(n758) );
  AOI22X1 U1053 ( .A(n548), .B(\memory[29][0] ), .C(n549), .D(\memory[28][0] ), 
        .Y(n757) );
  NOR2X1 U1054 ( .A(n762), .B(n763), .Y(n748) );
  NAND3X1 U1055 ( .A(n764), .B(n765), .C(n766), .Y(n763) );
  NOR2X1 U1056 ( .A(n767), .B(n768), .Y(n766) );
  OAI22X1 U1057 ( .A(n294), .B(n557), .C(n286), .D(n558), .Y(n768) );
  INVX1 U1058 ( .A(\memory[2][0] ), .Y(n286) );
  INVX1 U1059 ( .A(\memory[3][0] ), .Y(n294) );
  OAI22X1 U1060 ( .A(n278), .B(n559), .C(n269), .D(n560), .Y(n767) );
  INVX1 U1061 ( .A(\memory[0][0] ), .Y(n269) );
  INVX1 U1062 ( .A(\memory[1][0] ), .Y(n278) );
  AOI22X1 U1063 ( .A(n561), .B(\memory[4][0] ), .C(n562), .D(\memory[5][0] ), 
        .Y(n765) );
  AOI22X1 U1064 ( .A(n563), .B(\memory[6][0] ), .C(n564), .D(\memory[7][0] ), 
        .Y(n764) );
  NAND3X1 U1065 ( .A(n769), .B(n770), .C(n771), .Y(n762) );
  NOR2X1 U1066 ( .A(n772), .B(n773), .Y(n771) );
  OAI22X1 U1067 ( .A(n371), .B(n570), .C(n380), .D(n571), .Y(n773) );
  INVX1 U1068 ( .A(\memory[9][0] ), .Y(n380) );
  INVX1 U1069 ( .A(\memory[8][0] ), .Y(n371) );
  OAI22X1 U1070 ( .A(n389), .B(n572), .C(n398), .D(n573), .Y(n772) );
  INVX1 U1071 ( .A(\memory[11][0] ), .Y(n398) );
  INVX1 U1072 ( .A(\memory[10][0] ), .Y(n389) );
  AOI22X1 U1073 ( .A(n574), .B(\memory[15][0] ), .C(n575), .D(\memory[14][0] ), 
        .Y(n770) );
  AOI22X1 U1074 ( .A(n576), .B(\memory[13][0] ), .C(n577), .D(\memory[12][0] ), 
        .Y(n769) );
  INVX1 U1075 ( .A(n774), .Y(n1031) );
  MUX2X1 U1076 ( .B(n775), .A(OUT_OPCODE[1]), .S(n519), .Y(n774) );
  NAND2X1 U1077 ( .A(n776), .B(n777), .Y(n775) );
  NOR2X1 U1078 ( .A(n778), .B(n779), .Y(n777) );
  NAND3X1 U1079 ( .A(n780), .B(n781), .C(n782), .Y(n779) );
  NOR2X1 U1080 ( .A(n783), .B(n784), .Y(n782) );
  OAI22X1 U1081 ( .A(n481), .B(n529), .C(n484), .D(n530), .Y(n784) );
  INVX1 U1082 ( .A(\opcode[17][1] ), .Y(n484) );
  INVX1 U1083 ( .A(\opcode[16][1] ), .Y(n481) );
  OAI22X1 U1084 ( .A(n487), .B(n531), .C(n490), .D(n532), .Y(n783) );
  INVX1 U1085 ( .A(\opcode[19][1] ), .Y(n490) );
  INVX1 U1086 ( .A(\opcode[18][1] ), .Y(n487) );
  AOI22X1 U1087 ( .A(n533), .B(\opcode[23][1] ), .C(n534), .D(\opcode[22][1] ), 
        .Y(n781) );
  AOI22X1 U1088 ( .A(n535), .B(\opcode[21][1] ), .C(n536), .D(\opcode[20][1] ), 
        .Y(n780) );
  NAND3X1 U1089 ( .A(n785), .B(n786), .C(n787), .Y(n778) );
  NOR2X1 U1090 ( .A(n788), .B(n789), .Y(n787) );
  OAI22X1 U1091 ( .A(n107), .B(n542), .C(n102), .D(n543), .Y(n789) );
  INVX1 U1092 ( .A(\opcode[25][1] ), .Y(n102) );
  INVX1 U1093 ( .A(\opcode[24][1] ), .Y(n107) );
  OAI22X1 U1094 ( .A(n97), .B(n544), .C(n91), .D(n545), .Y(n788) );
  INVX1 U1095 ( .A(\opcode[27][1] ), .Y(n91) );
  INVX1 U1096 ( .A(\opcode[26][1] ), .Y(n97) );
  AOI22X1 U1097 ( .A(n546), .B(\opcode[31][1] ), .C(n547), .D(\opcode[30][1] ), 
        .Y(n786) );
  AOI22X1 U1098 ( .A(n548), .B(\opcode[29][1] ), .C(n549), .D(\opcode[28][1] ), 
        .Y(n785) );
  NOR2X1 U1099 ( .A(n790), .B(n791), .Y(n776) );
  NAND3X1 U1100 ( .A(n792), .B(n793), .C(n794), .Y(n791) );
  NOR2X1 U1101 ( .A(n795), .B(n796), .Y(n794) );
  OAI22X1 U1102 ( .A(n165), .B(n557), .C(n162), .D(n558), .Y(n796) );
  INVX1 U1103 ( .A(\opcode[2][1] ), .Y(n162) );
  INVX1 U1104 ( .A(\opcode[3][1] ), .Y(n165) );
  OAI22X1 U1105 ( .A(n159), .B(n559), .C(n155), .D(n560), .Y(n795) );
  INVX1 U1106 ( .A(\opcode[0][1] ), .Y(n155) );
  INVX1 U1107 ( .A(\opcode[1][1] ), .Y(n159) );
  AOI22X1 U1108 ( .A(n561), .B(\opcode[4][1] ), .C(n562), .D(\opcode[5][1] ), 
        .Y(n793) );
  AOI22X1 U1109 ( .A(n563), .B(\opcode[6][1] ), .C(n564), .D(\opcode[7][1] ), 
        .Y(n792) );
  NAND3X1 U1110 ( .A(n797), .B(n798), .C(n799), .Y(n790) );
  NOR2X1 U1111 ( .A(n800), .B(n801), .Y(n799) );
  OAI22X1 U1112 ( .A(n466), .B(n570), .C(n469), .D(n571), .Y(n801) );
  INVX1 U1113 ( .A(\opcode[9][1] ), .Y(n469) );
  INVX1 U1114 ( .A(\opcode[8][1] ), .Y(n466) );
  OAI22X1 U1115 ( .A(n472), .B(n572), .C(n476), .D(n573), .Y(n800) );
  INVX1 U1116 ( .A(\opcode[11][1] ), .Y(n476) );
  INVX1 U1117 ( .A(\opcode[10][1] ), .Y(n472) );
  AOI22X1 U1118 ( .A(n574), .B(\opcode[15][1] ), .C(n575), .D(\opcode[14][1] ), 
        .Y(n798) );
  AOI22X1 U1119 ( .A(n576), .B(\opcode[13][1] ), .C(n577), .D(\opcode[12][1] ), 
        .Y(n797) );
  INVX1 U1120 ( .A(n802), .Y(n1030) );
  MUX2X1 U1121 ( .B(n803), .A(OUT_OPCODE[0]), .S(n519), .Y(n802) );
  NAND3X1 U1122 ( .A(N195), .B(n85), .C(n72), .Y(n519) );
  NAND2X1 U1123 ( .A(n804), .B(n805), .Y(n803) );
  NOR2X1 U1124 ( .A(n806), .B(n807), .Y(n805) );
  NAND3X1 U1125 ( .A(n808), .B(n809), .C(n810), .Y(n807) );
  NOR2X1 U1126 ( .A(n811), .B(n812), .Y(n810) );
  OAI22X1 U1127 ( .A(n483), .B(n529), .C(n486), .D(n530), .Y(n812) );
  NAND2X1 U1128 ( .A(n813), .B(n814), .Y(n530) );
  INVX1 U1129 ( .A(\opcode[17][0] ), .Y(n486) );
  NAND2X1 U1130 ( .A(n815), .B(n814), .Y(n529) );
  INVX1 U1131 ( .A(\opcode[16][0] ), .Y(n483) );
  OAI22X1 U1132 ( .A(n489), .B(n531), .C(n492), .D(n532), .Y(n811) );
  NAND2X1 U1133 ( .A(n813), .B(n816), .Y(n532) );
  INVX1 U1134 ( .A(\opcode[19][0] ), .Y(n492) );
  NAND2X1 U1135 ( .A(n815), .B(n816), .Y(n531) );
  INVX1 U1136 ( .A(\opcode[18][0] ), .Y(n489) );
  AOI22X1 U1137 ( .A(n533), .B(\opcode[23][0] ), .C(n534), .D(\opcode[22][0] ), 
        .Y(n809) );
  AOI22X1 U1138 ( .A(n535), .B(\opcode[21][0] ), .C(n536), .D(\opcode[20][0] ), 
        .Y(n808) );
  INVX1 U1139 ( .A(n819), .Y(n815) );
  NAND3X1 U1140 ( .A(n820), .B(n821), .C(readptr[4]), .Y(n819) );
  INVX1 U1141 ( .A(n822), .Y(n813) );
  NAND3X1 U1142 ( .A(readptr[0]), .B(n821), .C(readptr[4]), .Y(n822) );
  NAND3X1 U1143 ( .A(n823), .B(n824), .C(n825), .Y(n806) );
  NOR2X1 U1144 ( .A(n826), .B(n827), .Y(n825) );
  OAI22X1 U1145 ( .A(n109), .B(n542), .C(n104), .D(n543), .Y(n827) );
  NAND2X1 U1146 ( .A(n814), .B(n828), .Y(n543) );
  INVX1 U1147 ( .A(\opcode[25][0] ), .Y(n104) );
  NAND2X1 U1148 ( .A(n814), .B(n829), .Y(n542) );
  INVX1 U1149 ( .A(\opcode[24][0] ), .Y(n109) );
  OAI22X1 U1150 ( .A(n99), .B(n544), .C(n94), .D(n545), .Y(n826) );
  NAND2X1 U1151 ( .A(n816), .B(n828), .Y(n545) );
  INVX1 U1152 ( .A(\opcode[27][0] ), .Y(n94) );
  NAND2X1 U1153 ( .A(n816), .B(n829), .Y(n544) );
  INVX1 U1154 ( .A(\opcode[26][0] ), .Y(n99) );
  AOI22X1 U1155 ( .A(n546), .B(\opcode[31][0] ), .C(n547), .D(\opcode[30][0] ), 
        .Y(n824) );
  AOI22X1 U1156 ( .A(n548), .B(\opcode[29][0] ), .C(n549), .D(\opcode[28][0] ), 
        .Y(n823) );
  INVX1 U1157 ( .A(n830), .Y(n829) );
  NAND3X1 U1158 ( .A(readptr[3]), .B(n820), .C(readptr[4]), .Y(n830) );
  INVX1 U1159 ( .A(n831), .Y(n828) );
  NAND3X1 U1160 ( .A(readptr[3]), .B(readptr[0]), .C(readptr[4]), .Y(n831) );
  NOR2X1 U1161 ( .A(n832), .B(n833), .Y(n804) );
  NAND3X1 U1162 ( .A(n834), .B(n835), .C(n836), .Y(n833) );
  NOR2X1 U1163 ( .A(n837), .B(n838), .Y(n836) );
  OAI22X1 U1164 ( .A(n163), .B(n557), .C(n160), .D(n558), .Y(n838) );
  NAND2X1 U1165 ( .A(n839), .B(n816), .Y(n558) );
  INVX1 U1166 ( .A(\opcode[2][0] ), .Y(n160) );
  NAND2X1 U1167 ( .A(n840), .B(n816), .Y(n557) );
  INVX1 U1168 ( .A(\opcode[3][0] ), .Y(n163) );
  OAI22X1 U1169 ( .A(n157), .B(n559), .C(n153), .D(n560), .Y(n837) );
  NAND2X1 U1170 ( .A(n839), .B(n814), .Y(n560) );
  INVX1 U1171 ( .A(\opcode[0][0] ), .Y(n153) );
  NAND2X1 U1172 ( .A(n840), .B(n814), .Y(n559) );
  INVX1 U1173 ( .A(\opcode[1][0] ), .Y(n157) );
  AOI22X1 U1174 ( .A(n561), .B(\opcode[4][0] ), .C(n562), .D(\opcode[5][0] ), 
        .Y(n835) );
  AOI22X1 U1175 ( .A(n563), .B(\opcode[6][0] ), .C(n564), .D(\opcode[7][0] ), 
        .Y(n834) );
  INVX1 U1176 ( .A(n841), .Y(n840) );
  NAND3X1 U1177 ( .A(n821), .B(n842), .C(readptr[0]), .Y(n841) );
  INVX1 U1178 ( .A(n843), .Y(n839) );
  NAND3X1 U1179 ( .A(n821), .B(n842), .C(n820), .Y(n843) );
  INVX1 U1180 ( .A(readptr[3]), .Y(n821) );
  NAND3X1 U1181 ( .A(n844), .B(n845), .C(n846), .Y(n832) );
  NOR2X1 U1182 ( .A(n847), .B(n848), .Y(n846) );
  OAI22X1 U1183 ( .A(n468), .B(n570), .C(n471), .D(n571), .Y(n848) );
  NAND2X1 U1184 ( .A(n849), .B(n814), .Y(n571) );
  INVX1 U1185 ( .A(\opcode[9][0] ), .Y(n471) );
  NAND2X1 U1186 ( .A(n850), .B(n814), .Y(n570) );
  NOR2X1 U1187 ( .A(readptr[1]), .B(readptr[2]), .Y(n814) );
  INVX1 U1188 ( .A(\opcode[8][0] ), .Y(n468) );
  OAI22X1 U1189 ( .A(n474), .B(n572), .C(n478), .D(n573), .Y(n847) );
  NAND2X1 U1190 ( .A(n849), .B(n816), .Y(n573) );
  INVX1 U1191 ( .A(\opcode[11][0] ), .Y(n478) );
  NAND2X1 U1192 ( .A(n850), .B(n816), .Y(n572) );
  NOR2X1 U1193 ( .A(n514), .B(readptr[2]), .Y(n816) );
  INVX1 U1194 ( .A(\opcode[10][0] ), .Y(n474) );
  AOI22X1 U1195 ( .A(n574), .B(\opcode[15][0] ), .C(n575), .D(\opcode[14][0] ), 
        .Y(n845) );
  NOR2X1 U1196 ( .A(n514), .B(n851), .Y(n817) );
  AOI22X1 U1197 ( .A(n576), .B(\opcode[13][0] ), .C(n577), .D(\opcode[12][0] ), 
        .Y(n844) );
  INVX1 U1198 ( .A(n852), .Y(n850) );
  NAND3X1 U1199 ( .A(n820), .B(n842), .C(readptr[3]), .Y(n852) );
  INVX1 U1200 ( .A(readptr[0]), .Y(n820) );
  NOR2X1 U1201 ( .A(n851), .B(readptr[1]), .Y(n818) );
  INVX1 U1202 ( .A(readptr[2]), .Y(n851) );
  INVX1 U1203 ( .A(n853), .Y(n849) );
  NAND3X1 U1204 ( .A(readptr[0]), .B(n842), .C(readptr[3]), .Y(n853) );
  INVX1 U1205 ( .A(readptr[4]), .Y(n842) );
  AND2X1 U1207 ( .A(N337), .B(n72), .Y(N347) );
  AND2X1 U1208 ( .A(N336), .B(n72), .Y(N346) );
  AND2X1 U1209 ( .A(N335), .B(n72), .Y(N345) );
  AND2X1 U1210 ( .A(N334), .B(n72), .Y(N344) );
  AND2X1 U1211 ( .A(N333), .B(n72), .Y(N343) );
  AND2X1 U1212 ( .A(N193), .B(n72), .Y(N342) );
  AND2X1 U1213 ( .A(N192), .B(n72), .Y(N341) );
  AND2X1 U1214 ( .A(N191), .B(n72), .Y(N340) );
  AND2X1 U1215 ( .A(N190), .B(n72), .Y(N339) );
  AND2X1 U1216 ( .A(N189), .B(n72), .Y(N338) );
  AND2X1 U1217 ( .A(R_ENABLE), .B(n304), .Y(N195) );
  NAND3X1 U1218 ( .A(n855), .B(n857), .C(n859), .Y(n304) );
  NOR2X1 U1219 ( .A(n861), .B(n863), .Y(n859) );
  XOR2X1 U1220 ( .A(writeptr[4]), .B(readptr[4]), .Y(n863) );
  XOR2X1 U1221 ( .A(n71), .B(readptr[3]), .Y(n861) );
  XOR2X1 U1222 ( .A(n514), .B(n67), .Y(n857) );
  INVX1 U1223 ( .A(readptr[1]), .Y(n514) );
  NOR2X1 U1224 ( .A(n864), .B(n865), .Y(n855) );
  XOR2X1 U1225 ( .A(n69), .B(readptr[0]), .Y(n865) );
  XOR2X1 U1226 ( .A(n65), .B(readptr[2]), .Y(n864) );
endmodule


module memoryblock_1 ( CLK, NEXT_BYTE, RCV_DATA, RCV_OPCODE, RST, W_ENABLE, 
        EOP, EMPTY, FULL, B_READY, PRGA_IN, PRGA_OPCODE );
  input [7:0] RCV_DATA;
  input [1:0] RCV_OPCODE;
  output [7:0] PRGA_IN;
  output [1:0] PRGA_OPCODE;
  input CLK, NEXT_BYTE, RST, W_ENABLE, EOP;
  output EMPTY, FULL, B_READY;
  wire   R_ENABLE;
  wire   [4:0] BYTE_COUNT;
  wire   [7:0] DATA;
  wire   [1:0] OUT_OPCODE;

  RBUFFER_1 U_0 ( .CLK(CLK), .RST(RST), .NEXT_BYTE(NEXT_BYTE), .DATA(DATA), 
        .OPCODE(OUT_OPCODE), .BYTE_COUNT(BYTE_COUNT), .EOP(EOP), .B_READY(
        B_READY), .R_ENABLE(R_ENABLE), .PRGA_IN(PRGA_IN), .PRGA_OPCODE(
        PRGA_OPCODE) );
  RFIFO_1 U_1 ( .CLK(CLK), .RST(RST), .W_ENABLE(W_ENABLE), .R_ENABLE(R_ENABLE), 
        .RCV_DATA(RCV_DATA), .RCV_OPCODE(RCV_OPCODE), .DATA(DATA), 
        .OUT_OPCODE(OUT_OPCODE), .BYTE_COUNT(BYTE_COUNT), .EMPTY(EMPTY), 
        .FULL(FULL) );
endmodule


module rx_CRC_CALC_1 ( CLK, RST, W_ENABLE, OPCODE, RCV_DATA, RX_CRC );
  input [1:0] OPCODE;
  input [7:0] RCV_DATA;
  output [15:0] RX_CRC;
  input CLK, RST, W_ENABLE;
  wire   n3, n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31,
         n33, n51, n52, n53, n54, n55, n57, n58, n59, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n101, n103, n105, n107, n109, n111, n113, n115, n117, n119,
         n121, n123, n125, n127, n129, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n32, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n56, n60, n79, n80, n81, n82, n100, n102, n104, n106, n108,
         n110, n112, n114, n116, n118, n120, n122, n124, n126, n128, n130,
         n131, n148, n149, n150, n151, n152, n153, n154, n155, n156;
  wire   [15:0] current_crc;
  wire   [15:0] cache_1;

  DFFPOSX1 \cache_1_reg[0]  ( .D(n129), .CLK(CLK), .Q(cache_1[0]) );
  DFFPOSX1 \cache_1_reg[8]  ( .D(n127), .CLK(CLK), .Q(cache_1[8]) );
  DFFPOSX1 \cache_1_reg[15]  ( .D(n125), .CLK(CLK), .Q(cache_1[15]) );
  DFFPOSX1 \cache_1_reg[1]  ( .D(n123), .CLK(CLK), .Q(cache_1[1]) );
  DFFPOSX1 \cache_1_reg[9]  ( .D(n121), .CLK(CLK), .Q(cache_1[9]) );
  DFFPOSX1 \cache_1_reg[2]  ( .D(n119), .CLK(CLK), .Q(cache_1[2]) );
  DFFPOSX1 \cache_1_reg[10]  ( .D(n117), .CLK(CLK), .Q(cache_1[10]) );
  DFFPOSX1 \cache_1_reg[3]  ( .D(n115), .CLK(CLK), .Q(cache_1[3]) );
  DFFPOSX1 \cache_1_reg[11]  ( .D(n113), .CLK(CLK), .Q(cache_1[11]) );
  DFFPOSX1 \cache_1_reg[4]  ( .D(n111), .CLK(CLK), .Q(cache_1[4]) );
  DFFPOSX1 \cache_1_reg[12]  ( .D(n109), .CLK(CLK), .Q(cache_1[12]) );
  DFFPOSX1 \cache_1_reg[5]  ( .D(n107), .CLK(CLK), .Q(cache_1[5]) );
  DFFPOSX1 \cache_1_reg[13]  ( .D(n105), .CLK(CLK), .Q(cache_1[13]) );
  DFFPOSX1 \cache_1_reg[6]  ( .D(n103), .CLK(CLK), .Q(cache_1[6]) );
  DFFPOSX1 \cache_1_reg[14]  ( .D(n101), .CLK(CLK), .Q(cache_1[14]) );
  DFFPOSX1 \cache_1_reg[7]  ( .D(n99), .CLK(CLK), .Q(cache_1[7]) );
  DFFPOSX1 \cache_2_reg[15]  ( .D(n98), .CLK(CLK), .Q(RX_CRC[15]) );
  DFFPOSX1 \cache_2_reg[14]  ( .D(n97), .CLK(CLK), .Q(RX_CRC[14]) );
  DFFPOSX1 \cache_2_reg[13]  ( .D(n96), .CLK(CLK), .Q(RX_CRC[13]) );
  DFFPOSX1 \cache_2_reg[12]  ( .D(n95), .CLK(CLK), .Q(RX_CRC[12]) );
  DFFPOSX1 \cache_2_reg[11]  ( .D(n94), .CLK(CLK), .Q(RX_CRC[11]) );
  DFFPOSX1 \cache_2_reg[10]  ( .D(n93), .CLK(CLK), .Q(RX_CRC[10]) );
  DFFPOSX1 \cache_2_reg[9]  ( .D(n92), .CLK(CLK), .Q(RX_CRC[9]) );
  DFFPOSX1 \cache_2_reg[8]  ( .D(n91), .CLK(CLK), .Q(RX_CRC[8]) );
  DFFPOSX1 \cache_2_reg[7]  ( .D(n90), .CLK(CLK), .Q(RX_CRC[7]) );
  DFFPOSX1 \cache_2_reg[6]  ( .D(n89), .CLK(CLK), .Q(RX_CRC[6]) );
  DFFPOSX1 \cache_2_reg[5]  ( .D(n88), .CLK(CLK), .Q(RX_CRC[5]) );
  DFFPOSX1 \cache_2_reg[4]  ( .D(n87), .CLK(CLK), .Q(RX_CRC[4]) );
  DFFPOSX1 \cache_2_reg[3]  ( .D(n86), .CLK(CLK), .Q(RX_CRC[3]) );
  DFFPOSX1 \cache_2_reg[2]  ( .D(n85), .CLK(CLK), .Q(RX_CRC[2]) );
  DFFPOSX1 \cache_2_reg[1]  ( .D(n84), .CLK(CLK), .Q(RX_CRC[1]) );
  DFFPOSX1 \cache_2_reg[0]  ( .D(n83), .CLK(CLK), .Q(RX_CRC[0]) );
  OAI21X1 U3 ( .A(n42), .B(n60), .C(n3), .Y(n83) );
  NAND2X1 U4 ( .A(RX_CRC[0]), .B(n43), .Y(n3) );
  OAI21X1 U5 ( .A(n41), .B(n102), .C(n5), .Y(n84) );
  NAND2X1 U6 ( .A(RX_CRC[1]), .B(n43), .Y(n5) );
  OAI21X1 U7 ( .A(n41), .B(n110), .C(n7), .Y(n85) );
  NAND2X1 U8 ( .A(RX_CRC[2]), .B(n43), .Y(n7) );
  OAI21X1 U9 ( .A(n41), .B(n118), .C(n9), .Y(n86) );
  NAND2X1 U10 ( .A(RX_CRC[3]), .B(n43), .Y(n9) );
  OAI21X1 U11 ( .A(n41), .B(n126), .C(n11), .Y(n87) );
  NAND2X1 U12 ( .A(RX_CRC[4]), .B(n43), .Y(n11) );
  OAI21X1 U13 ( .A(n41), .B(n148), .C(n13), .Y(n88) );
  NAND2X1 U14 ( .A(RX_CRC[5]), .B(n42), .Y(n13) );
  OAI21X1 U15 ( .A(n41), .B(n152), .C(n15), .Y(n89) );
  NAND2X1 U16 ( .A(RX_CRC[6]), .B(n42), .Y(n15) );
  OAI21X1 U17 ( .A(n41), .B(n156), .C(n17), .Y(n90) );
  NAND2X1 U18 ( .A(RX_CRC[7]), .B(n42), .Y(n17) );
  OAI21X1 U19 ( .A(n41), .B(n80), .C(n19), .Y(n91) );
  NAND2X1 U20 ( .A(RX_CRC[8]), .B(n42), .Y(n19) );
  OAI21X1 U21 ( .A(n41), .B(n106), .C(n21), .Y(n92) );
  NAND2X1 U22 ( .A(RX_CRC[9]), .B(n42), .Y(n21) );
  OAI21X1 U23 ( .A(n42), .B(n114), .C(n23), .Y(n93) );
  NAND2X1 U24 ( .A(RX_CRC[10]), .B(n42), .Y(n23) );
  OAI21X1 U25 ( .A(n42), .B(n122), .C(n25), .Y(n94) );
  NAND2X1 U26 ( .A(RX_CRC[11]), .B(n42), .Y(n25) );
  OAI21X1 U27 ( .A(n42), .B(n130), .C(n27), .Y(n95) );
  NAND2X1 U28 ( .A(RX_CRC[12]), .B(n42), .Y(n27) );
  OAI21X1 U29 ( .A(n42), .B(n150), .C(n29), .Y(n96) );
  NAND2X1 U30 ( .A(RX_CRC[13]), .B(n43), .Y(n29) );
  OAI21X1 U31 ( .A(n42), .B(n154), .C(n31), .Y(n97) );
  NAND2X1 U32 ( .A(RX_CRC[14]), .B(n43), .Y(n31) );
  OAI21X1 U33 ( .A(n42), .B(n82), .C(n33), .Y(n98) );
  NAND2X1 U34 ( .A(RX_CRC[15]), .B(n43), .Y(n33) );
  OAI22X1 U35 ( .A(n41), .B(n155), .C(n39), .D(n156), .Y(n99) );
  OAI22X1 U37 ( .A(n41), .B(n153), .C(n39), .D(n154), .Y(n101) );
  OAI22X1 U39 ( .A(n41), .B(n151), .C(n39), .D(n152), .Y(n103) );
  OAI22X1 U41 ( .A(n41), .B(n149), .C(n39), .D(n150), .Y(n105) );
  OAI22X1 U43 ( .A(n40), .B(n131), .C(n39), .D(n148), .Y(n107) );
  OAI22X1 U45 ( .A(n40), .B(n128), .C(n39), .D(n130), .Y(n109) );
  OAI22X1 U47 ( .A(n40), .B(n124), .C(n39), .D(n126), .Y(n111) );
  OAI22X1 U49 ( .A(n40), .B(n120), .C(n39), .D(n122), .Y(n113) );
  OAI22X1 U51 ( .A(n40), .B(n116), .C(n39), .D(n118), .Y(n115) );
  OAI22X1 U53 ( .A(n40), .B(n112), .C(n38), .D(n114), .Y(n117) );
  OAI22X1 U55 ( .A(n40), .B(n108), .C(n38), .D(n110), .Y(n119) );
  OAI22X1 U57 ( .A(n40), .B(n104), .C(n38), .D(n106), .Y(n121) );
  OAI22X1 U59 ( .A(n40), .B(n100), .C(n38), .D(n102), .Y(n123) );
  OAI22X1 U61 ( .A(n40), .B(n81), .C(n38), .D(n82), .Y(n125) );
  OAI22X1 U63 ( .A(n40), .B(n79), .C(n38), .D(n80), .Y(n127) );
  OAI22X1 U65 ( .A(n40), .B(n56), .C(n38), .D(n60), .Y(n129) );
  OAI22X1 U70 ( .A(n81), .B(n37), .C(n53), .D(n35), .Y(n132) );
  XOR2X1 U71 ( .A(n54), .B(current_crc[7]), .Y(n53) );
  OAI22X1 U72 ( .A(n35), .B(n151), .C(n153), .D(n37), .Y(n133) );
  OAI22X1 U73 ( .A(n35), .B(n131), .C(n149), .D(n52), .Y(n134) );
  OAI22X1 U74 ( .A(n51), .B(n124), .C(n128), .D(n37), .Y(n135) );
  OAI22X1 U75 ( .A(n35), .B(n116), .C(n120), .D(n52), .Y(n136) );
  OAI22X1 U77 ( .A(n51), .B(n108), .C(n112), .D(n37), .Y(n137) );
  OAI22X1 U78 ( .A(n104), .B(n37), .C(n55), .D(n51), .Y(n138) );
  XOR2X1 U79 ( .A(n100), .B(n45), .Y(n55) );
  OAI22X1 U80 ( .A(n79), .B(n52), .C(n57), .D(n35), .Y(n139) );
  XOR2X1 U81 ( .A(n58), .B(n59), .Y(n57) );
  XOR2X1 U82 ( .A(n56), .B(n45), .Y(n58) );
  OAI22X1 U84 ( .A(n155), .B(n37), .C(n46), .D(n51), .Y(n140) );
  OAI22X1 U86 ( .A(n151), .B(n52), .C(n61), .D(n35), .Y(n141) );
  XOR2X1 U87 ( .A(n62), .B(n63), .Y(n61) );
  OAI22X1 U89 ( .A(n131), .B(n37), .C(n64), .D(n51), .Y(n142) );
  OAI22X1 U91 ( .A(n124), .B(n52), .C(n65), .D(n35), .Y(n143) );
  XOR2X1 U92 ( .A(n66), .B(n67), .Y(n65) );
  OAI22X1 U94 ( .A(n116), .B(n37), .C(n68), .D(n51), .Y(n144) );
  OAI22X1 U96 ( .A(n108), .B(n52), .C(n69), .D(n35), .Y(n145) );
  XOR2X1 U97 ( .A(n70), .B(n71), .Y(n69) );
  OAI22X1 U99 ( .A(n100), .B(n37), .C(n72), .D(n51), .Y(n146) );
  XOR2X1 U100 ( .A(n73), .B(n74), .Y(n72) );
  XOR2X1 U101 ( .A(n75), .B(n76), .Y(n73) );
  OAI22X1 U103 ( .A(n56), .B(n52), .C(n54), .D(n35), .Y(n147) );
  XOR2X1 U104 ( .A(n77), .B(n78), .Y(n54) );
  XOR2X1 U105 ( .A(n45), .B(n71), .Y(n78) );
  XOR2X1 U106 ( .A(current_crc[8]), .B(RCV_DATA[0]), .Y(n71) );
  XOR2X1 U108 ( .A(n81), .B(RCV_DATA[7]), .Y(n75) );
  XOR2X1 U110 ( .A(n46), .B(n76), .Y(n77) );
  XOR2X1 U111 ( .A(n68), .B(n64), .Y(n76) );
  XNOR2X1 U112 ( .A(n63), .B(n67), .Y(n64) );
  XOR2X1 U113 ( .A(current_crc[11]), .B(RCV_DATA[3]), .Y(n67) );
  XNOR2X1 U114 ( .A(n128), .B(RCV_DATA[4]), .Y(n63) );
  XOR2X1 U116 ( .A(n70), .B(n48), .Y(n68) );
  XOR2X1 U118 ( .A(n112), .B(RCV_DATA[2]), .Y(n66) );
  XOR2X1 U120 ( .A(n104), .B(RCV_DATA[1]), .Y(n70) );
  XOR2X1 U123 ( .A(n59), .B(n47), .Y(n74) );
  XOR2X1 U125 ( .A(n149), .B(RCV_DATA[5]), .Y(n62) );
  XNOR2X1 U127 ( .A(n153), .B(RCV_DATA[6]), .Y(n59) );
  OAI21X1 U129 ( .A(n50), .B(n49), .C(n51), .Y(n52) );
  NAND3X1 U130 ( .A(OPCODE[0]), .B(n49), .C(W_ENABLE), .Y(n51) );
  DFFSR \current_crc_reg[14]  ( .D(n133), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[14]) );
  DFFSR \current_crc_reg[12]  ( .D(n135), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[12]) );
  DFFSR \current_crc_reg[10]  ( .D(n137), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[10]) );
  DFFSR \current_crc_reg[13]  ( .D(n134), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[13]) );
  DFFSR \current_crc_reg[11]  ( .D(n136), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[11]) );
  DFFSR \current_crc_reg[15]  ( .D(n132), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[15]) );
  DFFSR \current_crc_reg[8]  ( .D(n139), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[8]) );
  DFFSR \current_crc_reg[6]  ( .D(n141), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[6]) );
  DFFSR \current_crc_reg[4]  ( .D(n143), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[4]) );
  DFFSR \current_crc_reg[2]  ( .D(n145), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[2]) );
  DFFSR \current_crc_reg[0]  ( .D(n147), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[0]) );
  DFFSR \current_crc_reg[9]  ( .D(n138), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[9]) );
  DFFSR \current_crc_reg[7]  ( .D(n140), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[7]) );
  DFFSR \current_crc_reg[5]  ( .D(n142), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[5]) );
  DFFSR \current_crc_reg[3]  ( .D(n144), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[3]) );
  DFFSR \current_crc_reg[1]  ( .D(n146), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[1]) );
  INVX2 U36 ( .A(OPCODE[1]), .Y(n49) );
  INVX2 U38 ( .A(n32), .Y(n38) );
  INVX2 U69 ( .A(n51), .Y(n34) );
  BUFX2 U76 ( .A(n32), .Y(n40) );
  BUFX2 U83 ( .A(n32), .Y(n43) );
  INVX2 U85 ( .A(n32), .Y(n39) );
  OR2X2 U88 ( .A(n35), .B(RST), .Y(n32) );
  INVX2 U90 ( .A(n34), .Y(n35) );
  INVX2 U93 ( .A(n36), .Y(n37) );
  INVX2 U95 ( .A(n52), .Y(n36) );
  INVX2 U98 ( .A(RST), .Y(n44) );
  INVX1 U102 ( .A(OPCODE[0]), .Y(n50) );
  BUFX4 U107 ( .A(n32), .Y(n41) );
  BUFX4 U109 ( .A(n32), .Y(n42) );
  INVX2 U115 ( .A(n75), .Y(n45) );
  INVX2 U117 ( .A(n74), .Y(n46) );
  INVX2 U119 ( .A(n62), .Y(n47) );
  INVX2 U121 ( .A(n66), .Y(n48) );
  INVX2 U122 ( .A(current_crc[0]), .Y(n56) );
  INVX2 U124 ( .A(cache_1[0]), .Y(n60) );
  INVX2 U126 ( .A(current_crc[8]), .Y(n79) );
  INVX2 U128 ( .A(cache_1[8]), .Y(n80) );
  INVX2 U131 ( .A(current_crc[15]), .Y(n81) );
  INVX2 U132 ( .A(cache_1[15]), .Y(n82) );
  INVX2 U133 ( .A(current_crc[1]), .Y(n100) );
  INVX2 U134 ( .A(cache_1[1]), .Y(n102) );
  INVX2 U135 ( .A(current_crc[9]), .Y(n104) );
  INVX2 U136 ( .A(cache_1[9]), .Y(n106) );
  INVX2 U137 ( .A(current_crc[2]), .Y(n108) );
  INVX2 U138 ( .A(cache_1[2]), .Y(n110) );
  INVX2 U139 ( .A(current_crc[10]), .Y(n112) );
  INVX2 U140 ( .A(cache_1[10]), .Y(n114) );
  INVX2 U141 ( .A(current_crc[3]), .Y(n116) );
  INVX2 U142 ( .A(cache_1[3]), .Y(n118) );
  INVX2 U143 ( .A(current_crc[11]), .Y(n120) );
  INVX2 U144 ( .A(cache_1[11]), .Y(n122) );
  INVX2 U145 ( .A(current_crc[4]), .Y(n124) );
  INVX2 U146 ( .A(cache_1[4]), .Y(n126) );
  INVX2 U147 ( .A(current_crc[12]), .Y(n128) );
  INVX2 U148 ( .A(cache_1[12]), .Y(n130) );
  INVX2 U149 ( .A(current_crc[5]), .Y(n131) );
  INVX2 U150 ( .A(cache_1[5]), .Y(n148) );
  INVX2 U151 ( .A(current_crc[13]), .Y(n149) );
  INVX2 U152 ( .A(cache_1[13]), .Y(n150) );
  INVX2 U153 ( .A(current_crc[6]), .Y(n151) );
  INVX2 U154 ( .A(cache_1[6]), .Y(n152) );
  INVX2 U155 ( .A(current_crc[14]), .Y(n153) );
  INVX2 U156 ( .A(cache_1[14]), .Y(n154) );
  INVX2 U157 ( .A(current_crc[7]), .Y(n155) );
  INVX2 U158 ( .A(cache_1[7]), .Y(n156) );
endmodule


module rx_accumulator_1 ( CLK, RST, RCV_DATA, W_ENABLE, rx_CHECK_CRC );
  input [7:0] RCV_DATA;
  output [15:0] rx_CHECK_CRC;
  input CLK, RST, W_ENABLE;
  wire   n3, n4, n6, n7, n9, n10, n12, n13, n15, n16, n18, n19, n21, n22, n24,
         n25, n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51,
         n53, n55, n58, n40, n42, n44, n46, n48, n50, n52, n54, n56, n57, n59;

  OAI21X1 U2 ( .A(n40), .B(n59), .C(n3), .Y(n27) );
  NAND2X1 U3 ( .A(rx_CHECK_CRC[8]), .B(n40), .Y(n3) );
  OAI21X1 U4 ( .A(n42), .B(n59), .C(n4), .Y(n29) );
  NAND2X1 U5 ( .A(RCV_DATA[0]), .B(n42), .Y(n4) );
  OAI21X1 U7 ( .A(n40), .B(n57), .C(n6), .Y(n31) );
  NAND2X1 U8 ( .A(rx_CHECK_CRC[9]), .B(n40), .Y(n6) );
  OAI21X1 U9 ( .A(n42), .B(n57), .C(n7), .Y(n33) );
  NAND2X1 U10 ( .A(RCV_DATA[1]), .B(n42), .Y(n7) );
  OAI21X1 U12 ( .A(n40), .B(n56), .C(n9), .Y(n35) );
  NAND2X1 U13 ( .A(rx_CHECK_CRC[10]), .B(n40), .Y(n9) );
  OAI21X1 U14 ( .A(n42), .B(n56), .C(n10), .Y(n37) );
  NAND2X1 U15 ( .A(RCV_DATA[2]), .B(n42), .Y(n10) );
  OAI21X1 U17 ( .A(n40), .B(n54), .C(n12), .Y(n39) );
  NAND2X1 U18 ( .A(rx_CHECK_CRC[11]), .B(n40), .Y(n12) );
  OAI21X1 U19 ( .A(n42), .B(n54), .C(n13), .Y(n41) );
  NAND2X1 U20 ( .A(RCV_DATA[3]), .B(n42), .Y(n13) );
  OAI21X1 U22 ( .A(n40), .B(n52), .C(n15), .Y(n43) );
  NAND2X1 U23 ( .A(rx_CHECK_CRC[12]), .B(n40), .Y(n15) );
  OAI21X1 U24 ( .A(n42), .B(n52), .C(n16), .Y(n45) );
  NAND2X1 U25 ( .A(RCV_DATA[4]), .B(n42), .Y(n16) );
  OAI21X1 U27 ( .A(n40), .B(n50), .C(n18), .Y(n47) );
  NAND2X1 U28 ( .A(rx_CHECK_CRC[13]), .B(n40), .Y(n18) );
  OAI21X1 U29 ( .A(n42), .B(n50), .C(n19), .Y(n49) );
  NAND2X1 U30 ( .A(RCV_DATA[5]), .B(n42), .Y(n19) );
  OAI21X1 U32 ( .A(n40), .B(n48), .C(n21), .Y(n51) );
  NAND2X1 U33 ( .A(rx_CHECK_CRC[14]), .B(n40), .Y(n21) );
  OAI21X1 U34 ( .A(n42), .B(n48), .C(n22), .Y(n53) );
  NAND2X1 U35 ( .A(RCV_DATA[6]), .B(n42), .Y(n22) );
  OAI21X1 U37 ( .A(n40), .B(n46), .C(n24), .Y(n55) );
  NAND2X1 U38 ( .A(rx_CHECK_CRC[15]), .B(n40), .Y(n24) );
  OAI21X1 U41 ( .A(n42), .B(n46), .C(n25), .Y(n58) );
  NAND2X1 U42 ( .A(RCV_DATA[7]), .B(n42), .Y(n25) );
  DFFSR \present_CHECK_CRC_reg[7]  ( .D(n58), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[7]) );
  DFFSR \present_CHECK_CRC_reg[6]  ( .D(n53), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[6]) );
  DFFSR \present_CHECK_CRC_reg[5]  ( .D(n49), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[5]) );
  DFFSR \present_CHECK_CRC_reg[4]  ( .D(n45), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[4]) );
  DFFSR \present_CHECK_CRC_reg[3]  ( .D(n41), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[3]) );
  DFFSR \present_CHECK_CRC_reg[2]  ( .D(n37), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[2]) );
  DFFSR \present_CHECK_CRC_reg[1]  ( .D(n33), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[1]) );
  DFFSR \present_CHECK_CRC_reg[0]  ( .D(n29), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[0]) );
  DFFSR \present_CHECK_CRC_reg[15]  ( .D(n55), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[15]) );
  DFFSR \present_CHECK_CRC_reg[14]  ( .D(n51), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[14]) );
  DFFSR \present_CHECK_CRC_reg[13]  ( .D(n47), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[13]) );
  DFFSR \present_CHECK_CRC_reg[12]  ( .D(n43), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[12]) );
  DFFSR \present_CHECK_CRC_reg[11]  ( .D(n39), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[11]) );
  DFFSR \present_CHECK_CRC_reg[10]  ( .D(n35), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[10]) );
  DFFSR \present_CHECK_CRC_reg[9]  ( .D(n31), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[9]) );
  DFFSR \present_CHECK_CRC_reg[8]  ( .D(n27), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[8]) );
  INVX2 U6 ( .A(W_ENABLE), .Y(n40) );
  INVX2 U51 ( .A(n40), .Y(n42) );
  INVX2 U52 ( .A(RST), .Y(n44) );
  INVX2 U53 ( .A(rx_CHECK_CRC[7]), .Y(n46) );
  INVX2 U54 ( .A(rx_CHECK_CRC[6]), .Y(n48) );
  INVX2 U55 ( .A(rx_CHECK_CRC[5]), .Y(n50) );
  INVX2 U56 ( .A(rx_CHECK_CRC[4]), .Y(n52) );
  INVX2 U57 ( .A(rx_CHECK_CRC[3]), .Y(n54) );
  INVX2 U58 ( .A(rx_CHECK_CRC[2]), .Y(n56) );
  INVX2 U59 ( .A(rx_CHECK_CRC[1]), .Y(n57) );
  INVX2 U60 ( .A(rx_CHECK_CRC[0]), .Y(n59) );
endmodule


module rx_decode_1 ( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP, D_ORIG, BITSTUFF, 
        BS_ERROR );
  input CLK, RST, DP1_RX, SHIFT_ENABLE, EOP;
  output D_ORIG, BITSTUFF, BS_ERROR;
  wire   DP_hold1, DP_hold2, N29, N30, N31, N32, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n6, n8, n9, n10, n12, n13,
         n14, n15, n16;
  wire   [3:0] state;

  DFFSR DP_hold2_reg ( .D(n44), .CLK(CLK), .R(1'b1), .S(n6), .Q(DP_hold2) );
  DFFSR DP_hold1_reg ( .D(n43), .CLK(CLK), .R(1'b1), .S(n6), .Q(DP_hold1) );
  OR2X2 U10 ( .A(n8), .B(state[1]), .Y(n36) );
  NAND2X1 U20 ( .A(n17), .B(n18), .Y(n43) );
  AOI22X1 U21 ( .A(DP_hold1), .B(n12), .C(DP1_RX), .D(n19), .Y(n17) );
  NAND2X1 U22 ( .A(n20), .B(n18), .Y(n44) );
  AOI22X1 U23 ( .A(n10), .B(DP_hold1), .C(DP_hold2), .D(n21), .Y(n20) );
  NAND2X1 U24 ( .A(SHIFT_ENABLE), .B(n19), .Y(n21) );
  XNOR2X1 U25 ( .A(DP_hold1), .B(DP_hold2), .Y(D_ORIG) );
  NOR2X1 U26 ( .A(n22), .B(EOP), .Y(N32) );
  AOI21X1 U27 ( .A(n23), .B(BITSTUFF), .C(BS_ERROR), .Y(n22) );
  NAND3X1 U28 ( .A(state[3]), .B(n16), .C(n25), .Y(n24) );
  NOR2X1 U29 ( .A(state[2]), .B(state[1]), .Y(n25) );
  NOR2X1 U30 ( .A(n19), .B(state[3]), .Y(BITSTUFF) );
  NOR2X1 U31 ( .A(n26), .B(n14), .Y(N31) );
  AOI21X1 U32 ( .A(state[2]), .B(n27), .C(n28), .Y(n26) );
  OAI21X1 U33 ( .A(n29), .B(n30), .C(n31), .Y(n28) );
  NAND2X1 U34 ( .A(state[0]), .B(n23), .Y(n30) );
  NAND2X1 U35 ( .A(state[1]), .B(n15), .Y(n29) );
  OAI21X1 U36 ( .A(state[1]), .B(n32), .C(SHIFT_ENABLE), .Y(n27) );
  NOR2X1 U37 ( .A(n33), .B(n14), .Y(N30) );
  AOI21X1 U38 ( .A(state[1]), .B(n34), .C(n35), .Y(n33) );
  OAI21X1 U39 ( .A(n16), .B(n36), .C(n31), .Y(n35) );
  NAND2X1 U40 ( .A(n12), .B(n32), .Y(n31) );
  NAND2X1 U41 ( .A(n13), .B(n16), .Y(n19) );
  OAI21X1 U42 ( .A(n32), .B(n37), .C(SHIFT_ENABLE), .Y(n34) );
  NAND2X1 U43 ( .A(n16), .B(n15), .Y(n37) );
  NOR2X1 U44 ( .A(n38), .B(n14), .Y(N29) );
  NOR2X1 U45 ( .A(EOP), .B(state[3]), .Y(n18) );
  AOI21X1 U46 ( .A(state[0]), .B(n9), .C(n39), .Y(n38) );
  OAI21X1 U47 ( .A(n8), .B(n40), .C(n41), .Y(n39) );
  NAND3X1 U48 ( .A(n13), .B(n32), .C(SHIFT_ENABLE), .Y(n41) );
  NAND2X1 U49 ( .A(n42), .B(n16), .Y(n40) );
  NAND2X1 U50 ( .A(state[2]), .B(state[1]), .Y(n42) );
  NOR2X1 U51 ( .A(n32), .B(n9), .Y(n23) );
  XOR2X1 U52 ( .A(DP1_RX), .B(DP_hold2), .Y(n32) );
  DFFSR \state_reg[3]  ( .D(N32), .CLK(CLK), .R(n6), .S(1'b1), .Q(state[3]) );
  DFFSR \state_reg[0]  ( .D(N29), .CLK(CLK), .R(n6), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[2]  ( .D(N31), .CLK(CLK), .R(n6), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[1]  ( .D(N30), .CLK(CLK), .R(n6), .S(1'b1), .Q(state[1]) );
  INVX2 U8 ( .A(RST), .Y(n6) );
  INVX2 U11 ( .A(n23), .Y(n8) );
  INVX2 U12 ( .A(SHIFT_ENABLE), .Y(n9) );
  INVX2 U13 ( .A(n21), .Y(n10) );
  INVX2 U14 ( .A(n24), .Y(BS_ERROR) );
  INVX2 U15 ( .A(n19), .Y(n12) );
  INVX2 U16 ( .A(n42), .Y(n13) );
  INVX2 U17 ( .A(n18), .Y(n14) );
  INVX2 U18 ( .A(state[2]), .Y(n15) );
  INVX2 U19 ( .A(state[0]), .Y(n16) );
endmodule


module rx_edgedetect_1 ( CLK, RST, DP1_RX, D_EDGE );
  input CLK, RST, DP1_RX;
  output D_EDGE;
  wire   DP_hold1, DP_hold2, n4, n2;

  DFFSR DP_hold1_reg ( .D(DP1_RX), .CLK(CLK), .R(1'b1), .S(n2), .Q(DP_hold1)
         );
  DFFSR DP_hold2_reg ( .D(DP_hold1), .CLK(CLK), .R(1'b1), .S(n2), .Q(DP_hold2)
         );
  NOR2X1 U6 ( .A(RST), .B(n4), .Y(D_EDGE) );
  XNOR2X1 U7 ( .A(DP_hold2), .B(DP_hold1), .Y(n4) );
  INVX2 U4 ( .A(RST), .Y(n2) );
endmodule


module rx_eopdetect_1 ( DP1_RX, DM1_RX, EOP );
  input DP1_RX, DM1_RX;
  output EOP;


  NOR2X1 U1 ( .A(DP1_RX), .B(DM1_RX), .Y(EOP) );
endmodule


module rx_rcu_1 ( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR, 
        RX_CRC, RX_CHECK_CRC, RCV_DATA, RCVING, W_ENABLE, R_ERROR, CRC_ERROR, 
        OPCODE );
  input [15:0] RX_CRC;
  input [15:0] RX_CHECK_CRC;
  input [7:0] RCV_DATA;
  output [1:0] OPCODE;
  input CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR;
  output RCVING, W_ENABLE, R_ERROR, CRC_ERROR;
  wire   n192, nxtR_ERROR, curR_ERROR, curCRC_ERROR, n9, n11, n12, n14, n15,
         n16, n20, n21, n22, n27, n29, n31, n32, n33, n34, n36, n37, n38, n39,
         n40, n41, n42, n45, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56,
         n57, n59, n60, n61, n62, n63, n65, n66, n67, n70, n71, n72, n74, n75,
         n77, n78, n79, n80, n81, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n94, n95, n96, n97, n98, n99, n100, n102, n103, n105, n106, n107,
         n109, n111, n113, n116, n117, n119, n120, n121, n122, n123, n125,
         n126, n127, n129, n133, n134, n136, n137, n138, n139, n140, n142,
         n144, n145, n146, n147, n150, n151, n161, n162, n163, n1, n2, n3, n19,
         n23, n24, n25, n28, n30, n35, n43, n44, n49, n58, n64, n68, n69, n73,
         n76, n82, n93, n101, n104, n108, n110, n112, n114, n115, n118, n124,
         n128, n130, n131, n132, n135, n141, n143, n148, n149, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  wire   [3:0] state;
  wire   [3:0] count;
  wire   [3:0] nextstate;

  DFFPOSX1 curCRC_ERROR_reg ( .D(n151), .CLK(CLK), .Q(curCRC_ERROR) );
  DFFPOSX1 curR_ERROR_reg ( .D(n150), .CLK(CLK), .Q(curR_ERROR) );
  DFFPOSX1 CRC_ERROR_reg ( .D(n169), .CLK(CLK), .Q(CRC_ERROR) );
  OAI21X1 U5 ( .A(EOP), .B(n43), .C(n14), .Y(n12) );
  AOI22X1 U6 ( .A(BS_ERROR), .B(n15), .C(n16), .D(n30), .Y(n14) );
  OAI21X1 U7 ( .A(n191), .B(n25), .C(n20), .Y(n16) );
  AOI22X1 U8 ( .A(n21), .B(D_EDGE), .C(n1), .D(n22), .Y(n20) );
  OAI21X1 U9 ( .A(n181), .B(n189), .C(n182), .Y(n22) );
  NOR2X1 U11 ( .A(n181), .B(n175), .Y(n21) );
  OAI21X1 U12 ( .A(n27), .B(n183), .C(n29), .Y(n15) );
  OAI21X1 U13 ( .A(n3), .B(n31), .C(n32), .Y(n11) );
  NAND2X1 U15 ( .A(n176), .B(n36), .Y(n31) );
  NAND2X1 U16 ( .A(n37), .B(n38), .Y(nextstate[2]) );
  NOR2X1 U17 ( .A(n39), .B(n40), .Y(n38) );
  OAI21X1 U18 ( .A(n25), .B(n41), .C(n34), .Y(n40) );
  OAI21X1 U19 ( .A(n3), .B(n42), .C(n35), .Y(n41) );
  NAND2X1 U20 ( .A(n177), .B(n186), .Y(n42) );
  NAND2X1 U21 ( .A(n45), .B(n46), .Y(n39) );
  NOR2X1 U22 ( .A(n47), .B(n48), .Y(n37) );
  OAI22X1 U23 ( .A(n23), .B(n30), .C(n50), .D(n189), .Y(n48) );
  OAI21X1 U24 ( .A(n35), .B(n51), .C(n52), .Y(n47) );
  OAI21X1 U25 ( .A(n53), .B(n54), .C(n55), .Y(n52) );
  AOI22X1 U26 ( .A(n56), .B(n57), .C(n36), .D(n191), .Y(n51) );
  NOR2X1 U27 ( .A(D_EDGE), .B(n181), .Y(n56) );
  OAI21X1 U28 ( .A(n168), .B(n191), .C(n59), .Y(nextstate[1]) );
  OAI21X1 U30 ( .A(n62), .B(n63), .C(n189), .Y(n60) );
  OAI21X1 U31 ( .A(n29), .B(n178), .C(n65), .Y(n63) );
  OAI21X1 U33 ( .A(n43), .B(n67), .C(n172), .Y(n62) );
  NAND2X1 U34 ( .A(n179), .B(n191), .Y(n67) );
  OAI22X1 U35 ( .A(n70), .B(n71), .C(n30), .D(n72), .Y(nextstate[0]) );
  OAI21X1 U36 ( .A(n181), .B(n24), .C(n74), .Y(n72) );
  NAND3X1 U37 ( .A(n189), .B(n181), .C(n75), .Y(n74) );
  OAI21X1 U38 ( .A(n19), .B(n191), .C(n77), .Y(n75) );
  AOI22X1 U39 ( .A(n66), .B(n78), .C(n79), .D(n80), .Y(n77) );
  OAI22X1 U42 ( .A(state[0]), .B(n182), .C(n81), .D(n181), .Y(n71) );
  AOI22X1 U43 ( .A(EOP), .B(n78), .C(D_EDGE), .D(n171), .Y(n81) );
  OAI21X1 U45 ( .A(state[2]), .B(n84), .C(n85), .Y(n70) );
  NOR2X1 U46 ( .A(n35), .B(n36), .Y(n85) );
  AOI22X1 U47 ( .A(n86), .B(n66), .C(D_EDGE), .D(n78), .Y(n84) );
  NOR2X1 U48 ( .A(n179), .B(EOP), .Y(n66) );
  NOR2X1 U50 ( .A(BS_ERROR), .B(n19), .Y(n86) );
  AOI21X1 U52 ( .A(CRC_ERROR), .B(RST), .C(n88), .Y(n87) );
  OAI21X1 U53 ( .A(n89), .B(n90), .C(n91), .Y(n88) );
  NAND2X1 U54 ( .A(curCRC_ERROR), .B(n92), .Y(n90) );
  NAND2X1 U55 ( .A(n44), .B(n30), .Y(n89) );
  OAI21X1 U56 ( .A(n44), .B(n188), .C(n94), .Y(n150) );
  AOI21X1 U57 ( .A(n9), .B(n44), .C(n170), .Y(n94) );
  NAND3X1 U59 ( .A(n96), .B(n30), .C(curR_ERROR), .Y(n95) );
  OAI21X1 U60 ( .A(n1), .B(n181), .C(n97), .Y(n96) );
  OAI21X1 U61 ( .A(n176), .B(n25), .C(n98), .Y(n9) );
  OAI21X1 U64 ( .A(n1), .B(n80), .C(n175), .Y(n100) );
  OAI21X1 U65 ( .A(n54), .B(n173), .C(EOP), .Y(n99) );
  OAI21X1 U69 ( .A(n103), .B(n187), .C(n91), .Y(n151) );
  NAND3X1 U70 ( .A(n3), .B(n44), .C(n105), .Y(n91) );
  NOR2X1 U71 ( .A(n25), .B(n102), .Y(n105) );
  NAND3X1 U72 ( .A(n35), .B(n186), .C(n177), .Y(n102) );
  AOI21X1 U76 ( .A(n92), .B(n30), .C(RST), .Y(n103) );
  OAI21X1 U77 ( .A(n181), .B(n19), .C(n97), .Y(n92) );
  NAND2X1 U78 ( .A(n27), .B(n83), .Y(n97) );
  NOR2X1 U79 ( .A(D_EDGE), .B(state[2]), .Y(n83) );
  OAI21X1 U81 ( .A(n107), .B(n184), .C(n109), .Y(n161) );
  NAND3X1 U82 ( .A(n160), .B(n184), .C(count[0]), .Y(n109) );
  AOI21X1 U83 ( .A(n111), .B(n180), .C(n113), .Y(n107) );
  OAI21X1 U84 ( .A(n157), .B(n185), .C(n116), .Y(n162) );
  NAND3X1 U85 ( .A(n117), .B(n185), .C(n158), .Y(n116) );
  OAI21X1 U87 ( .A(n120), .B(n186), .C(n121), .Y(n163) );
  NAND3X1 U88 ( .A(n117), .B(n186), .C(n122), .Y(n121) );
  NOR2X1 U89 ( .A(n123), .B(n185), .Y(n122) );
  AOI21X1 U90 ( .A(n111), .B(n185), .C(n119), .Y(n120) );
  OAI21X1 U91 ( .A(n158), .B(n166), .C(n46), .Y(n119) );
  NAND3X1 U93 ( .A(count[1]), .B(count[0]), .C(n125), .Y(n123) );
  AOI22X1 U95 ( .A(n113), .B(count[0]), .C(n180), .D(n160), .Y(n126) );
  NAND3X1 U97 ( .A(n117), .B(n190), .C(SHIFT_ENABLE), .Y(n127) );
  OAI21X1 U100 ( .A(n125), .B(n166), .C(n46), .Y(n113) );
  NAND2X1 U101 ( .A(EOP), .B(n129), .Y(n46) );
  NOR2X1 U103 ( .A(n55), .B(n167), .Y(n111) );
  NOR2X1 U104 ( .A(n186), .B(n106), .Y(n55) );
  NAND3X1 U105 ( .A(n184), .B(n185), .C(n180), .Y(n106) );
  NOR2X1 U110 ( .A(BITSTUFF), .B(n159), .Y(n125) );
  NAND3X1 U115 ( .A(n134), .B(n164), .C(n79), .Y(n33) );
  NAND3X1 U117 ( .A(n136), .B(n137), .C(n138), .Y(n80) );
  NOR2X1 U119 ( .A(RCV_DATA[6]), .B(RCV_DATA[5]), .Y(n140) );
  NOR2X1 U120 ( .A(RCV_DATA[4]), .B(RCV_DATA[3]), .Y(n139) );
  NOR2X1 U121 ( .A(RCV_DATA[2]), .B(RCV_DATA[1]), .Y(n137) );
  NOR2X1 U122 ( .A(RCV_DATA[0]), .B(n165), .Y(n136) );
  NAND3X1 U124 ( .A(n168), .B(n61), .C(n50), .Y(RCVING) );
  NOR2X1 U125 ( .A(n129), .B(n142), .Y(n50) );
  OAI21X1 U126 ( .A(n183), .B(n174), .C(n133), .Y(n142) );
  NAND3X1 U127 ( .A(state[2]), .B(n30), .C(n27), .Y(n133) );
  OAI21X1 U129 ( .A(n35), .B(n25), .C(n34), .Y(n144) );
  NAND3X1 U130 ( .A(state[2]), .B(n30), .C(n78), .Y(n34) );
  NAND3X1 U133 ( .A(n43), .B(n29), .C(n172), .Y(n129) );
  NOR2X1 U135 ( .A(n19), .B(n183), .Y(n53) );
  NAND3X1 U137 ( .A(n30), .B(n181), .C(n57), .Y(n29) );
  NOR2X1 U141 ( .A(n30), .B(state[2]), .Y(n134) );
  NOR2X1 U143 ( .A(n175), .B(n171), .Y(n78) );
  OAI21X1 U144 ( .A(n181), .B(n23), .C(n30), .Y(n146) );
  OAI21X1 U148 ( .A(n147), .B(n1), .C(n35), .Y(n145) );
  NOR2X1 U149 ( .A(state[0]), .B(n181), .Y(n147) );
  OAI21X1 U150 ( .A(n30), .B(n25), .C(n61), .Y(n192) );
  NAND3X1 U151 ( .A(n35), .B(state[2]), .C(n57), .Y(n61) );
  NOR2X1 U155 ( .A(n174), .B(n181), .Y(n36) );
  NOR2X1 U158 ( .A(state[0]), .B(n1), .Y(n79) );
  OR2X2 U3 ( .A(n9), .B(n170), .Y(nxtR_ERROR) );
  OR2X2 U4 ( .A(n11), .B(n12), .Y(nextstate[3]) );
  AND2X2 U14 ( .A(n33), .B(n34), .Y(n32) );
  AND2X2 U29 ( .A(n60), .B(n61), .Y(n59) );
  AND2X2 U62 ( .A(n99), .B(n45), .Y(n98) );
  OR2X2 U63 ( .A(n183), .B(n100), .Y(n45) );
  AND2X2 U99 ( .A(n111), .B(n46), .Y(n117) );
  AND2X2 U114 ( .A(n33), .B(n133), .Y(n65) );
  AND2X2 U118 ( .A(n139), .B(n140), .Y(n138) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        state[0]) );
  DFFSR R_ERROR_reg ( .D(nxtR_ERROR), .CLK(CLK), .R(n44), .S(1'b1), .Q(R_ERROR) );
  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        state[2]) );
  DFFSR \count_reg[0]  ( .D(n156), .CLK(CLK), .R(n44), .S(1'b1), .Q(count[0])
         );
  DFFSR \count_reg[1]  ( .D(n161), .CLK(CLK), .R(n44), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n162), .CLK(CLK), .R(n44), .S(1'b1), .Q(count[2])
         );
  DFFSR \count_reg[3]  ( .D(n163), .CLK(CLK), .R(n44), .S(1'b1), .Q(count[3])
         );
  BUFX2 U10 ( .A(state[3]), .Y(n1) );
  INVX2 U32 ( .A(state[0]), .Y(n175) );
  AND2X2 U40 ( .A(n146), .B(n145), .Y(n2) );
  NAND2X1 U41 ( .A(n152), .B(n149), .Y(n3) );
  INVX2 U75 ( .A(n1), .Y(n171) );
  OR2X2 U80 ( .A(n175), .B(n1), .Y(n19) );
  INVX2 U86 ( .A(n19), .Y(n57) );
  OR2X2 U92 ( .A(n171), .B(state[0]), .Y(n23) );
  INVX2 U94 ( .A(n23), .Y(n27) );
  NAND2X1 U96 ( .A(n167), .B(n2), .Y(OPCODE[1]) );
  OR2X2 U98 ( .A(n175), .B(n171), .Y(n24) );
  INVX2 U102 ( .A(state[2]), .Y(n181) );
  OR2X2 U106 ( .A(n174), .B(n181), .Y(n25) );
  OAI21X1 U107 ( .A(n30), .B(n25), .C(n61), .Y(OPCODE[0]) );
  INVX2 U108 ( .A(n65), .Y(n28) );
  OR2X2 U109 ( .A(n28), .B(n192), .Y(W_ENABLE) );
  INVX2 U111 ( .A(RST), .Y(n44) );
  INVX2 U112 ( .A(n134), .Y(n183) );
  INVX2 U113 ( .A(state[1]), .Y(n30) );
  INVX1 U116 ( .A(n30), .Y(n35) );
  OR2X2 U123 ( .A(n24), .B(n183), .Y(n43) );
  INVX1 U128 ( .A(n43), .Y(n54) );
  XNOR2X1 U131 ( .A(RX_CHECK_CRC[10]), .B(RX_CRC[10]), .Y(n69) );
  XNOR2X1 U132 ( .A(RX_CHECK_CRC[9]), .B(RX_CRC[9]), .Y(n68) );
  XOR2X1 U134 ( .A(RX_CHECK_CRC[7]), .B(RX_CRC[7]), .Y(n58) );
  XOR2X1 U136 ( .A(RX_CHECK_CRC[8]), .B(RX_CRC[8]), .Y(n49) );
  NOR2X1 U138 ( .A(n58), .B(n49), .Y(n64) );
  NAND3X1 U139 ( .A(n69), .B(n68), .C(n64), .Y(n108) );
  XNOR2X1 U140 ( .A(RX_CHECK_CRC[14]), .B(RX_CRC[14]), .Y(n101) );
  XNOR2X1 U142 ( .A(RX_CHECK_CRC[13]), .B(RX_CRC[13]), .Y(n93) );
  XOR2X1 U145 ( .A(RX_CHECK_CRC[11]), .B(RX_CRC[11]), .Y(n76) );
  XOR2X1 U146 ( .A(RX_CHECK_CRC[12]), .B(RX_CRC[12]), .Y(n73) );
  NOR2X1 U147 ( .A(n76), .B(n73), .Y(n82) );
  NAND3X1 U152 ( .A(n101), .B(n93), .C(n82), .Y(n104) );
  NOR2X1 U153 ( .A(n108), .B(n104), .Y(n152) );
  NOR2X1 U154 ( .A(n153), .B(RX_CHECK_CRC[0]), .Y(n110) );
  OAI22X1 U156 ( .A(RX_CRC[1]), .B(n110), .C(n110), .D(n155), .Y(n128) );
  AND2X1 U157 ( .A(RX_CHECK_CRC[0]), .B(n153), .Y(n112) );
  OAI22X1 U159 ( .A(n112), .B(n154), .C(RX_CHECK_CRC[1]), .D(n112), .Y(n124)
         );
  XOR2X1 U160 ( .A(RX_CHECK_CRC[15]), .B(RX_CRC[15]), .Y(n115) );
  XOR2X1 U161 ( .A(RX_CHECK_CRC[2]), .B(RX_CRC[2]), .Y(n114) );
  NOR2X1 U162 ( .A(n115), .B(n114), .Y(n118) );
  NAND3X1 U163 ( .A(n128), .B(n124), .C(n118), .Y(n148) );
  XNOR2X1 U164 ( .A(RX_CHECK_CRC[6]), .B(RX_CRC[6]), .Y(n141) );
  XNOR2X1 U165 ( .A(RX_CHECK_CRC[5]), .B(RX_CRC[5]), .Y(n135) );
  XOR2X1 U166 ( .A(RX_CHECK_CRC[3]), .B(RX_CRC[3]), .Y(n131) );
  XOR2X1 U167 ( .A(RX_CHECK_CRC[4]), .B(RX_CRC[4]), .Y(n130) );
  NOR2X1 U168 ( .A(n131), .B(n130), .Y(n132) );
  NAND3X1 U169 ( .A(n141), .B(n135), .C(n132), .Y(n143) );
  NOR2X1 U170 ( .A(n148), .B(n143), .Y(n149) );
  INVX2 U171 ( .A(RX_CRC[0]), .Y(n153) );
  INVX2 U172 ( .A(RX_CRC[1]), .Y(n154) );
  INVX2 U173 ( .A(RX_CHECK_CRC[1]), .Y(n155) );
  INVX2 U174 ( .A(n126), .Y(n156) );
  INVX2 U175 ( .A(n119), .Y(n157) );
  INVX2 U176 ( .A(n123), .Y(n158) );
  INVX2 U177 ( .A(SHIFT_ENABLE), .Y(n159) );
  INVX2 U178 ( .A(n127), .Y(n160) );
  INVX2 U179 ( .A(n80), .Y(n164) );
  INVX2 U180 ( .A(RCV_DATA[7]), .Y(n165) );
  INVX2 U181 ( .A(n111), .Y(n166) );
  INVX2 U182 ( .A(n129), .Y(n167) );
  INVX2 U183 ( .A(n144), .Y(n168) );
  INVX2 U184 ( .A(n87), .Y(n169) );
  INVX2 U185 ( .A(n95), .Y(n170) );
  INVX2 U186 ( .A(n53), .Y(n172) );
  INVX2 U187 ( .A(n29), .Y(n173) );
  INVX2 U188 ( .A(n79), .Y(n174) );
  INVX2 U189 ( .A(n102), .Y(n176) );
  INVX2 U190 ( .A(n106), .Y(n177) );
  INVX2 U191 ( .A(n66), .Y(n178) );
  INVX2 U192 ( .A(n55), .Y(n179) );
  INVX2 U193 ( .A(count[0]), .Y(n180) );
  INVX2 U194 ( .A(n83), .Y(n182) );
  INVX2 U195 ( .A(count[1]), .Y(n184) );
  INVX2 U196 ( .A(count[2]), .Y(n185) );
  INVX2 U197 ( .A(count[3]), .Y(n186) );
  INVX2 U198 ( .A(curCRC_ERROR), .Y(n187) );
  INVX2 U199 ( .A(curR_ERROR), .Y(n188) );
  INVX2 U200 ( .A(BS_ERROR), .Y(n189) );
  INVX2 U201 ( .A(BITSTUFF), .Y(n190) );
  INVX2 U202 ( .A(EOP), .Y(n191) );
endmodule


module rx_shift_reg_1 ( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF, RCV_DATA );
  output [7:0] RCV_DATA;
  input CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF;
  wire   n2, n4, n6, n8, n10, n12, n14, n16, n18, n19, n21, n23, n24, n26, n27,
         n29, n30, n32, n33, n35, n36, n38, n39, n41, n42, n44, n17, n20, n22,
         n25, n28, n31, n34, n37, n40, n43, n45;
  wire   [7:0] present_val;

  DFFPOSX1 \RCV_DATA_reg[7]  ( .D(n42), .CLK(CLK), .Q(RCV_DATA[7]) );
  DFFPOSX1 \RCV_DATA_reg[6]  ( .D(n39), .CLK(CLK), .Q(RCV_DATA[6]) );
  DFFPOSX1 \RCV_DATA_reg[5]  ( .D(n36), .CLK(CLK), .Q(RCV_DATA[5]) );
  DFFPOSX1 \RCV_DATA_reg[4]  ( .D(n33), .CLK(CLK), .Q(RCV_DATA[4]) );
  DFFPOSX1 \RCV_DATA_reg[3]  ( .D(n30), .CLK(CLK), .Q(RCV_DATA[3]) );
  DFFPOSX1 \RCV_DATA_reg[2]  ( .D(n27), .CLK(CLK), .Q(RCV_DATA[2]) );
  DFFPOSX1 \RCV_DATA_reg[1]  ( .D(n24), .CLK(CLK), .Q(RCV_DATA[1]) );
  DFFPOSX1 \RCV_DATA_reg[0]  ( .D(n21), .CLK(CLK), .Q(RCV_DATA[0]) );
  OAI21X1 U2 ( .A(RST), .B(n43), .C(n2), .Y(n21) );
  NAND2X1 U3 ( .A(RCV_DATA[0]), .B(RST), .Y(n2) );
  OAI22X1 U4 ( .A(n20), .B(n43), .C(n4), .D(n40), .Y(n23) );
  OAI21X1 U6 ( .A(RST), .B(n40), .C(n6), .Y(n24) );
  NAND2X1 U7 ( .A(RCV_DATA[1]), .B(RST), .Y(n6) );
  OAI22X1 U8 ( .A(n20), .B(n40), .C(n4), .D(n37), .Y(n26) );
  OAI21X1 U10 ( .A(RST), .B(n37), .C(n8), .Y(n27) );
  NAND2X1 U11 ( .A(RCV_DATA[2]), .B(RST), .Y(n8) );
  OAI22X1 U12 ( .A(n20), .B(n37), .C(n4), .D(n34), .Y(n29) );
  OAI21X1 U14 ( .A(RST), .B(n34), .C(n10), .Y(n30) );
  NAND2X1 U15 ( .A(RCV_DATA[3]), .B(RST), .Y(n10) );
  OAI22X1 U16 ( .A(n20), .B(n34), .C(n4), .D(n31), .Y(n32) );
  OAI21X1 U18 ( .A(RST), .B(n31), .C(n12), .Y(n33) );
  NAND2X1 U19 ( .A(RCV_DATA[4]), .B(RST), .Y(n12) );
  OAI22X1 U20 ( .A(n20), .B(n31), .C(n4), .D(n28), .Y(n35) );
  OAI21X1 U22 ( .A(RST), .B(n28), .C(n14), .Y(n36) );
  NAND2X1 U23 ( .A(RCV_DATA[5]), .B(RST), .Y(n14) );
  OAI22X1 U24 ( .A(n20), .B(n28), .C(n4), .D(n25), .Y(n38) );
  OAI21X1 U26 ( .A(RST), .B(n25), .C(n16), .Y(n39) );
  NAND2X1 U27 ( .A(RCV_DATA[6]), .B(RST), .Y(n16) );
  OAI22X1 U28 ( .A(n20), .B(n25), .C(n4), .D(n22), .Y(n41) );
  OAI21X1 U30 ( .A(RST), .B(n22), .C(n18), .Y(n42) );
  NAND2X1 U31 ( .A(RCV_DATA[7]), .B(RST), .Y(n18) );
  OAI21X1 U32 ( .A(n20), .B(n22), .C(n19), .Y(n44) );
  NAND2X1 U33 ( .A(D_ORIG), .B(n20), .Y(n19) );
  NAND2X1 U36 ( .A(SHIFT_ENABLE), .B(n45), .Y(n4) );
  DFFSR \present_val_reg[7]  ( .D(n44), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[7]) );
  DFFSR \present_val_reg[6]  ( .D(n41), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[6]) );
  DFFSR \present_val_reg[5]  ( .D(n38), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[5]) );
  DFFSR \present_val_reg[4]  ( .D(n35), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[4]) );
  DFFSR \present_val_reg[3]  ( .D(n32), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[3]) );
  DFFSR \present_val_reg[2]  ( .D(n29), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[2]) );
  DFFSR \present_val_reg[1]  ( .D(n26), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[1]) );
  DFFSR \present_val_reg[0]  ( .D(n23), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[0]) );
  INVX2 U5 ( .A(n4), .Y(n20) );
  INVX2 U37 ( .A(RST), .Y(n17) );
  INVX2 U38 ( .A(present_val[7]), .Y(n22) );
  INVX2 U39 ( .A(present_val[6]), .Y(n25) );
  INVX2 U40 ( .A(present_val[5]), .Y(n28) );
  INVX2 U41 ( .A(present_val[4]), .Y(n31) );
  INVX2 U42 ( .A(present_val[3]), .Y(n34) );
  INVX2 U43 ( .A(present_val[2]), .Y(n37) );
  INVX2 U44 ( .A(present_val[1]), .Y(n40) );
  INVX2 U45 ( .A(present_val[0]), .Y(n43) );
  INVX2 U46 ( .A(BITSTUFF), .Y(n45) );
endmodule


module rx_timer_1 ( CLK, RST, D_EDGE, RCVING, SHIFT_ENABLE );
  input CLK, RST, D_EDGE, RCVING;
  output SHIFT_ENABLE;
  wire   state, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n6, n7,
         n8, n9, n10, n11, n12, n24, n25;
  wire   [3:0] count;
  wire   [3:0] nextcount;

  AND2X2 U9 ( .A(n25), .B(state), .Y(n19) );
  NOR2X1 U17 ( .A(n13), .B(n14), .Y(nextcount[3]) );
  AOI22X1 U18 ( .A(n15), .B(n16), .C(n17), .D(count[3]), .Y(n13) );
  XOR2X1 U19 ( .A(n18), .B(n16), .Y(n17) );
  NOR2X1 U20 ( .A(count[3]), .B(n11), .Y(n15) );
  AOI21X1 U21 ( .A(n19), .B(n20), .C(n24), .Y(nextcount[2]) );
  XOR2X1 U22 ( .A(n21), .B(count[2]), .Y(n20) );
  NOR2X1 U23 ( .A(n22), .B(n14), .Y(nextcount[1]) );
  NAND2X1 U24 ( .A(state), .B(n23), .Y(nextcount[0]) );
  OAI21X1 U25 ( .A(D_EDGE), .B(n10), .C(RCVING), .Y(n23) );
  NAND3X1 U28 ( .A(RCVING), .B(n25), .C(state), .Y(n14) );
  OAI21X1 U29 ( .A(n22), .B(n12), .C(n21), .Y(n18) );
  NAND2X1 U30 ( .A(count[0]), .B(count[1]), .Y(n21) );
  XOR2X1 U31 ( .A(n12), .B(n22), .Y(n16) );
  XNOR2X1 U32 ( .A(count[0]), .B(count[1]), .Y(n22) );
  DFFSR state_reg ( .D(RCVING), .CLK(CLK), .R(n8), .S(1'b1), .Q(state) );
  DFFSR \count_reg[2]  ( .D(nextcount[2]), .CLK(CLK), .R(n8), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[0]  ( .D(nextcount[0]), .CLK(CLK), .R(n8), .S(1'b1), .Q(
        count[0]) );
  DFFSR \count_reg[3]  ( .D(nextcount[3]), .CLK(CLK), .R(n8), .S(1'b1), .Q(
        count[3]) );
  DFFSR \count_reg[1]  ( .D(nextcount[1]), .CLK(CLK), .R(n8), .S(1'b1), .Q(
        count[1]) );
  INVX2 U8 ( .A(RST), .Y(n8) );
  AND2X2 U10 ( .A(n6), .B(n7), .Y(SHIFT_ENABLE) );
  NOR2X1 U11 ( .A(n16), .B(n18), .Y(n6) );
  AND2X2 U12 ( .A(n9), .B(count[3]), .Y(n7) );
  INVX2 U13 ( .A(n14), .Y(n9) );
  INVX2 U14 ( .A(count[0]), .Y(n10) );
  INVX2 U15 ( .A(n18), .Y(n11) );
  INVX2 U16 ( .A(count[2]), .Y(n12) );
  INVX2 U26 ( .A(RCVING), .Y(n24) );
  INVX2 U27 ( .A(D_EDGE), .Y(n25) );
endmodule


module receiver_block_rewire_1 ( CLK, DM1_RX, DP1_RX, RST, BS_ERROR, CRC_ERROR, 
        EOP_external, OPCODE, RCV_DATA, R_ERROR, W_ENABLE );
  output [1:0] OPCODE;
  output [7:0] RCV_DATA;
  input CLK, DM1_RX, DP1_RX, RST;
  output BS_ERROR, CRC_ERROR, EOP_external, R_ERROR, W_ENABLE;
  wire   SHIFT_ENABLE, BITSTUFF, D_ORIG, D_EDGE, RCVING, n1, n2;
  wire   [15:0] RX_CRC;
  wire   [15:0] rx_CHECK_CRC;

  rx_CRC_CALC_1 U_2 ( .CLK(CLK), .RST(n1), .W_ENABLE(W_ENABLE), .OPCODE(OPCODE), .RCV_DATA(RCV_DATA), .RX_CRC(RX_CRC) );
  rx_accumulator_1 U_3 ( .CLK(CLK), .RST(n1), .RCV_DATA(RCV_DATA), .W_ENABLE(
        W_ENABLE), .rx_CHECK_CRC(rx_CHECK_CRC) );
  rx_decode_1 U_1 ( .CLK(CLK), .RST(n1), .DP1_RX(DP1_RX), .SHIFT_ENABLE(
        SHIFT_ENABLE), .EOP(EOP_external), .D_ORIG(D_ORIG), .BITSTUFF(BITSTUFF), .BS_ERROR(BS_ERROR) );
  rx_edgedetect_1 U_0 ( .CLK(CLK), .RST(n1), .DP1_RX(DP1_RX), .D_EDGE(D_EDGE)
         );
  rx_eopdetect_1 U_4 ( .DP1_RX(DP1_RX), .DM1_RX(DM1_RX), .EOP(EOP_external) );
  rx_rcu_1 U_5 ( .CLK(CLK), .RST(n1), .D_EDGE(D_EDGE), .EOP(EOP_external), 
        .SHIFT_ENABLE(SHIFT_ENABLE), .BITSTUFF(BITSTUFF), .BS_ERROR(BS_ERROR), 
        .RX_CRC(RX_CRC), .RX_CHECK_CRC(rx_CHECK_CRC), .RCV_DATA(RCV_DATA), 
        .RCVING(RCVING), .W_ENABLE(W_ENABLE), .R_ERROR(R_ERROR), .CRC_ERROR(
        CRC_ERROR), .OPCODE(OPCODE) );
  rx_shift_reg_1 U_6 ( .CLK(CLK), .RST(n1), .SHIFT_ENABLE(SHIFT_ENABLE), 
        .D_ORIG(D_ORIG), .BITSTUFF(BITSTUFF), .RCV_DATA(RCV_DATA) );
  rx_timer_1 U_7 ( .CLK(CLK), .RST(n1), .D_EDGE(D_EDGE), .RCVING(RCVING), 
        .SHIFT_ENABLE(SHIFT_ENABLE) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module tx_CRC_CALC_1 ( CLK, RST, EOP, T_STROBE, PRGA_OPCODE, PRGA_OUT, TX_CRC
 );
  input [1:0] PRGA_OPCODE;
  input [7:0] PRGA_OUT;
  output [15:0] TX_CRC;
  input CLK, RST, EOP, T_STROBE;
  wire   n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n1,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n79, n80, n81;

  OAI22X1 U39 ( .A(n25), .B(n20), .C(n38), .D(n19), .Y(n63) );
  XNOR2X1 U40 ( .A(n40), .B(n80), .Y(n38) );
  OAI22X1 U41 ( .A(n79), .B(n20), .C(n19), .D(n37), .Y(n64) );
  OAI22X1 U42 ( .A(n36), .B(n20), .C(n19), .D(n35), .Y(n65) );
  OAI22X1 U43 ( .A(n34), .B(n20), .C(n19), .D(n33), .Y(n66) );
  OAI22X1 U44 ( .A(n32), .B(n20), .C(n19), .D(n31), .Y(n67) );
  OAI22X1 U45 ( .A(n29), .B(n20), .C(n19), .D(n28), .Y(n68) );
  OAI22X1 U46 ( .A(n27), .B(n20), .C(n41), .D(n19), .Y(n69) );
  XNOR2X1 U47 ( .A(TX_CRC[1]), .B(n42), .Y(n41) );
  OAI22X1 U48 ( .A(n24), .B(n20), .C(n43), .D(n19), .Y(n70) );
  XOR2X1 U49 ( .A(n44), .B(n45), .Y(n43) );
  XNOR2X1 U50 ( .A(TX_CRC[0]), .B(n42), .Y(n44) );
  OAI22X1 U51 ( .A(n80), .B(n20), .C(n46), .D(n19), .Y(n71) );
  OAI22X1 U52 ( .A(n20), .B(n37), .C(n47), .D(n19), .Y(n72) );
  XNOR2X1 U53 ( .A(n48), .B(n49), .Y(n47) );
  OAI22X1 U54 ( .A(n20), .B(n35), .C(n50), .D(n39), .Y(n73) );
  OAI22X1 U55 ( .A(n20), .B(n33), .C(n51), .D(n39), .Y(n74) );
  XNOR2X1 U56 ( .A(n52), .B(n53), .Y(n51) );
  OAI22X1 U57 ( .A(n20), .B(n31), .C(n54), .D(n39), .Y(n75) );
  OAI22X1 U58 ( .A(n20), .B(n28), .C(n55), .D(n39), .Y(n76) );
  XOR2X1 U59 ( .A(n56), .B(n57), .Y(n55) );
  OAI22X1 U60 ( .A(n20), .B(n26), .C(n58), .D(n39), .Y(n77) );
  XOR2X1 U61 ( .A(n59), .B(n60), .Y(n58) );
  XOR2X1 U62 ( .A(n42), .B(n46), .Y(n59) );
  OAI22X1 U63 ( .A(n20), .B(n23), .C(n40), .D(n39), .Y(n78) );
  XOR2X1 U64 ( .A(n61), .B(n62), .Y(n40) );
  XOR2X1 U65 ( .A(n57), .B(n42), .Y(n62) );
  XNOR2X1 U66 ( .A(n25), .B(PRGA_OUT[7]), .Y(n42) );
  XNOR2X1 U67 ( .A(n24), .B(PRGA_OUT[0]), .Y(n57) );
  XOR2X1 U68 ( .A(n46), .B(n60), .Y(n61) );
  XOR2X1 U69 ( .A(n54), .B(n50), .Y(n60) );
  XNOR2X1 U70 ( .A(n53), .B(n48), .Y(n50) );
  XOR2X1 U71 ( .A(TX_CRC[12]), .B(PRGA_OUT[4]), .Y(n48) );
  XOR2X1 U72 ( .A(TX_CRC[11]), .B(PRGA_OUT[3]), .Y(n53) );
  XNOR2X1 U73 ( .A(n56), .B(n30), .Y(n54) );
  XOR2X1 U74 ( .A(TX_CRC[10]), .B(PRGA_OUT[2]), .Y(n52) );
  XNOR2X1 U75 ( .A(TX_CRC[9]), .B(PRGA_OUT[1]), .Y(n56) );
  XNOR2X1 U76 ( .A(n49), .B(n45), .Y(n46) );
  XNOR2X1 U77 ( .A(n79), .B(PRGA_OUT[6]), .Y(n45) );
  XOR2X1 U78 ( .A(TX_CRC[13]), .B(PRGA_OUT[5]), .Y(n49) );
  NAND3X1 U80 ( .A(PRGA_OPCODE[0]), .B(n81), .C(T_STROBE), .Y(n39) );
  DFFSR \current_crc_reg[6]  ( .D(n72), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[6]) );
  DFFSR \current_crc_reg[5]  ( .D(n73), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[5]) );
  DFFSR \current_crc_reg[4]  ( .D(n74), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[4]) );
  DFFSR \current_crc_reg[3]  ( .D(n75), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[3]) );
  DFFSR \current_crc_reg[2]  ( .D(n76), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[2]) );
  DFFSR \current_crc_reg[1]  ( .D(n77), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[1]) );
  DFFSR \current_crc_reg[0]  ( .D(n78), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[0]) );
  DFFSR \current_crc_reg[15]  ( .D(n63), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[15]) );
  DFFSR \current_crc_reg[14]  ( .D(n64), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[14]) );
  DFFSR \current_crc_reg[13]  ( .D(n65), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[13]) );
  DFFSR \current_crc_reg[12]  ( .D(n66), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[12]) );
  DFFSR \current_crc_reg[11]  ( .D(n67), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[11]) );
  DFFSR \current_crc_reg[10]  ( .D(n68), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[10]) );
  DFFSR \current_crc_reg[9]  ( .D(n69), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[9]) );
  DFFSR \current_crc_reg[8]  ( .D(n70), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[8]) );
  DFFSR \current_crc_reg[7]  ( .D(n71), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[7]) );
  AND2X2 U3 ( .A(n19), .B(n22), .Y(n1) );
  INVX2 U20 ( .A(n1), .Y(n20) );
  INVX2 U21 ( .A(RST), .Y(n21) );
  INVX2 U22 ( .A(n18), .Y(n19) );
  INVX2 U23 ( .A(n39), .Y(n18) );
  INVX2 U24 ( .A(EOP), .Y(n22) );
  INVX2 U25 ( .A(TX_CRC[0]), .Y(n23) );
  INVX2 U26 ( .A(TX_CRC[8]), .Y(n24) );
  INVX2 U27 ( .A(TX_CRC[15]), .Y(n25) );
  INVX2 U28 ( .A(TX_CRC[1]), .Y(n26) );
  INVX2 U29 ( .A(TX_CRC[9]), .Y(n27) );
  INVX2 U30 ( .A(TX_CRC[2]), .Y(n28) );
  INVX2 U31 ( .A(TX_CRC[10]), .Y(n29) );
  INVX2 U32 ( .A(n52), .Y(n30) );
  INVX2 U33 ( .A(TX_CRC[3]), .Y(n31) );
  INVX2 U34 ( .A(TX_CRC[11]), .Y(n32) );
  INVX2 U35 ( .A(TX_CRC[4]), .Y(n33) );
  INVX2 U36 ( .A(TX_CRC[12]), .Y(n34) );
  INVX2 U37 ( .A(TX_CRC[5]), .Y(n35) );
  INVX2 U38 ( .A(TX_CRC[13]), .Y(n36) );
  INVX2 U79 ( .A(TX_CRC[6]), .Y(n37) );
  INVX2 U81 ( .A(TX_CRC[14]), .Y(n79) );
  INVX2 U82 ( .A(TX_CRC[7]), .Y(n80) );
  INVX2 U83 ( .A(PRGA_OPCODE[1]), .Y(n81) );
endmodule


module tx_encode_1 ( clk, rst, SHIFT_ENABLE_E, d_encode, EOP, t_bitstuff, 
        dp_tx_out, dm_tx_out );
  input clk, rst, SHIFT_ENABLE_E, d_encode, EOP;
  output t_bitstuff, dp_tx_out, dm_tx_out;
  wire   DE_holdout, DE_holdout_BS, DE_holdout_last, DE_holdout_nxt, dm_tx_nxt,
         n1, n3, n5, n6, n9, n12, n13, n14, n15, n18, n19, n20, n22, n23, n24,
         n26, n27, n32, n33, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n61, n64, n16, n17, n21, n25, n28, n29,
         n30, n31, n34, n35, n42, n53, n54, n56, n57, n58, n59, n60, n63;
  wire   [3:0] state;
  wire   [3:0] nextstate;

  DFFSR DE_holdout_reg ( .D(DE_holdout_nxt), .CLK(clk), .R(1'b1), .S(n16), .Q(
        DE_holdout) );
  DFFPOSX1 DE_holdout_last_reg ( .D(n61), .CLK(clk), .Q(DE_holdout_last) );
  DFFSR dp_tx_out_reg ( .D(DE_holdout_nxt), .CLK(clk), .R(1'b1), .S(n16), .Q(
        dp_tx_out) );
  AOI21X1 U3 ( .A(state[3]), .B(n1), .C(n30), .Y(nextstate[3]) );
  OAI21X1 U4 ( .A(n3), .B(n60), .C(n5), .Y(nextstate[2]) );
  AOI21X1 U5 ( .A(n6), .B(n17), .C(n34), .Y(n5) );
  NOR2X1 U7 ( .A(state[2]), .B(n59), .Y(n6) );
  AOI21X1 U8 ( .A(n35), .B(n59), .C(n12), .Y(n3) );
  OAI21X1 U9 ( .A(state[1]), .B(n9), .C(n13), .Y(nextstate[1]) );
  AOI21X1 U10 ( .A(state[1]), .B(n14), .C(n34), .Y(n13) );
  OAI21X1 U11 ( .A(state[0]), .B(n15), .C(n21), .Y(n14) );
  NAND3X1 U12 ( .A(SHIFT_ENABLE_E), .B(n35), .C(state[0]), .Y(n9) );
  OAI21X1 U14 ( .A(n58), .B(n21), .C(n18), .Y(nextstate[0]) );
  OAI21X1 U15 ( .A(n19), .B(n20), .C(SHIFT_ENABLE_E), .Y(n18) );
  OAI21X1 U16 ( .A(n31), .B(n22), .C(n23), .Y(n20) );
  NAND2X1 U17 ( .A(n24), .B(n42), .Y(n22) );
  NOR2X1 U18 ( .A(state[0]), .B(n15), .Y(n19) );
  NAND3X1 U19 ( .A(d_encode), .B(n26), .C(n27), .Y(n15) );
  XNOR2X1 U20 ( .A(n54), .B(n53), .Y(n27) );
  NOR2X1 U22 ( .A(n31), .B(SHIFT_ENABLE_E), .Y(n12) );
  OAI22X1 U23 ( .A(n16), .B(n54), .C(rst), .D(n53), .Y(n61) );
  OAI22X1 U26 ( .A(n25), .B(n63), .C(n53), .D(n32), .Y(n64) );
  NAND2X1 U28 ( .A(n34), .B(SHIFT_ENABLE_E), .Y(n32) );
  NAND3X1 U30 ( .A(n24), .B(n58), .C(n26), .Y(n23) );
  NOR2X1 U31 ( .A(state[3]), .B(n33), .Y(t_bitstuff) );
  OAI21X1 U32 ( .A(n57), .B(n56), .C(n36), .Y(dm_tx_nxt) );
  AOI22X1 U33 ( .A(n37), .B(n24), .C(n38), .D(n39), .Y(n36) );
  NOR2X1 U34 ( .A(n24), .B(n31), .Y(n38) );
  NOR2X1 U36 ( .A(EOP), .B(state[3]), .Y(n26) );
  NOR2X1 U37 ( .A(EOP), .B(n40), .Y(n37) );
  AOI22X1 U38 ( .A(state[0]), .B(n41), .C(n28), .D(n58), .Y(n40) );
  XNOR2X1 U40 ( .A(DE_holdout_BS), .B(n44), .Y(n41) );
  OAI21X1 U41 ( .A(n57), .B(n56), .C(n45), .Y(DE_holdout_nxt) );
  OAI21X1 U42 ( .A(n46), .B(n47), .C(n30), .Y(n45) );
  OAI21X1 U44 ( .A(n24), .B(n39), .C(n48), .Y(n47) );
  NAND3X1 U45 ( .A(n43), .B(n58), .C(n24), .Y(n48) );
  XOR2X1 U46 ( .A(DE_holdout), .B(SHIFT_ENABLE_E), .Y(n43) );
  XNOR2X1 U47 ( .A(n49), .B(n53), .Y(n39) );
  NAND2X1 U49 ( .A(SHIFT_ENABLE_E), .B(n42), .Y(n49) );
  OAI21X1 U51 ( .A(n33), .B(n50), .C(n51), .Y(n46) );
  AOI21X1 U52 ( .A(n52), .B(n29), .C(state[3]), .Y(n51) );
  NOR2X1 U54 ( .A(n63), .B(n33), .Y(n52) );
  NAND2X1 U55 ( .A(n44), .B(n63), .Y(n50) );
  NAND2X1 U57 ( .A(SHIFT_ENABLE_E), .B(d_encode), .Y(n44) );
  NAND2X1 U58 ( .A(state[0]), .B(n24), .Y(n33) );
  NOR2X1 U59 ( .A(n60), .B(n59), .Y(n24) );
  NAND3X1 U62 ( .A(n59), .B(n60), .C(n58), .Y(n1) );
  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(clk), .R(n16), .S(1'b1), .Q(
        state[3]) );
  DFFSR dm_tx_out_reg ( .D(dm_tx_nxt), .CLK(clk), .R(n16), .S(1'b1), .Q(
        dm_tx_out) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n16), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n16), .S(1'b1), .Q(
        state[1]) );
  DFFSR DE_holdout_BS_reg ( .D(n64), .CLK(clk), .R(n16), .S(1'b1), .Q(
        DE_holdout_BS) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n16), .S(1'b1), .Q(
        state[2]) );
  INVX2 U29 ( .A(rst), .Y(n16) );
  INVX2 U35 ( .A(n9), .Y(n17) );
  INVX2 U39 ( .A(n12), .Y(n21) );
  INVX2 U43 ( .A(n32), .Y(n25) );
  INVX2 U48 ( .A(n43), .Y(n28) );
  INVX2 U50 ( .A(n44), .Y(n29) );
  INVX2 U53 ( .A(EOP), .Y(n30) );
  INVX2 U56 ( .A(n26), .Y(n31) );
  INVX2 U60 ( .A(n23), .Y(n34) );
  INVX2 U61 ( .A(n15), .Y(n35) );
  INVX2 U63 ( .A(d_encode), .Y(n42) );
  INVX2 U64 ( .A(DE_holdout), .Y(n53) );
  INVX2 U65 ( .A(DE_holdout_last), .Y(n54) );
  INVX2 U66 ( .A(state[3]), .Y(n56) );
  INVX2 U68 ( .A(n1), .Y(n57) );
  INVX2 U69 ( .A(state[0]), .Y(n58) );
  INVX2 U70 ( .A(state[1]), .Y(n59) );
  INVX2 U71 ( .A(state[2]), .Y(n60) );
  INVX2 U72 ( .A(DE_holdout_BS), .Y(n63) );
endmodule


module tx_shiftreg_1 ( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe, 
        send_data, d_encode );
  input [7:0] send_data;
  input clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe;
  output d_encode;
  wire   n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n11, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n54;
  wire   [7:1] present_val;
  wire   [2:0] count;

  DFFSR \count_reg[0]  ( .D(n53), .CLK(clk), .R(1'b1), .S(n14), .Q(count[0])
         );
  DFFSR \count_reg[1]  ( .D(n51), .CLK(clk), .R(1'b1), .S(n14), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n52), .CLK(clk), .R(1'b1), .S(n14), .Q(count[2])
         );
  OAI21X1 U30 ( .A(n13), .B(n54), .C(n29), .Y(n43) );
  AOI22X1 U31 ( .A(send_data[0]), .B(n17), .C(present_val[1]), .D(n15), .Y(n29) );
  OAI21X1 U32 ( .A(n13), .B(n21), .C(n30), .Y(n44) );
  NAND2X1 U33 ( .A(send_data[7]), .B(n17), .Y(n30) );
  OAI21X1 U34 ( .A(n13), .B(n22), .C(n31), .Y(n45) );
  AOI22X1 U35 ( .A(send_data[6]), .B(n17), .C(present_val[7]), .D(n15), .Y(n31) );
  OAI21X1 U36 ( .A(n13), .B(n23), .C(n32), .Y(n46) );
  AOI22X1 U37 ( .A(send_data[5]), .B(n17), .C(present_val[6]), .D(n15), .Y(n32) );
  OAI21X1 U38 ( .A(n13), .B(n24), .C(n33), .Y(n47) );
  AOI22X1 U39 ( .A(send_data[4]), .B(n17), .C(present_val[5]), .D(n15), .Y(n33) );
  OAI21X1 U40 ( .A(n13), .B(n25), .C(n34), .Y(n48) );
  AOI22X1 U41 ( .A(send_data[3]), .B(n17), .C(present_val[4]), .D(n15), .Y(n34) );
  OAI21X1 U42 ( .A(n13), .B(n26), .C(n35), .Y(n49) );
  AOI22X1 U43 ( .A(send_data[2]), .B(n17), .C(present_val[3]), .D(n15), .Y(n35) );
  OAI21X1 U44 ( .A(n27), .B(n13), .C(n36), .Y(n50) );
  AOI22X1 U45 ( .A(send_data[1]), .B(n17), .C(present_val[2]), .D(n15), .Y(n36) );
  OAI21X1 U46 ( .A(n37), .B(n38), .C(n39), .Y(n51) );
  OAI21X1 U47 ( .A(n18), .B(n11), .C(count[1]), .Y(n39) );
  NAND2X1 U48 ( .A(count[0]), .B(n19), .Y(n38) );
  OAI21X1 U49 ( .A(n17), .B(n20), .C(n40), .Y(n52) );
  NAND3X1 U50 ( .A(count[1]), .B(count[0]), .C(n15), .Y(n40) );
  OAI22X1 U51 ( .A(n18), .B(n13), .C(count[0]), .D(n37), .Y(n53) );
  NAND2X1 U52 ( .A(n13), .B(n41), .Y(n37) );
  OAI21X1 U53 ( .A(t_bitstuff), .B(n16), .C(n41), .Y(n28) );
  NAND3X1 U54 ( .A(SHIFT_ENABLE_R), .B(count[0]), .C(n42), .Y(n41) );
  NOR2X1 U55 ( .A(n19), .B(n20), .Y(n42) );
  DFFSR \present_val_reg[7]  ( .D(n44), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[7]) );
  DFFSR \present_val_reg[1]  ( .D(n50), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[1]) );
  DFFSR \present_val_reg[6]  ( .D(n45), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[6]) );
  DFFSR \present_val_reg[5]  ( .D(n46), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[5]) );
  DFFSR \present_val_reg[4]  ( .D(n47), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[4]) );
  DFFSR \present_val_reg[3]  ( .D(n48), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[3]) );
  DFFSR \present_val_reg[2]  ( .D(n49), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[2]) );
  DFFSR \present_val_reg[0]  ( .D(n43), .CLK(clk), .R(n14), .S(1'b1), .Q(
        d_encode) );
  INVX4 U3 ( .A(n11), .Y(n13) );
  INVX2 U15 ( .A(rst), .Y(n14) );
  INVX2 U16 ( .A(n41), .Y(n17) );
  INVX2 U17 ( .A(n28), .Y(n11) );
  INVX2 U18 ( .A(n37), .Y(n15) );
  INVX2 U19 ( .A(SHIFT_ENABLE_R), .Y(n16) );
  INVX2 U20 ( .A(count[0]), .Y(n18) );
  INVX2 U21 ( .A(count[1]), .Y(n19) );
  INVX2 U22 ( .A(count[2]), .Y(n20) );
  INVX2 U23 ( .A(present_val[7]), .Y(n21) );
  INVX2 U24 ( .A(present_val[6]), .Y(n22) );
  INVX2 U25 ( .A(present_val[5]), .Y(n23) );
  INVX2 U26 ( .A(present_val[4]), .Y(n24) );
  INVX2 U27 ( .A(present_val[3]), .Y(n25) );
  INVX2 U28 ( .A(present_val[2]), .Y(n26) );
  INVX2 U29 ( .A(present_val[1]), .Y(n27) );
  INVX2 U56 ( .A(d_encode), .Y(n54) );
endmodule


module tx_tcu_1_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module tx_tcu_1 ( clk, rst, p_ready, t_bitstuff, PRGA_OUT, prga_opcode, t_crc, 
        sending, EOP, next_byte, send_data, t_strobe );
  input [7:0] PRGA_OUT;
  input [1:0] prga_opcode;
  input [15:0] t_crc;
  output [7:0] send_data;
  input clk, rst, p_ready, t_bitstuff;
  output sending, EOP, next_byte, t_strobe;
  wire   N59, N60, N61, N62, N63, N64, N65, N84, N85, N86, N87, N88, N89, N90,
         N188, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n194, n195, n196, n197, n198,
         n199, n200, \r81/carry[6] , \r81/carry[5] , \r81/carry[4] ,
         \r81/carry[3] , \r81/carry[2] , \r81/carry[1] , \r81/B[0] , n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n174, n175;
  wire   [2:0] state;
  wire   [6:0] count;
  wire   [2:0] nextstate;
  wire   [7:0] flop_data;
  wire   [7:0] current_send_data;

  DFFPOSX1 \flop_data_reg[7]  ( .D(n152), .CLK(clk), .Q(flop_data[7]) );
  DFFPOSX1 \current_send_data_reg[7]  ( .D(n173), .CLK(clk), .Q(
        current_send_data[7]) );
  DFFPOSX1 \flop_data_reg[6]  ( .D(n153), .CLK(clk), .Q(flop_data[6]) );
  DFFPOSX1 \current_send_data_reg[6]  ( .D(n172), .CLK(clk), .Q(
        current_send_data[6]) );
  DFFPOSX1 \flop_data_reg[5]  ( .D(n154), .CLK(clk), .Q(flop_data[5]) );
  DFFPOSX1 \current_send_data_reg[5]  ( .D(n171), .CLK(clk), .Q(
        current_send_data[5]) );
  DFFPOSX1 \flop_data_reg[4]  ( .D(n155), .CLK(clk), .Q(flop_data[4]) );
  DFFPOSX1 \current_send_data_reg[4]  ( .D(n170), .CLK(clk), .Q(
        current_send_data[4]) );
  DFFPOSX1 \flop_data_reg[3]  ( .D(n156), .CLK(clk), .Q(flop_data[3]) );
  DFFPOSX1 \current_send_data_reg[3]  ( .D(n169), .CLK(clk), .Q(
        current_send_data[3]) );
  DFFPOSX1 \flop_data_reg[2]  ( .D(n157), .CLK(clk), .Q(flop_data[2]) );
  DFFPOSX1 \current_send_data_reg[2]  ( .D(n168), .CLK(clk), .Q(
        current_send_data[2]) );
  DFFPOSX1 \flop_data_reg[1]  ( .D(n174), .CLK(clk), .Q(flop_data[1]) );
  DFFPOSX1 \current_send_data_reg[1]  ( .D(n167), .CLK(clk), .Q(
        current_send_data[1]) );
  DFFPOSX1 \flop_data_reg[0]  ( .D(n175), .CLK(clk), .Q(flop_data[0]) );
  DFFPOSX1 \current_send_data_reg[0]  ( .D(n166), .CLK(clk), .Q(
        current_send_data[0]) );
  DFFPOSX1 \send_data_reg[7]  ( .D(n165), .CLK(clk), .Q(send_data[7]) );
  DFFPOSX1 \send_data_reg[6]  ( .D(n164), .CLK(clk), .Q(send_data[6]) );
  DFFPOSX1 \send_data_reg[5]  ( .D(n163), .CLK(clk), .Q(send_data[5]) );
  DFFPOSX1 \send_data_reg[4]  ( .D(n162), .CLK(clk), .Q(send_data[4]) );
  DFFPOSX1 \send_data_reg[3]  ( .D(n161), .CLK(clk), .Q(send_data[3]) );
  DFFPOSX1 \send_data_reg[2]  ( .D(n160), .CLK(clk), .Q(send_data[2]) );
  DFFPOSX1 \send_data_reg[1]  ( .D(n159), .CLK(clk), .Q(send_data[1]) );
  DFFPOSX1 \send_data_reg[0]  ( .D(n158), .CLK(clk), .Q(send_data[0]) );
  tx_tcu_1_DW01_inc_0 r80 ( .A({N188, count[5:0]}), .SUM({N65, N64, N63, N62, 
        N61, N60, N59}) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n15), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n15), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n15), .S(1'b1), .Q(
        state[0]) );
  DFFSR \count_reg[3]  ( .D(n196), .CLK(clk), .R(n15), .S(1'b1), .Q(count[3])
         );
  DFFSR \count_reg[2]  ( .D(n195), .CLK(clk), .R(n15), .S(1'b1), .Q(count[2])
         );
  DFFSR \count_reg[1]  ( .D(n194), .CLK(clk), .R(n15), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[0]  ( .D(n200), .CLK(clk), .R(n15), .S(1'b1), .Q(count[0])
         );
  DFFSR \count_reg[4]  ( .D(n197), .CLK(clk), .R(n15), .S(1'b1), .Q(count[4])
         );
  DFFSR \count_reg[5]  ( .D(n198), .CLK(clk), .R(n15), .S(1'b1), .Q(count[5])
         );
  DFFSR \count_reg[6]  ( .D(n199), .CLK(clk), .R(n15), .S(1'b1), .Q(N188) );
  INVX2 U13 ( .A(n12), .Y(n15) );
  BUFX2 U14 ( .A(rst), .Y(n13) );
  BUFX2 U15 ( .A(rst), .Y(n12) );
  BUFX2 U16 ( .A(rst), .Y(n14) );
  INVX2 U17 ( .A(N188), .Y(n11) );
  XOR2X1 U18 ( .A(N188), .B(\r81/carry[6] ), .Y(N90) );
  AND2X1 U19 ( .A(count[5]), .B(\r81/carry[5] ), .Y(\r81/carry[6] ) );
  XOR2X1 U20 ( .A(\r81/carry[5] ), .B(count[5]), .Y(N89) );
  AND2X1 U21 ( .A(count[4]), .B(\r81/carry[4] ), .Y(\r81/carry[5] ) );
  XOR2X1 U22 ( .A(\r81/carry[4] ), .B(count[4]), .Y(N88) );
  AND2X1 U23 ( .A(count[3]), .B(\r81/carry[3] ), .Y(\r81/carry[4] ) );
  XOR2X1 U24 ( .A(\r81/carry[3] ), .B(count[3]), .Y(N87) );
  AND2X1 U25 ( .A(count[2]), .B(\r81/carry[2] ), .Y(\r81/carry[3] ) );
  XOR2X1 U26 ( .A(\r81/carry[2] ), .B(count[2]), .Y(N86) );
  AND2X1 U27 ( .A(count[1]), .B(\r81/carry[1] ), .Y(\r81/carry[2] ) );
  XOR2X1 U28 ( .A(\r81/carry[1] ), .B(count[1]), .Y(N85) );
  AND2X1 U29 ( .A(count[0]), .B(\r81/B[0] ), .Y(\r81/carry[1] ) );
  XOR2X1 U30 ( .A(\r81/B[0] ), .B(count[0]), .Y(N84) );
  NOR2X1 U31 ( .A(n16), .B(n17), .Y(t_strobe) );
  NAND2X1 U32 ( .A(n18), .B(n19), .Y(n17) );
  NAND2X1 U33 ( .A(n11), .B(n20), .Y(n16) );
  OR2X1 U34 ( .A(n21), .B(n22), .Y(sending) );
  OAI21X1 U35 ( .A(N188), .B(n23), .C(n24), .Y(n22) );
  NAND3X1 U36 ( .A(n25), .B(n26), .C(n27), .Y(n21) );
  NAND3X1 U37 ( .A(n28), .B(n27), .C(n29), .Y(nextstate[2]) );
  AOI22X1 U38 ( .A(n30), .B(p_ready), .C(n31), .D(n32), .Y(n29) );
  NOR2X1 U39 ( .A(state[1]), .B(state[0]), .Y(n30) );
  NAND3X1 U40 ( .A(n33), .B(n34), .C(n35), .Y(nextstate[1]) );
  AOI22X1 U41 ( .A(n36), .B(n18), .C(n31), .D(n37), .Y(n35) );
  INVX1 U42 ( .A(n38), .Y(n36) );
  NAND3X1 U43 ( .A(n39), .B(n40), .C(p_ready), .Y(n33) );
  NAND3X1 U44 ( .A(n41), .B(n28), .C(n42), .Y(nextstate[0]) );
  AOI21X1 U45 ( .A(n18), .B(n38), .C(n43), .Y(n42) );
  OAI21X1 U46 ( .A(n44), .B(n27), .C(n45), .Y(n43) );
  NAND3X1 U47 ( .A(p_ready), .B(n37), .C(n31), .Y(n45) );
  AND2X1 U48 ( .A(n46), .B(n47), .Y(n31) );
  INVX1 U49 ( .A(n48), .Y(n44) );
  NAND3X1 U50 ( .A(n19), .B(n11), .C(count[0]), .Y(n38) );
  INVX1 U51 ( .A(n49), .Y(n28) );
  AND2X1 U52 ( .A(n26), .B(n25), .Y(n41) );
  OAI21X1 U53 ( .A(n50), .B(n51), .C(n52), .Y(next_byte) );
  MUX2X1 U54 ( .B(n53), .A(n54), .S(n55), .Y(n152) );
  INVX1 U55 ( .A(n56), .Y(n153) );
  MUX2X1 U56 ( .B(PRGA_OUT[6]), .A(flop_data[6]), .S(n55), .Y(n56) );
  INVX1 U57 ( .A(n57), .Y(n154) );
  MUX2X1 U58 ( .B(PRGA_OUT[5]), .A(flop_data[5]), .S(n55), .Y(n57) );
  INVX1 U59 ( .A(n58), .Y(n155) );
  MUX2X1 U60 ( .B(PRGA_OUT[4]), .A(flop_data[4]), .S(n55), .Y(n58) );
  INVX1 U61 ( .A(n59), .Y(n156) );
  MUX2X1 U62 ( .B(PRGA_OUT[3]), .A(flop_data[3]), .S(n55), .Y(n59) );
  INVX1 U63 ( .A(n60), .Y(n157) );
  MUX2X1 U64 ( .B(PRGA_OUT[2]), .A(flop_data[2]), .S(n55), .Y(n60) );
  INVX1 U65 ( .A(n61), .Y(n174) );
  MUX2X1 U66 ( .B(PRGA_OUT[1]), .A(flop_data[1]), .S(n55), .Y(n61) );
  INVX1 U67 ( .A(n62), .Y(n175) );
  MUX2X1 U68 ( .B(PRGA_OUT[0]), .A(flop_data[0]), .S(n55), .Y(n62) );
  NAND3X1 U69 ( .A(n63), .B(n23), .C(n64), .Y(n55) );
  AND2X1 U70 ( .A(n24), .B(n52), .Y(n64) );
  MUX2X1 U71 ( .B(n65), .A(n66), .S(n40), .Y(n52) );
  NOR2X1 U72 ( .A(p_ready), .B(n67), .Y(n66) );
  NOR2X1 U73 ( .A(n14), .B(n65), .Y(n63) );
  INVX1 U74 ( .A(t_bitstuff), .Y(\r81/B[0] ) );
  OAI21X1 U75 ( .A(n20), .B(n68), .C(n69), .Y(n200) );
  AOI22X1 U76 ( .A(N59), .B(n70), .C(N84), .D(n71), .Y(n69) );
  OAI21X1 U77 ( .A(n11), .B(n68), .C(n72), .Y(n199) );
  AOI22X1 U78 ( .A(N65), .B(n70), .C(N90), .D(n71), .Y(n72) );
  OAI21X1 U79 ( .A(n73), .B(n68), .C(n74), .Y(n198) );
  AOI22X1 U80 ( .A(N64), .B(n70), .C(N89), .D(n71), .Y(n74) );
  OAI21X1 U81 ( .A(n75), .B(n68), .C(n76), .Y(n197) );
  AOI22X1 U82 ( .A(N63), .B(n70), .C(N88), .D(n71), .Y(n76) );
  OAI21X1 U83 ( .A(n77), .B(n68), .C(n78), .Y(n196) );
  AOI22X1 U84 ( .A(N62), .B(n70), .C(N87), .D(n71), .Y(n78) );
  OAI21X1 U85 ( .A(n79), .B(n68), .C(n80), .Y(n195) );
  AOI22X1 U86 ( .A(N61), .B(n70), .C(N86), .D(n71), .Y(n80) );
  OAI21X1 U87 ( .A(n81), .B(n68), .C(n82), .Y(n194) );
  AOI22X1 U88 ( .A(N60), .B(n70), .C(N85), .D(n71), .Y(n82) );
  OAI21X1 U89 ( .A(n32), .B(n51), .C(n34), .Y(n71) );
  OR2X1 U90 ( .A(n25), .B(n48), .Y(n34) );
  NAND3X1 U91 ( .A(state[0]), .B(n83), .C(state[1]), .Y(n25) );
  INVX1 U92 ( .A(n37), .Y(n32) );
  NAND2X1 U93 ( .A(n48), .B(n50), .Y(n37) );
  AND2X1 U94 ( .A(prga_opcode[1]), .B(prga_opcode[0]), .Y(n50) );
  AND2X1 U95 ( .A(n68), .B(n84), .Y(n70) );
  OAI21X1 U96 ( .A(n48), .B(n27), .C(n85), .Y(n84) );
  NOR2X1 U97 ( .A(n18), .B(n49), .Y(n85) );
  NOR2X1 U98 ( .A(n86), .B(n87), .Y(n48) );
  NAND3X1 U99 ( .A(count[4]), .B(count[1]), .C(count[5]), .Y(n87) );
  NAND3X1 U100 ( .A(count[0]), .B(count[3]), .C(n88), .Y(n86) );
  NOR2X1 U101 ( .A(N188), .B(n79), .Y(n88) );
  NAND2X1 U102 ( .A(n18), .B(t_bitstuff), .Y(n68) );
  INVX1 U103 ( .A(count[1]), .Y(n81) );
  OAI21X1 U104 ( .A(n89), .B(n90), .C(n91), .Y(n173) );
  INVX1 U105 ( .A(current_send_data[7]), .Y(n90) );
  OAI21X1 U106 ( .A(n89), .B(n92), .C(n93), .Y(n172) );
  INVX1 U107 ( .A(current_send_data[6]), .Y(n92) );
  OAI21X1 U108 ( .A(n89), .B(n94), .C(n95), .Y(n171) );
  INVX1 U109 ( .A(current_send_data[5]), .Y(n94) );
  OAI21X1 U110 ( .A(n89), .B(n96), .C(n97), .Y(n170) );
  INVX1 U111 ( .A(current_send_data[4]), .Y(n96) );
  OAI21X1 U112 ( .A(n89), .B(n98), .C(n99), .Y(n169) );
  INVX1 U113 ( .A(current_send_data[3]), .Y(n98) );
  OAI21X1 U114 ( .A(n89), .B(n100), .C(n101), .Y(n168) );
  INVX1 U115 ( .A(current_send_data[2]), .Y(n100) );
  OAI21X1 U116 ( .A(n89), .B(n102), .C(n103), .Y(n167) );
  INVX1 U117 ( .A(current_send_data[1]), .Y(n102) );
  OAI21X1 U118 ( .A(n89), .B(n104), .C(n105), .Y(n166) );
  INVX1 U119 ( .A(current_send_data[0]), .Y(n104) );
  AOI21X1 U120 ( .A(state[0]), .B(state[1]), .C(n13), .Y(n89) );
  NAND2X1 U121 ( .A(n106), .B(n91), .Y(n165) );
  NOR2X1 U122 ( .A(n107), .B(n108), .Y(n91) );
  OAI21X1 U123 ( .A(n53), .B(n109), .C(n110), .Y(n108) );
  NAND2X1 U124 ( .A(t_crc[15]), .B(n111), .Y(n110) );
  INVX1 U125 ( .A(n112), .Y(n109) );
  INVX1 U126 ( .A(PRGA_OUT[7]), .Y(n53) );
  OAI22X1 U127 ( .A(n54), .B(n113), .C(n114), .D(n115), .Y(n107) );
  NAND2X1 U128 ( .A(n116), .B(state[0]), .Y(n115) );
  OAI21X1 U129 ( .A(N188), .B(t_crc[7]), .C(n15), .Y(n114) );
  INVX1 U130 ( .A(n117), .Y(n113) );
  INVX1 U131 ( .A(flop_data[7]), .Y(n54) );
  AOI22X1 U132 ( .A(n118), .B(current_send_data[7]), .C(send_data[7]), .D(n12), 
        .Y(n106) );
  NAND2X1 U133 ( .A(n119), .B(n93), .Y(n164) );
  AND2X1 U134 ( .A(n120), .B(n121), .Y(n93) );
  AOI22X1 U135 ( .A(t_crc[6]), .B(n122), .C(n117), .D(flop_data[6]), .Y(n121)
         );
  AOI22X1 U136 ( .A(t_crc[14]), .B(n111), .C(n112), .D(PRGA_OUT[6]), .Y(n120)
         );
  AOI22X1 U137 ( .A(n118), .B(current_send_data[6]), .C(send_data[6]), .D(n12), 
        .Y(n119) );
  NAND2X1 U138 ( .A(n123), .B(n95), .Y(n163) );
  AND2X1 U139 ( .A(n124), .B(n125), .Y(n95) );
  AOI22X1 U140 ( .A(t_crc[5]), .B(n122), .C(n117), .D(flop_data[5]), .Y(n125)
         );
  AOI22X1 U141 ( .A(t_crc[13]), .B(n111), .C(n112), .D(PRGA_OUT[5]), .Y(n124)
         );
  AOI22X1 U142 ( .A(n118), .B(current_send_data[5]), .C(send_data[5]), .D(n13), 
        .Y(n123) );
  NAND2X1 U143 ( .A(n126), .B(n97), .Y(n162) );
  AND2X1 U144 ( .A(n127), .B(n128), .Y(n97) );
  AOI22X1 U145 ( .A(t_crc[4]), .B(n122), .C(n117), .D(flop_data[4]), .Y(n128)
         );
  AOI22X1 U146 ( .A(t_crc[12]), .B(n111), .C(n112), .D(PRGA_OUT[4]), .Y(n127)
         );
  AOI22X1 U147 ( .A(n118), .B(current_send_data[4]), .C(send_data[4]), .D(n13), 
        .Y(n126) );
  NAND2X1 U148 ( .A(n129), .B(n99), .Y(n161) );
  AND2X1 U149 ( .A(n130), .B(n131), .Y(n99) );
  AOI22X1 U150 ( .A(t_crc[3]), .B(n122), .C(n117), .D(flop_data[3]), .Y(n131)
         );
  AOI22X1 U151 ( .A(t_crc[11]), .B(n111), .C(n112), .D(PRGA_OUT[3]), .Y(n130)
         );
  AOI22X1 U152 ( .A(n118), .B(current_send_data[3]), .C(send_data[3]), .D(n13), 
        .Y(n129) );
  NAND2X1 U153 ( .A(n132), .B(n101), .Y(n160) );
  AND2X1 U154 ( .A(n133), .B(n134), .Y(n101) );
  AOI22X1 U155 ( .A(t_crc[2]), .B(n122), .C(n117), .D(flop_data[2]), .Y(n134)
         );
  AOI22X1 U156 ( .A(t_crc[10]), .B(n111), .C(n112), .D(PRGA_OUT[2]), .Y(n133)
         );
  AOI22X1 U157 ( .A(n118), .B(current_send_data[2]), .C(send_data[2]), .D(n13), 
        .Y(n132) );
  NAND2X1 U158 ( .A(n135), .B(n103), .Y(n159) );
  AND2X1 U159 ( .A(n136), .B(n137), .Y(n103) );
  AOI22X1 U160 ( .A(t_crc[1]), .B(n122), .C(n117), .D(flop_data[1]), .Y(n137)
         );
  AOI22X1 U161 ( .A(t_crc[9]), .B(n111), .C(n112), .D(PRGA_OUT[1]), .Y(n136)
         );
  AOI22X1 U162 ( .A(n118), .B(current_send_data[1]), .C(send_data[1]), .D(n13), 
        .Y(n135) );
  NAND2X1 U163 ( .A(n138), .B(n105), .Y(n158) );
  AND2X1 U164 ( .A(n139), .B(n140), .Y(n105) );
  AOI22X1 U165 ( .A(t_crc[0]), .B(n122), .C(n117), .D(flop_data[0]), .Y(n140)
         );
  NOR2X1 U166 ( .A(n24), .B(n13), .Y(n117) );
  NOR2X1 U167 ( .A(n46), .B(n18), .Y(n24) );
  NOR2X1 U168 ( .A(n40), .B(n67), .Y(n18) );
  INVX1 U169 ( .A(n39), .Y(n67) );
  NOR2X1 U170 ( .A(state[1]), .B(state[2]), .Y(n39) );
  INVX1 U171 ( .A(n51), .Y(n46) );
  INVX1 U172 ( .A(n141), .Y(n122) );
  NAND3X1 U173 ( .A(n116), .B(state[0]), .C(n142), .Y(n141) );
  NOR2X1 U174 ( .A(n14), .B(N188), .Y(n142) );
  AOI22X1 U175 ( .A(t_crc[8]), .B(n111), .C(n112), .D(PRGA_OUT[0]), .Y(n139)
         );
  NOR2X1 U176 ( .A(n26), .B(n13), .Y(n112) );
  NAND2X1 U177 ( .A(n65), .B(n40), .Y(n26) );
  NOR2X1 U178 ( .A(n83), .B(n143), .Y(n65) );
  INVX1 U179 ( .A(state[1]), .Y(n143) );
  NOR2X1 U180 ( .A(n27), .B(n14), .Y(n111) );
  NAND2X1 U181 ( .A(n116), .B(n40), .Y(n27) );
  AOI22X1 U182 ( .A(n118), .B(current_send_data[0]), .C(send_data[0]), .D(n12), 
        .Y(n138) );
  INVX1 U183 ( .A(n144), .Y(n118) );
  NAND3X1 U184 ( .A(state[0]), .B(n15), .C(state[1]), .Y(n144) );
  OAI21X1 U185 ( .A(n51), .B(n47), .C(n145), .Y(EOP) );
  NAND3X1 U186 ( .A(N188), .B(n146), .C(n49), .Y(n145) );
  NOR2X1 U187 ( .A(n23), .B(n147), .Y(n49) );
  OAI21X1 U188 ( .A(n148), .B(n149), .C(state[0]), .Y(n147) );
  NAND3X1 U189 ( .A(count[2]), .B(N188), .C(count[3]), .Y(n149) );
  NAND3X1 U190 ( .A(n75), .B(n73), .C(n150), .Y(n148) );
  NOR2X1 U191 ( .A(count[1]), .B(count[0]), .Y(n150) );
  INVX1 U192 ( .A(count[5]), .Y(n73) );
  INVX1 U193 ( .A(count[4]), .Y(n75) );
  INVX1 U194 ( .A(n116), .Y(n23) );
  NOR2X1 U195 ( .A(n83), .B(state[1]), .Y(n116) );
  NAND3X1 U196 ( .A(n19), .B(n20), .C(N188), .Y(n47) );
  INVX1 U197 ( .A(count[0]), .Y(n20) );
  NOR2X1 U198 ( .A(n146), .B(count[1]), .Y(n19) );
  NAND3X1 U199 ( .A(n79), .B(n77), .C(n151), .Y(n146) );
  NOR2X1 U200 ( .A(count[5]), .B(count[4]), .Y(n151) );
  INVX1 U201 ( .A(count[3]), .Y(n77) );
  INVX1 U202 ( .A(count[2]), .Y(n79) );
  NAND3X1 U203 ( .A(n40), .B(n83), .C(state[1]), .Y(n51) );
  INVX1 U204 ( .A(state[2]), .Y(n83) );
  INVX1 U205 ( .A(state[0]), .Y(n40) );
endmodule


module tx_timer_1 ( CLK, RST, SENDING, SHIFT_ENABLE_R, SHIFT_ENABLE_E );
  input CLK, RST, SENDING;
  output SHIFT_ENABLE_R, SHIFT_ENABLE_E;
  wire   state, nxt_SHIFT_ENABLE_E, n12, n13, n14, n15, n16, n17, n18, n19, n7,
         n8, n9, n10, n11;
  wire   [3:0] count;
  wire   [3:0] nextcount;
  assign SHIFT_ENABLE_R = nxt_SHIFT_ENABLE_E;

  NOR2X1 U14 ( .A(n12), .B(n13), .Y(nextcount[3]) );
  XNOR2X1 U15 ( .A(count[3]), .B(n14), .Y(n12) );
  NOR2X1 U16 ( .A(n15), .B(n9), .Y(n14) );
  AOI21X1 U17 ( .A(n16), .B(state), .C(n11), .Y(nextcount[2]) );
  XNOR2X1 U18 ( .A(n15), .B(n9), .Y(n16) );
  NAND2X1 U19 ( .A(count[1]), .B(count[0]), .Y(n15) );
  NOR2X1 U20 ( .A(n17), .B(n13), .Y(nextcount[1]) );
  NAND3X1 U21 ( .A(SENDING), .B(n18), .C(state), .Y(n13) );
  XNOR2X1 U22 ( .A(count[0]), .B(count[1]), .Y(n17) );
  OAI21X1 U23 ( .A(count[0]), .B(n11), .C(state), .Y(nextcount[0]) );
  NOR2X1 U24 ( .A(n18), .B(n19), .Y(nxt_SHIFT_ENABLE_E) );
  NAND3X1 U25 ( .A(count[3]), .B(SENDING), .C(state), .Y(n19) );
  NAND3X1 U26 ( .A(n10), .B(n9), .C(n8), .Y(n18) );
  DFFSR state_reg ( .D(SENDING), .CLK(CLK), .R(n7), .S(1'b1), .Q(state) );
  DFFSR \count_reg[2]  ( .D(nextcount[2]), .CLK(CLK), .R(n7), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[0]  ( .D(nextcount[0]), .CLK(CLK), .R(n7), .S(1'b1), .Q(
        count[0]) );
  DFFSR \count_reg[3]  ( .D(nextcount[3]), .CLK(CLK), .R(n7), .S(1'b1), .Q(
        count[3]) );
  DFFSR \count_reg[1]  ( .D(nextcount[1]), .CLK(CLK), .R(n7), .S(1'b1), .Q(
        count[1]) );
  DFFSR SHIFT_ENABLE_E_reg ( .D(nxt_SHIFT_ENABLE_E), .CLK(CLK), .R(n7), .S(
        1'b1), .Q(SHIFT_ENABLE_E) );
  INVX2 U9 ( .A(RST), .Y(n7) );
  INVX2 U10 ( .A(count[0]), .Y(n8) );
  INVX2 U11 ( .A(count[2]), .Y(n9) );
  INVX2 U12 ( .A(count[1]), .Y(n10) );
  INVX2 U13 ( .A(SENDING), .Y(n11) );
endmodule


module transmitter_block_1 ( PRGA_OUT, clk, p_ready, prga_opcode, rst, SENDING, 
        dm_tx_out, dp_tx_out, NEXT_BYTE );
  input [7:0] PRGA_OUT;
  input [1:0] prga_opcode;
  input clk, p_ready, rst;
  output SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE;
  wire   t_strobe, EOP, SHIFT_ENABLE_E, d_encode, t_bitstuff, SHIFT_ENABLE_R;
  wire   [15:0] TX_CRC;
  wire   [7:0] send_data;

  tx_CRC_CALC_1 U_1 ( .CLK(clk), .RST(rst), .EOP(EOP), .T_STROBE(t_strobe), 
        .PRGA_OPCODE(prga_opcode), .PRGA_OUT(PRGA_OUT), .TX_CRC(TX_CRC) );
  tx_encode_1 U_0 ( .clk(clk), .rst(rst), .SHIFT_ENABLE_E(SHIFT_ENABLE_E), 
        .d_encode(d_encode), .EOP(EOP), .t_bitstuff(t_bitstuff), .dp_tx_out(
        dp_tx_out), .dm_tx_out(dm_tx_out) );
  tx_shiftreg_1 U_2 ( .clk(clk), .rst(rst), .SHIFT_ENABLE_R(SHIFT_ENABLE_R), 
        .t_bitstuff(t_bitstuff), .t_strobe(t_strobe), .send_data(send_data), 
        .d_encode(d_encode) );
  tx_tcu_1 U_3 ( .clk(clk), .rst(rst), .p_ready(p_ready), .t_bitstuff(
        t_bitstuff), .PRGA_OUT(PRGA_OUT), .prga_opcode(prga_opcode), .t_crc(
        TX_CRC), .sending(SENDING), .EOP(EOP), .next_byte(NEXT_BYTE), 
        .send_data(send_data), .t_strobe(t_strobe) );
  tx_timer_1 U_4 ( .CLK(clk), .RST(rst), .SENDING(SENDING), .SHIFT_ENABLE_R(
        SHIFT_ENABLE_R), .SHIFT_ENABLE_E(SHIFT_ENABLE_E) );
endmodule


module RMEDT_REWIRE_1 ( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN, DATA_IN, BS_ERROR, 
        CRC_ERROR, EMPTY, FULL, KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, 
        R_ERROR, SENDING, dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE, DATA, 
        ADDR );
  input [7:0] DATA_IN;
  output [7:0] DATA;
  output [7:0] ADDR;
  input CLK, DM1_RX, DP1_RX, RST, SERIAL_IN;
  output BS_ERROR, CRC_ERROR, EMPTY, FULL, KEY_ERROR, PROG_ERROR, PARITY_ERROR,
         RBUF_FULL, R_ERROR, SENDING, dm_tx_out, dp_tx_out, W_ENABLE_R,
         R_ENABLE;
  wire   B_READY, PDATA_READY, EOP_external, NEXT_BYTE, W_ENABLE, n1, n2;
  wire   [7:0] PRGA_IN;
  wire   [1:0] PRGA_OPCODE;
  wire   [7:0] PROCESSED_DATA;
  wire   [7:0] RCV_DATA;
  wire   [1:0] OPCODE;

  EDBlock_1 U_0 ( .BYTE(PRGA_IN), .BYTE_READY(B_READY), .CLK(CLK), .OPCODE(
        PRGA_OPCODE), .RST(n1), .SERIAL_IN(SERIAL_IN), .DATA_IN(DATA_IN), 
        .KEY_ERROR(KEY_ERROR), .PARITY_ERROR(PARITY_ERROR), .PDATA_READY(
        PDATA_READY), .PROCESSED_DATA(PROCESSED_DATA), .PROG_ERROR(PROG_ERROR), 
        .RBUF_FULL(RBUF_FULL), .W_ENABLE(W_ENABLE_R), .R_ENABLE(R_ENABLE), 
        .DATA(DATA), .ADDR(ADDR) );
  memoryblock_1 U_1 ( .CLK(CLK), .NEXT_BYTE(NEXT_BYTE), .RCV_DATA(RCV_DATA), 
        .RCV_OPCODE(OPCODE), .RST(n1), .W_ENABLE(W_ENABLE), .EOP(EOP_external), 
        .EMPTY(EMPTY), .FULL(FULL), .B_READY(B_READY), .PRGA_IN(PRGA_IN), 
        .PRGA_OPCODE(PRGA_OPCODE) );
  receiver_block_rewire_1 U_2 ( .CLK(CLK), .DM1_RX(DM1_RX), .DP1_RX(DP1_RX), 
        .RST(n1), .BS_ERROR(BS_ERROR), .CRC_ERROR(CRC_ERROR), .EOP_external(
        EOP_external), .OPCODE(OPCODE), .RCV_DATA(RCV_DATA), .R_ERROR(R_ERROR), 
        .W_ENABLE(W_ENABLE) );
  transmitter_block_1 U_3 ( .PRGA_OUT(PROCESSED_DATA), .clk(CLK), .p_ready(
        PDATA_READY), .prga_opcode(PRGA_OPCODE), .rst(n1), .SENDING(SENDING), 
        .dm_tx_out(dm_tx_out), .dp_tx_out(dp_tx_out), .NEXT_BYTE(NEXT_BYTE) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module KSA_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module KSA_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module KSA_0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_0_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module KSA_0_DW01_add_3 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [7:1] carry;

  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n6), .YC(carry[2]), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(carry[4]), .B(n1), .Y(SUM[4]) );
  NAND2X1 U3 ( .A(carry[4]), .B(B[4]), .Y(n2) );
  NAND2X1 U4 ( .A(carry[4]), .B(A[4]), .Y(n3) );
  NAND2X1 U5 ( .A(B[4]), .B(A[4]), .Y(n4) );
  NAND3X1 U6 ( .A(n3), .B(n2), .C(n4), .Y(carry[5]) );
  XOR2X1 U7 ( .A(B[7]), .B(A[7]), .Y(n5) );
  XOR2X1 U8 ( .A(carry[7]), .B(n5), .Y(SUM[7]) );
  AND2X2 U9 ( .A(B[0]), .B(A[0]), .Y(n6) );
  XOR2X1 U10 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module KSA_0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(A[5]), .B(n10), .Y(n2) );
  XOR2X1 U3 ( .A(n2), .B(carry[5]), .Y(SUM[5]) );
  NAND2X1 U4 ( .A(A[5]), .B(n10), .Y(n3) );
  NAND2X1 U5 ( .A(A[5]), .B(carry[5]), .Y(n4) );
  NAND2X1 U6 ( .A(n10), .B(carry[5]), .Y(n5) );
  NAND3X1 U7 ( .A(n3), .B(n4), .C(n5), .Y(carry[6]) );
  XOR2X1 U8 ( .A(A[6]), .B(n11), .Y(n6) );
  XOR2X1 U9 ( .A(n6), .B(carry[6]), .Y(SUM[6]) );
  NAND2X1 U10 ( .A(A[6]), .B(n11), .Y(n7) );
  NAND2X1 U11 ( .A(A[6]), .B(carry[6]), .Y(n8) );
  NAND2X1 U12 ( .A(n11), .B(carry[6]), .Y(n9) );
  NAND3X1 U13 ( .A(n7), .B(n8), .C(n9), .Y(carry[7]) );
  BUFX2 U14 ( .A(B[5]), .Y(n10) );
  BUFX2 U15 ( .A(B[6]), .Y(n11) );
  XOR2X1 U16 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module KSA_0 ( KEY, CLK, RST, KEY_ERROR, BYTE_READY, BYTE, OPCODE, DATA_IN, 
        PROCESSED_DATA, PDATA_READY, W_ENABLE, R_ENABLE, ADDR, DATA );
  input [63:0] KEY;
  input [7:0] BYTE;
  input [1:0] OPCODE;
  input [7:0] DATA_IN;
  output [7:0] PROCESSED_DATA;
  output [7:0] ADDR;
  output [7:0] DATA;
  input CLK, RST, KEY_ERROR, BYTE_READY;
  output PDATA_READY, W_ENABLE, R_ENABLE;
  wire   permuteComplete, \keyTable[0][7] , \keyTable[0][6] , \keyTable[0][5] ,
         \keyTable[0][4] , \keyTable[0][3] , \keyTable[0][2] ,
         \keyTable[0][1] , \keyTable[0][0] , \keyTable[1][7] ,
         \keyTable[1][6] , \keyTable[1][5] , \keyTable[1][4] ,
         \keyTable[1][3] , \keyTable[1][2] , \keyTable[1][1] ,
         \keyTable[1][0] , \keyTable[2][7] , \keyTable[2][6] ,
         \keyTable[2][5] , \keyTable[2][4] , \keyTable[2][3] ,
         \keyTable[2][2] , \keyTable[2][1] , \keyTable[2][0] ,
         \keyTable[3][7] , \keyTable[3][6] , \keyTable[3][5] ,
         \keyTable[3][4] , \keyTable[3][3] , \keyTable[3][2] ,
         \keyTable[3][1] , \keyTable[3][0] , \keyTable[4][7] ,
         \keyTable[4][6] , \keyTable[4][5] , \keyTable[4][4] ,
         \keyTable[4][3] , \keyTable[4][2] , \keyTable[4][1] ,
         \keyTable[4][0] , \keyTable[5][7] , \keyTable[5][6] ,
         \keyTable[5][5] , \keyTable[5][4] , \keyTable[5][3] ,
         \keyTable[5][2] , \keyTable[5][1] , \keyTable[5][0] ,
         \keyTable[6][7] , \keyTable[6][6] , \keyTable[6][5] ,
         \keyTable[6][4] , \keyTable[6][3] , \keyTable[6][2] ,
         \keyTable[6][1] , \keyTable[6][0] , \keyTable[7][7] ,
         \keyTable[7][6] , \keyTable[7][5] , \keyTable[7][4] ,
         \keyTable[7][3] , \keyTable[7][2] , \keyTable[7][1] ,
         \keyTable[7][0] , fw_enable, fr_enable, N407, N408, N409, N410, N411,
         N412, N413, N414, N424, N425, N426, N427, N428, N429, N430, N431,
         N442, N443, N444, N445, N446, N447, N448, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N496, N497, N498, N499, N500, N501, N502, N503, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N456, N455, N454, N453, N452, N451, N450, N449, n3,
         n4, n5, n6, n7, n8, n9, n10, n12, n14, n15, n16, n17, n20, n22, n24,
         n27, n29, n32, n34, n37, n39, n42, n44, n47, n216, n218, n220, n230,
         n235, n237, n238, n239, n240, n241, n244, n246, n247, n249, n250,
         n252, n253, n255, n256, n258, n259, n261, n262, n264, n265, n267,
         n268, n270, n271, n275, n277, n280, n282, n285, n287, n290, n292,
         n295, n297, n300, n302, n305, n307, n311, n317, n318, n326, n327,
         n329, n331, n333, n335, n337, n339, n341, n343, n345, n347, n349,
         n351, n353, n355, n357, n359, n361, n363, n365, n367, n369, n371,
         n373, n375, n377, n379, n381, n383, n385, n387, n389, n391, n393,
         n395, n397, n399, n401, n403, n405, n407, n409, n411, n413, n415,
         n417, n419, n421, n423, n425, n427, n429, n431, n433, n435, n437,
         n439, n441, n443, n445, n447, n449, n451, n453, n455, n458, n459,
         n462, n463, n465, n467, n469, n471, n473, n475, n480, n482, n488,
         n498, n500, n501, n503, n504, n505, n506, n507, n509, n512, n514,
         n516, n518, n520, n522, n524, n528, n540, n541, n542, n543, n545,
         n547, n549, n551, n553, n555, n557, n562, n569, n571, n572, n575,
         n577, n579, n581, n592, n594, n600, n604, n605, n606, n610, n612,
         n614, n616, n618, n624, n626, n629, n630, n632, n636, n637, n638,
         n648, n649, n650, n651, n692, n701, n746, n748, n750, n752, n754,
         n756, n758, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n864, n865, n866, n867, n868, n869, n870, n871, n883, n884,
         n885, n886, n887, n888, n889, n890, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602;
  wire   [4:0] state;
  wire   [7:0] si;
  wire   [7:0] sj;
  wire   [7:0] currentProcessedData;
  wire   [4:0] nextState;
  wire   [7:0] inti;
  wire   [7:0] intj;
  wire   [2:0] keyi;
  wire   [7:0] temp;
  wire   [7:0] extratemp;
  wire   [7:0] nextProcessedData;
  wire   [7:0] delaydata;
  wire   [7:0] prefillCounter;
  wire   [7:0] faddr;
  wire   [7:0] fdata;
  tri   [7:0] nfaddr;
  tri   [7:0] nfdata;

  DFFPOSX1 \prefillCounter_reg[0]  ( .D(n986), .CLK(CLK), .Q(prefillCounter[0]) );
  DFFPOSX1 permuteComplete_reg ( .D(n1002), .CLK(CLK), .Q(permuteComplete) );
  DFFPOSX1 \extratemp_reg[7]  ( .D(n482), .CLK(CLK), .Q(extratemp[7]) );
  DFFPOSX1 \extratemp_reg[6]  ( .D(n480), .CLK(CLK), .Q(extratemp[6]) );
  DFFPOSX1 \extratemp_reg[5]  ( .D(n475), .CLK(CLK), .Q(extratemp[5]) );
  DFFPOSX1 \extratemp_reg[4]  ( .D(n473), .CLK(CLK), .Q(extratemp[4]) );
  DFFPOSX1 \extratemp_reg[3]  ( .D(n471), .CLK(CLK), .Q(extratemp[3]) );
  DFFPOSX1 \extratemp_reg[2]  ( .D(n469), .CLK(CLK), .Q(extratemp[2]) );
  DFFPOSX1 \extratemp_reg[1]  ( .D(n467), .CLK(CLK), .Q(extratemp[1]) );
  DFFPOSX1 \extratemp_reg[0]  ( .D(n465), .CLK(CLK), .Q(extratemp[0]) );
  DFFPOSX1 \keyTable_reg[7][0]  ( .D(n1093), .CLK(CLK), .Q(\keyTable[7][0] )
         );
  DFFPOSX1 \keyTable_reg[7][1]  ( .D(n1092), .CLK(CLK), .Q(\keyTable[7][1] )
         );
  DFFPOSX1 \keyTable_reg[7][2]  ( .D(n1091), .CLK(CLK), .Q(\keyTable[7][2] )
         );
  DFFPOSX1 \keyTable_reg[7][3]  ( .D(n1090), .CLK(CLK), .Q(\keyTable[7][3] )
         );
  DFFPOSX1 \keyTable_reg[7][4]  ( .D(n1089), .CLK(CLK), .Q(\keyTable[7][4] )
         );
  DFFPOSX1 \keyTable_reg[7][5]  ( .D(n1088), .CLK(CLK), .Q(\keyTable[7][5] )
         );
  DFFPOSX1 \keyTable_reg[7][6]  ( .D(n1087), .CLK(CLK), .Q(\keyTable[7][6] )
         );
  DFFPOSX1 \keyTable_reg[7][7]  ( .D(n1086), .CLK(CLK), .Q(\keyTable[7][7] )
         );
  DFFPOSX1 \keyTable_reg[6][0]  ( .D(n1085), .CLK(CLK), .Q(\keyTable[6][0] )
         );
  DFFPOSX1 \keyTable_reg[6][1]  ( .D(n1084), .CLK(CLK), .Q(\keyTable[6][1] )
         );
  DFFPOSX1 \keyTable_reg[6][2]  ( .D(n1083), .CLK(CLK), .Q(\keyTable[6][2] )
         );
  DFFPOSX1 \keyTable_reg[6][3]  ( .D(n1082), .CLK(CLK), .Q(\keyTable[6][3] )
         );
  DFFPOSX1 \keyTable_reg[6][4]  ( .D(n1081), .CLK(CLK), .Q(\keyTable[6][4] )
         );
  DFFPOSX1 \keyTable_reg[6][5]  ( .D(n1080), .CLK(CLK), .Q(\keyTable[6][5] )
         );
  DFFPOSX1 \keyTable_reg[6][6]  ( .D(n1079), .CLK(CLK), .Q(\keyTable[6][6] )
         );
  DFFPOSX1 \keyTable_reg[6][7]  ( .D(n1078), .CLK(CLK), .Q(\keyTable[6][7] )
         );
  DFFPOSX1 \keyTable_reg[5][0]  ( .D(n1077), .CLK(CLK), .Q(\keyTable[5][0] )
         );
  DFFPOSX1 \keyTable_reg[5][1]  ( .D(n1076), .CLK(CLK), .Q(\keyTable[5][1] )
         );
  DFFPOSX1 \keyTable_reg[5][2]  ( .D(n1075), .CLK(CLK), .Q(\keyTable[5][2] )
         );
  DFFPOSX1 \keyTable_reg[5][3]  ( .D(n1074), .CLK(CLK), .Q(\keyTable[5][3] )
         );
  DFFPOSX1 \keyTable_reg[5][4]  ( .D(n1073), .CLK(CLK), .Q(\keyTable[5][4] )
         );
  DFFPOSX1 \keyTable_reg[5][5]  ( .D(n1072), .CLK(CLK), .Q(\keyTable[5][5] )
         );
  DFFPOSX1 \keyTable_reg[5][6]  ( .D(n1071), .CLK(CLK), .Q(\keyTable[5][6] )
         );
  DFFPOSX1 \keyTable_reg[5][7]  ( .D(n1070), .CLK(CLK), .Q(\keyTable[5][7] )
         );
  DFFPOSX1 \keyTable_reg[4][0]  ( .D(n1069), .CLK(CLK), .Q(\keyTable[4][0] )
         );
  DFFPOSX1 \keyTable_reg[4][1]  ( .D(n1068), .CLK(CLK), .Q(\keyTable[4][1] )
         );
  DFFPOSX1 \keyTable_reg[4][2]  ( .D(n1067), .CLK(CLK), .Q(\keyTable[4][2] )
         );
  DFFPOSX1 \keyTable_reg[4][3]  ( .D(n1066), .CLK(CLK), .Q(\keyTable[4][3] )
         );
  DFFPOSX1 \keyTable_reg[4][4]  ( .D(n1065), .CLK(CLK), .Q(\keyTable[4][4] )
         );
  DFFPOSX1 \keyTable_reg[4][5]  ( .D(n1064), .CLK(CLK), .Q(\keyTable[4][5] )
         );
  DFFPOSX1 \keyTable_reg[4][6]  ( .D(n1063), .CLK(CLK), .Q(\keyTable[4][6] )
         );
  DFFPOSX1 \keyTable_reg[4][7]  ( .D(n1062), .CLK(CLK), .Q(\keyTable[4][7] )
         );
  DFFPOSX1 \keyTable_reg[3][0]  ( .D(n1061), .CLK(CLK), .Q(\keyTable[3][0] )
         );
  DFFPOSX1 \keyTable_reg[3][1]  ( .D(n1060), .CLK(CLK), .Q(\keyTable[3][1] )
         );
  DFFPOSX1 \keyTable_reg[3][2]  ( .D(n1059), .CLK(CLK), .Q(\keyTable[3][2] )
         );
  DFFPOSX1 \keyTable_reg[3][3]  ( .D(n1058), .CLK(CLK), .Q(\keyTable[3][3] )
         );
  DFFPOSX1 \keyTable_reg[3][4]  ( .D(n1057), .CLK(CLK), .Q(\keyTable[3][4] )
         );
  DFFPOSX1 \keyTable_reg[3][5]  ( .D(n1056), .CLK(CLK), .Q(\keyTable[3][5] )
         );
  DFFPOSX1 \keyTable_reg[3][6]  ( .D(n1055), .CLK(CLK), .Q(\keyTable[3][6] )
         );
  DFFPOSX1 \keyTable_reg[3][7]  ( .D(n1054), .CLK(CLK), .Q(\keyTable[3][7] )
         );
  DFFPOSX1 \keyTable_reg[2][0]  ( .D(n1053), .CLK(CLK), .Q(\keyTable[2][0] )
         );
  DFFPOSX1 \keyTable_reg[2][1]  ( .D(n1052), .CLK(CLK), .Q(\keyTable[2][1] )
         );
  DFFPOSX1 \keyTable_reg[2][2]  ( .D(n1051), .CLK(CLK), .Q(\keyTable[2][2] )
         );
  DFFPOSX1 \keyTable_reg[2][3]  ( .D(n1050), .CLK(CLK), .Q(\keyTable[2][3] )
         );
  DFFPOSX1 \keyTable_reg[2][4]  ( .D(n1049), .CLK(CLK), .Q(\keyTable[2][4] )
         );
  DFFPOSX1 \keyTable_reg[2][5]  ( .D(n1048), .CLK(CLK), .Q(\keyTable[2][5] )
         );
  DFFPOSX1 \keyTable_reg[2][6]  ( .D(n1047), .CLK(CLK), .Q(\keyTable[2][6] )
         );
  DFFPOSX1 \keyTable_reg[2][7]  ( .D(n1046), .CLK(CLK), .Q(\keyTable[2][7] )
         );
  DFFPOSX1 \keyTable_reg[1][0]  ( .D(n1045), .CLK(CLK), .Q(\keyTable[1][0] )
         );
  DFFPOSX1 \keyTable_reg[1][1]  ( .D(n1044), .CLK(CLK), .Q(\keyTable[1][1] )
         );
  DFFPOSX1 \keyTable_reg[1][2]  ( .D(n1043), .CLK(CLK), .Q(\keyTable[1][2] )
         );
  DFFPOSX1 \keyTable_reg[1][3]  ( .D(n1042), .CLK(CLK), .Q(\keyTable[1][3] )
         );
  DFFPOSX1 \keyTable_reg[1][4]  ( .D(n1041), .CLK(CLK), .Q(\keyTable[1][4] )
         );
  DFFPOSX1 \keyTable_reg[1][5]  ( .D(n1040), .CLK(CLK), .Q(\keyTable[1][5] )
         );
  DFFPOSX1 \keyTable_reg[1][6]  ( .D(n1039), .CLK(CLK), .Q(\keyTable[1][6] )
         );
  DFFPOSX1 \keyTable_reg[0][6]  ( .D(n1038), .CLK(CLK), .Q(\keyTable[0][6] )
         );
  DFFPOSX1 \keyTable_reg[0][5]  ( .D(n1037), .CLK(CLK), .Q(\keyTable[0][5] )
         );
  DFFPOSX1 \keyTable_reg[0][4]  ( .D(n1036), .CLK(CLK), .Q(\keyTable[0][4] )
         );
  DFFPOSX1 \keyTable_reg[0][3]  ( .D(n1035), .CLK(CLK), .Q(\keyTable[0][3] )
         );
  DFFPOSX1 \keyTable_reg[0][2]  ( .D(n1034), .CLK(CLK), .Q(\keyTable[0][2] )
         );
  DFFPOSX1 \keyTable_reg[0][1]  ( .D(n1033), .CLK(CLK), .Q(\keyTable[0][1] )
         );
  DFFPOSX1 \keyTable_reg[0][0]  ( .D(n1032), .CLK(CLK), .Q(\keyTable[0][0] )
         );
  DFFPOSX1 \keyTable_reg[1][7]  ( .D(n1031), .CLK(CLK), .Q(\keyTable[1][7] )
         );
  DFFPOSX1 \keyTable_reg[0][7]  ( .D(n1030), .CLK(CLK), .Q(\keyTable[0][7] )
         );
  DFFPOSX1 \prefillCounter_reg[7]  ( .D(n987), .CLK(CLK), .Q(prefillCounter[7]) );
  DFFPOSX1 \prefillCounter_reg[1]  ( .D(n988), .CLK(CLK), .Q(prefillCounter[1]) );
  DFFPOSX1 \prefillCounter_reg[2]  ( .D(n989), .CLK(CLK), .Q(prefillCounter[2]) );
  DFFPOSX1 \prefillCounter_reg[3]  ( .D(n990), .CLK(CLK), .Q(prefillCounter[3]) );
  DFFPOSX1 \prefillCounter_reg[4]  ( .D(n991), .CLK(CLK), .Q(prefillCounter[4]) );
  DFFPOSX1 \prefillCounter_reg[5]  ( .D(n992), .CLK(CLK), .Q(prefillCounter[5]) );
  DFFPOSX1 \prefillCounter_reg[6]  ( .D(n993), .CLK(CLK), .Q(prefillCounter[6]) );
  DFFPOSX1 \temp_reg[7]  ( .D(n1029), .CLK(CLK), .Q(temp[7]) );
  DFFPOSX1 \temp_reg[0]  ( .D(n1022), .CLK(CLK), .Q(temp[0]) );
  DFFPOSX1 \temp_reg[1]  ( .D(n1023), .CLK(CLK), .Q(temp[1]) );
  DFFPOSX1 \temp_reg[2]  ( .D(n1024), .CLK(CLK), .Q(temp[2]) );
  DFFPOSX1 \temp_reg[3]  ( .D(n1025), .CLK(CLK), .Q(temp[3]) );
  DFFPOSX1 \temp_reg[4]  ( .D(n1026), .CLK(CLK), .Q(temp[4]) );
  DFFPOSX1 \temp_reg[5]  ( .D(n1027), .CLK(CLK), .Q(temp[5]) );
  DFFPOSX1 \temp_reg[6]  ( .D(n1028), .CLK(CLK), .Q(temp[6]) );
  DFFPOSX1 \delaydata_reg[7]  ( .D(n383), .CLK(CLK), .Q(delaydata[7]) );
  DFFPOSX1 \delaydata_reg[0]  ( .D(n411), .CLK(CLK), .Q(delaydata[0]) );
  DFFPOSX1 \delaydata_reg[1]  ( .D(n407), .CLK(CLK), .Q(delaydata[1]) );
  DFFPOSX1 \delaydata_reg[2]  ( .D(n403), .CLK(CLK), .Q(delaydata[2]) );
  DFFPOSX1 \delaydata_reg[3]  ( .D(n399), .CLK(CLK), .Q(delaydata[3]) );
  DFFPOSX1 \delaydata_reg[4]  ( .D(n395), .CLK(CLK), .Q(delaydata[4]) );
  DFFPOSX1 \delaydata_reg[5]  ( .D(n391), .CLK(CLK), .Q(delaydata[5]) );
  DFFPOSX1 \delaydata_reg[6]  ( .D(n387), .CLK(CLK), .Q(delaydata[6]) );
  DFFPOSX1 \intj_reg[7]  ( .D(n1018), .CLK(CLK), .Q(intj[7]) );
  DFFPOSX1 \intj_reg[0]  ( .D(n1011), .CLK(CLK), .Q(intj[0]) );
  DFFPOSX1 \intj_reg[1]  ( .D(n1012), .CLK(CLK), .Q(intj[1]) );
  DFFPOSX1 \intj_reg[2]  ( .D(n1013), .CLK(CLK), .Q(intj[2]) );
  DFFPOSX1 \intj_reg[3]  ( .D(n1014), .CLK(CLK), .Q(intj[3]) );
  DFFPOSX1 \intj_reg[4]  ( .D(n1015), .CLK(CLK), .Q(intj[4]) );
  DFFPOSX1 \intj_reg[5]  ( .D(n1016), .CLK(CLK), .Q(intj[5]) );
  DFFPOSX1 \intj_reg[6]  ( .D(n1017), .CLK(CLK), .Q(intj[6]) );
  DFFPOSX1 \keyi_reg[2]  ( .D(n1019), .CLK(CLK), .Q(keyi[2]) );
  DFFPOSX1 \keyi_reg[1]  ( .D(n1020), .CLK(CLK), .Q(keyi[1]) );
  DFFPOSX1 \keyi_reg[0]  ( .D(n1021), .CLK(CLK), .Q(keyi[0]) );
  DFFPOSX1 \inti_reg[7]  ( .D(n437), .CLK(CLK), .Q(inti[7]) );
  DFFPOSX1 \inti_reg[0]  ( .D(n423), .CLK(CLK), .Q(inti[0]) );
  DFFPOSX1 \inti_reg[1]  ( .D(n425), .CLK(CLK), .Q(inti[1]) );
  DFFPOSX1 \inti_reg[2]  ( .D(n427), .CLK(CLK), .Q(inti[2]) );
  DFFPOSX1 \inti_reg[3]  ( .D(n429), .CLK(CLK), .Q(inti[3]) );
  DFFPOSX1 \inti_reg[4]  ( .D(n431), .CLK(CLK), .Q(inti[4]) );
  DFFPOSX1 \inti_reg[5]  ( .D(n433), .CLK(CLK), .Q(inti[5]) );
  DFFPOSX1 \inti_reg[6]  ( .D(n435), .CLK(CLK), .Q(inti[6]) );
  DFFPOSX1 \PROCESSED_DATA_reg[0]  ( .D(n1094), .CLK(CLK), .Q(
        PROCESSED_DATA[0]) );
  DFFPOSX1 \PROCESSED_DATA_reg[1]  ( .D(n1095), .CLK(CLK), .Q(
        PROCESSED_DATA[1]) );
  DFFPOSX1 \PROCESSED_DATA_reg[2]  ( .D(n1096), .CLK(CLK), .Q(
        PROCESSED_DATA[2]) );
  DFFPOSX1 \PROCESSED_DATA_reg[3]  ( .D(n1097), .CLK(CLK), .Q(
        PROCESSED_DATA[3]) );
  DFFPOSX1 \PROCESSED_DATA_reg[4]  ( .D(n1098), .CLK(CLK), .Q(
        PROCESSED_DATA[4]) );
  DFFPOSX1 \PROCESSED_DATA_reg[5]  ( .D(n1099), .CLK(CLK), .Q(
        PROCESSED_DATA[5]) );
  DFFPOSX1 \PROCESSED_DATA_reg[6]  ( .D(n1100), .CLK(CLK), .Q(
        PROCESSED_DATA[6]) );
  DFFPOSX1 \PROCESSED_DATA_reg[7]  ( .D(n1101), .CLK(CLK), .Q(
        PROCESSED_DATA[7]) );
  DFFPOSX1 \faddr_reg[7]  ( .D(n1102), .CLK(CLK), .Q(faddr[7]) );
  DFFPOSX1 \ADDR_reg[7]  ( .D(n1103), .CLK(CLK), .Q(ADDR[7]) );
  DFFPOSX1 \faddr_reg[6]  ( .D(n1104), .CLK(CLK), .Q(faddr[6]) );
  DFFPOSX1 \ADDR_reg[6]  ( .D(n1105), .CLK(CLK), .Q(ADDR[6]) );
  DFFPOSX1 \faddr_reg[5]  ( .D(n1106), .CLK(CLK), .Q(faddr[5]) );
  DFFPOSX1 \ADDR_reg[5]  ( .D(n1107), .CLK(CLK), .Q(ADDR[5]) );
  DFFPOSX1 \faddr_reg[4]  ( .D(n1108), .CLK(CLK), .Q(faddr[4]) );
  DFFPOSX1 \ADDR_reg[4]  ( .D(n1109), .CLK(CLK), .Q(ADDR[4]) );
  DFFPOSX1 \faddr_reg[3]  ( .D(n1110), .CLK(CLK), .Q(faddr[3]) );
  DFFPOSX1 \ADDR_reg[3]  ( .D(n1111), .CLK(CLK), .Q(ADDR[3]) );
  DFFPOSX1 \faddr_reg[2]  ( .D(n1112), .CLK(CLK), .Q(faddr[2]) );
  DFFPOSX1 \ADDR_reg[2]  ( .D(n1113), .CLK(CLK), .Q(ADDR[2]) );
  DFFPOSX1 \faddr_reg[1]  ( .D(n1114), .CLK(CLK), .Q(faddr[1]) );
  DFFPOSX1 \ADDR_reg[1]  ( .D(n1115), .CLK(CLK), .Q(ADDR[1]) );
  DFFPOSX1 \faddr_reg[0]  ( .D(n1116), .CLK(CLK), .Q(faddr[0]) );
  DFFPOSX1 \ADDR_reg[0]  ( .D(n1117), .CLK(CLK), .Q(ADDR[0]) );
  DFFPOSX1 \fdata_reg[7]  ( .D(n1118), .CLK(CLK), .Q(fdata[7]) );
  DFFPOSX1 \fdata_reg[6]  ( .D(n1119), .CLK(CLK), .Q(fdata[6]) );
  DFFPOSX1 \fdata_reg[5]  ( .D(n1120), .CLK(CLK), .Q(fdata[5]) );
  DFFPOSX1 \fdata_reg[4]  ( .D(n1121), .CLK(CLK), .Q(fdata[4]) );
  DFFPOSX1 \fdata_reg[3]  ( .D(n1122), .CLK(CLK), .Q(fdata[3]) );
  DFFPOSX1 \fdata_reg[2]  ( .D(n1123), .CLK(CLK), .Q(fdata[2]) );
  DFFPOSX1 \fdata_reg[1]  ( .D(n1124), .CLK(CLK), .Q(fdata[1]) );
  DFFPOSX1 \fdata_reg[0]  ( .D(n1125), .CLK(CLK), .Q(fdata[0]) );
  DFFPOSX1 fw_enable_reg ( .D(n1126), .CLK(CLK), .Q(fw_enable) );
  DFFPOSX1 fr_enable_reg ( .D(n1127), .CLK(CLK), .Q(fr_enable) );
  DFFPOSX1 W_ENABLE_reg ( .D(n1128), .CLK(CLK), .Q(W_ENABLE) );
  DFFPOSX1 R_ENABLE_reg ( .D(n1129), .CLK(CLK), .Q(R_ENABLE) );
  DFFPOSX1 \DATA_reg[7]  ( .D(n1130), .CLK(CLK), .Q(DATA[7]) );
  DFFPOSX1 \DATA_reg[6]  ( .D(n1131), .CLK(CLK), .Q(DATA[6]) );
  DFFPOSX1 \DATA_reg[5]  ( .D(n1132), .CLK(CLK), .Q(DATA[5]) );
  DFFPOSX1 \DATA_reg[4]  ( .D(n1133), .CLK(CLK), .Q(DATA[4]) );
  DFFPOSX1 \DATA_reg[3]  ( .D(n1134), .CLK(CLK), .Q(DATA[3]) );
  DFFPOSX1 \DATA_reg[2]  ( .D(n1135), .CLK(CLK), .Q(DATA[2]) );
  DFFPOSX1 \DATA_reg[1]  ( .D(n1136), .CLK(CLK), .Q(DATA[1]) );
  DFFPOSX1 \DATA_reg[0]  ( .D(n1137), .CLK(CLK), .Q(DATA[0]) );
  NOR2X1 U3 ( .A(n1602), .B(n577), .Y(n1153) );
  AOI22X1 U7 ( .A(n271), .B(extratemp[7]), .C(n604), .D(temp[7]), .Y(n1601) );
  OAI21X1 U8 ( .A(n463), .B(n976), .C(n1600), .Y(n1602) );
  AOI22X1 U9 ( .A(DATA_IN[7]), .B(n1599), .C(prefillCounter[7]), .D(n275), .Y(
        n1600) );
  NOR2X1 U10 ( .A(n1598), .B(n575), .Y(n1152) );
  AOI22X1 U12 ( .A(n271), .B(extratemp[6]), .C(n604), .D(temp[6]), .Y(n1597)
         );
  OAI21X1 U13 ( .A(n463), .B(n977), .C(n1596), .Y(n1598) );
  AOI22X1 U14 ( .A(DATA_IN[6]), .B(n1599), .C(prefillCounter[6]), .D(n275), 
        .Y(n1596) );
  NOR2X1 U15 ( .A(n1595), .B(n572), .Y(n1151) );
  AOI22X1 U17 ( .A(n271), .B(extratemp[5]), .C(n604), .D(temp[5]), .Y(n1594)
         );
  OAI21X1 U18 ( .A(n463), .B(n978), .C(n1593), .Y(n1595) );
  AOI22X1 U19 ( .A(DATA_IN[5]), .B(n1599), .C(prefillCounter[5]), .D(n275), 
        .Y(n1593) );
  NOR2X1 U20 ( .A(n1592), .B(n571), .Y(n1150) );
  AOI22X1 U22 ( .A(n271), .B(extratemp[4]), .C(n604), .D(temp[4]), .Y(n1591)
         );
  OAI21X1 U23 ( .A(n463), .B(n979), .C(n1590), .Y(n1592) );
  AOI22X1 U24 ( .A(DATA_IN[4]), .B(n1599), .C(prefillCounter[4]), .D(n275), 
        .Y(n1590) );
  NOR2X1 U25 ( .A(n1589), .B(n569), .Y(n1149) );
  AOI22X1 U27 ( .A(n271), .B(extratemp[3]), .C(n604), .D(temp[3]), .Y(n1588)
         );
  OAI21X1 U28 ( .A(n463), .B(n980), .C(n1587), .Y(n1589) );
  AOI22X1 U29 ( .A(DATA_IN[3]), .B(n1599), .C(prefillCounter[3]), .D(n275), 
        .Y(n1587) );
  NOR2X1 U30 ( .A(n1586), .B(n562), .Y(n1148) );
  AOI22X1 U32 ( .A(n271), .B(extratemp[2]), .C(n604), .D(temp[2]), .Y(n1585)
         );
  OAI21X1 U33 ( .A(n463), .B(n981), .C(n1584), .Y(n1586) );
  AOI22X1 U34 ( .A(DATA_IN[2]), .B(n1599), .C(prefillCounter[2]), .D(n275), 
        .Y(n1584) );
  NOR2X1 U35 ( .A(n1583), .B(n557), .Y(n1147) );
  AOI22X1 U37 ( .A(n271), .B(extratemp[1]), .C(n604), .D(temp[1]), .Y(n1582)
         );
  OAI21X1 U38 ( .A(n463), .B(n982), .C(n1581), .Y(n1583) );
  AOI22X1 U39 ( .A(DATA_IN[1]), .B(n1599), .C(prefillCounter[1]), .D(n275), 
        .Y(n1581) );
  NOR2X1 U40 ( .A(n1580), .B(n555), .Y(n1146) );
  AOI22X1 U42 ( .A(n271), .B(extratemp[0]), .C(n604), .D(temp[0]), .Y(n1579)
         );
  OAI21X1 U43 ( .A(n463), .B(n983), .C(n1578), .Y(n1580) );
  AOI22X1 U44 ( .A(DATA_IN[0]), .B(n1599), .C(prefillCounter[0]), .D(n275), 
        .Y(n1578) );
  NOR2X1 U46 ( .A(n1576), .B(n1575), .Y(n1145) );
  NAND2X1 U47 ( .A(n1574), .B(n1573), .Y(n1575) );
  AOI22X1 U48 ( .A(sj[7]), .B(n1572), .C(N448), .D(n282), .Y(n1573) );
  AOI22X1 U49 ( .A(intj[7]), .B(n280), .C(N503), .D(n268), .Y(n1574) );
  NAND2X1 U50 ( .A(n1570), .B(n1569), .Y(n1576) );
  AOI22X1 U51 ( .A(temp[7]), .B(n39), .C(inti[7]), .D(n1567), .Y(n1569) );
  AOI22X1 U52 ( .A(prefillCounter[7]), .B(n275), .C(faddr[7]), .D(n300), .Y(
        n1570) );
  NOR2X1 U53 ( .A(n1565), .B(n1564), .Y(n1144) );
  NAND2X1 U54 ( .A(n1563), .B(n1562), .Y(n1564) );
  AOI22X1 U55 ( .A(sj[6]), .B(n1572), .C(N447), .D(n282), .Y(n1562) );
  AOI22X1 U56 ( .A(intj[6]), .B(n280), .C(N502), .D(n268), .Y(n1563) );
  NAND2X1 U57 ( .A(n1561), .B(n1560), .Y(n1565) );
  AOI22X1 U58 ( .A(temp[6]), .B(n39), .C(inti[6]), .D(n1567), .Y(n1560) );
  AOI22X1 U59 ( .A(prefillCounter[6]), .B(n275), .C(faddr[6]), .D(n300), .Y(
        n1561) );
  NOR2X1 U60 ( .A(n1559), .B(n1558), .Y(n1143) );
  NAND2X1 U61 ( .A(n1557), .B(n1556), .Y(n1558) );
  AOI22X1 U62 ( .A(sj[5]), .B(n1572), .C(N446), .D(n282), .Y(n1556) );
  AOI22X1 U63 ( .A(intj[5]), .B(n280), .C(N501), .D(n268), .Y(n1557) );
  NAND2X1 U64 ( .A(n1555), .B(n1554), .Y(n1559) );
  AOI22X1 U65 ( .A(temp[5]), .B(n39), .C(inti[5]), .D(n1567), .Y(n1554) );
  AOI22X1 U66 ( .A(prefillCounter[5]), .B(n275), .C(faddr[5]), .D(n300), .Y(
        n1555) );
  NOR2X1 U67 ( .A(n1553), .B(n1552), .Y(n1142) );
  NAND2X1 U68 ( .A(n1551), .B(n1550), .Y(n1552) );
  AOI22X1 U69 ( .A(sj[4]), .B(n1572), .C(N445), .D(n282), .Y(n1550) );
  AOI22X1 U70 ( .A(intj[4]), .B(n280), .C(N500), .D(n268), .Y(n1551) );
  NAND2X1 U71 ( .A(n1549), .B(n1548), .Y(n1553) );
  AOI22X1 U72 ( .A(temp[4]), .B(n39), .C(inti[4]), .D(n1567), .Y(n1548) );
  AOI22X1 U73 ( .A(prefillCounter[4]), .B(n275), .C(faddr[4]), .D(n300), .Y(
        n1549) );
  NOR2X1 U74 ( .A(n1547), .B(n1546), .Y(n1141) );
  NAND2X1 U75 ( .A(n1545), .B(n1544), .Y(n1546) );
  AOI22X1 U76 ( .A(sj[3]), .B(n1572), .C(N444), .D(n282), .Y(n1544) );
  AOI22X1 U77 ( .A(intj[3]), .B(n280), .C(N499), .D(n268), .Y(n1545) );
  NAND2X1 U78 ( .A(n1543), .B(n1542), .Y(n1547) );
  AOI22X1 U79 ( .A(temp[3]), .B(n39), .C(inti[3]), .D(n1567), .Y(n1542) );
  AOI22X1 U80 ( .A(prefillCounter[3]), .B(n275), .C(faddr[3]), .D(n300), .Y(
        n1543) );
  NOR2X1 U81 ( .A(n1541), .B(n1540), .Y(n1140) );
  NAND2X1 U82 ( .A(n1539), .B(n1538), .Y(n1540) );
  AOI22X1 U83 ( .A(sj[2]), .B(n1572), .C(N443), .D(n282), .Y(n1538) );
  AOI22X1 U84 ( .A(intj[2]), .B(n280), .C(N498), .D(n268), .Y(n1539) );
  NAND2X1 U85 ( .A(n1537), .B(n1536), .Y(n1541) );
  AOI22X1 U86 ( .A(temp[2]), .B(n39), .C(inti[2]), .D(n1567), .Y(n1536) );
  AOI22X1 U87 ( .A(prefillCounter[2]), .B(n275), .C(faddr[2]), .D(n300), .Y(
        n1537) );
  NOR2X1 U88 ( .A(n1535), .B(n1534), .Y(n1139) );
  NAND2X1 U89 ( .A(n1533), .B(n1532), .Y(n1534) );
  AOI22X1 U90 ( .A(sj[1]), .B(n1572), .C(N442), .D(n282), .Y(n1532) );
  AOI22X1 U91 ( .A(intj[1]), .B(n280), .C(N497), .D(n268), .Y(n1533) );
  NAND2X1 U92 ( .A(n1531), .B(n1530), .Y(n1535) );
  AOI22X1 U93 ( .A(temp[1]), .B(n39), .C(inti[1]), .D(n1567), .Y(n1530) );
  AOI22X1 U94 ( .A(prefillCounter[1]), .B(n275), .C(faddr[1]), .D(n300), .Y(
        n1531) );
  NOR2X1 U95 ( .A(n1529), .B(n1528), .Y(n1138) );
  NAND2X1 U96 ( .A(n1527), .B(n1526), .Y(n1528) );
  AOI22X1 U97 ( .A(sj[0]), .B(n1572), .C(n932), .D(n282), .Y(n1526) );
  OAI21X1 U98 ( .A(n1525), .B(n1524), .C(n1523), .Y(n1572) );
  AOI22X1 U99 ( .A(intj[0]), .B(n280), .C(N496), .D(n268), .Y(n1527) );
  NAND2X1 U100 ( .A(n1522), .B(n1521), .Y(n1529) );
  AOI22X1 U101 ( .A(temp[0]), .B(n39), .C(inti[0]), .D(n1567), .Y(n1521) );
  OAI21X1 U102 ( .A(n1520), .B(n1519), .C(n516), .Y(n1567) );
  AOI22X1 U104 ( .A(prefillCounter[0]), .B(n275), .C(faddr[0]), .D(n300), .Y(
        n1522) );
  OAI21X1 U106 ( .A(n252), .B(n630), .C(n277), .Y(n1516) );
  OAI21X1 U108 ( .A(n1515), .B(n1514), .C(n1513), .Y(n1517) );
  AOI21X1 U109 ( .A(n1512), .B(n1511), .C(n553), .Y(n1513) );
  NOR2X1 U110 ( .A(KEY_ERROR), .B(n1510), .Y(n1512) );
  OAI21X1 U111 ( .A(n373), .B(n1509), .C(n371), .Y(n1514) );
  NAND3X1 U112 ( .A(n1508), .B(n1507), .C(n1506), .Y(nextState[3]) );
  AOI21X1 U113 ( .A(n600), .B(n629), .C(n1505), .Y(n1506) );
  NAND2X1 U114 ( .A(n1504), .B(n1503), .Y(n1505) );
  AOI22X1 U115 ( .A(n1502), .B(n371), .C(n547), .D(n1501), .Y(n1508) );
  NAND3X1 U116 ( .A(n1500), .B(n1499), .C(n1498), .Y(nextState[2]) );
  NOR2X1 U117 ( .A(n1497), .B(n1496), .Y(n1498) );
  OAI21X1 U118 ( .A(n1495), .B(n1525), .C(n1507), .Y(n1496) );
  AOI21X1 U119 ( .A(n1494), .B(permuteComplete), .C(n1493), .Y(n1507) );
  NAND2X1 U120 ( .A(n249), .B(n1492), .Y(n1493) );
  OAI22X1 U121 ( .A(n1519), .B(n1491), .C(KEY_ERROR), .D(n1490), .Y(n1497) );
  AOI22X1 U122 ( .A(n1489), .B(n1488), .C(n1487), .D(n1486), .Y(n1490) );
  NOR2X1 U123 ( .A(n1485), .B(n373), .Y(n1489) );
  NOR2X1 U124 ( .A(n271), .B(n618), .Y(n1499) );
  NOR2X1 U125 ( .A(n616), .B(n1484), .Y(n1500) );
  NAND3X1 U126 ( .A(n1483), .B(n1482), .C(n1481), .Y(nextState[1]) );
  NOR2X1 U127 ( .A(n1480), .B(n1479), .Y(n1481) );
  OAI21X1 U128 ( .A(n1478), .B(n1477), .C(n220), .Y(n1479) );
  NAND3X1 U129 ( .A(n1475), .B(n413), .C(n1474), .Y(n1477) );
  NOR2X1 U130 ( .A(prefillCounter[2]), .B(prefillCounter[1]), .Y(n1474) );
  NAND3X1 U131 ( .A(n1473), .B(n922), .C(n1472), .Y(n1478) );
  NOR2X1 U132 ( .A(prefillCounter[4]), .B(prefillCounter[3]), .Y(n1472) );
  NOR2X1 U133 ( .A(prefillCounter[7]), .B(prefillCounter[6]), .Y(n1473) );
  AOI22X1 U135 ( .A(n1471), .B(state[0]), .C(n1470), .D(n371), .Y(n1483) );
  OAI21X1 U137 ( .A(n542), .B(n1486), .C(n1469), .Y(n1470) );
  NAND2X1 U138 ( .A(n1501), .B(n1468), .Y(n1469) );
  OAI21X1 U139 ( .A(n1467), .B(n1486), .C(n1466), .Y(n1468) );
  OAI21X1 U140 ( .A(n1485), .B(n373), .C(n594), .Y(n1466) );
  NAND3X1 U143 ( .A(n379), .B(n377), .C(BYTE_READY), .Y(n1486) );
  NOR2X1 U145 ( .A(state[1]), .B(n1519), .Y(n1471) );
  NAND3X1 U146 ( .A(n1464), .B(n1463), .C(n1462), .Y(nextState[0]) );
  NOR2X1 U147 ( .A(n282), .B(n1461), .Y(n1462) );
  OAI21X1 U148 ( .A(KEY_ERROR), .B(n1460), .C(n1482), .Y(n1461) );
  NOR2X1 U149 ( .A(n1459), .B(n1458), .Y(n1482) );
  OAI21X1 U150 ( .A(permuteComplete), .B(n592), .C(n1457), .Y(n1458) );
  NAND3X1 U151 ( .A(n1492), .B(n1456), .C(n1455), .Y(n1459) );
  AOI21X1 U152 ( .A(n1488), .B(n1510), .C(n1454), .Y(n1460) );
  OAI21X1 U153 ( .A(n252), .B(n1453), .C(n1452), .Y(n1454) );
  NAND3X1 U154 ( .A(BYTE_READY), .B(n1487), .C(n375), .Y(n1452) );
  NAND2X1 U156 ( .A(OPCODE[0]), .B(n377), .Y(n1509) );
  NAND2X1 U158 ( .A(BYTE_READY), .B(n1451), .Y(n1510) );
  OAI21X1 U159 ( .A(OPCODE[0]), .B(OPCODE[1]), .C(n1465), .Y(n1451) );
  NAND2X1 U160 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n1465) );
  NOR2X1 U161 ( .A(n553), .B(n271), .Y(n1463) );
  NOR2X1 U162 ( .A(n1475), .B(n1450), .Y(n1464) );
  OAI21X1 U163 ( .A(n318), .B(n415), .C(n1449), .Y(n1137) );
  NAND2X1 U164 ( .A(DATA[0]), .B(n305), .Y(n1449) );
  OAI21X1 U165 ( .A(n326), .B(n462), .C(n1448), .Y(n1136) );
  NAND2X1 U166 ( .A(DATA[1]), .B(n327), .Y(n1448) );
  OAI21X1 U167 ( .A(n326), .B(n459), .C(n1447), .Y(n1135) );
  NAND2X1 U168 ( .A(DATA[2]), .B(n327), .Y(n1447) );
  OAI21X1 U169 ( .A(n326), .B(n458), .C(n1446), .Y(n1134) );
  NAND2X1 U170 ( .A(DATA[3]), .B(n327), .Y(n1446) );
  OAI21X1 U171 ( .A(n326), .B(n455), .C(n1445), .Y(n1133) );
  NAND2X1 U172 ( .A(DATA[4]), .B(RST), .Y(n1445) );
  OAI21X1 U173 ( .A(n326), .B(n453), .C(n1444), .Y(n1132) );
  NAND2X1 U174 ( .A(DATA[5]), .B(n327), .Y(n1444) );
  OAI21X1 U175 ( .A(n326), .B(n451), .C(n1443), .Y(n1131) );
  NAND2X1 U176 ( .A(DATA[6]), .B(n327), .Y(n1443) );
  OAI21X1 U177 ( .A(n326), .B(n449), .C(n1442), .Y(n1130) );
  NAND2X1 U178 ( .A(DATA[7]), .B(n327), .Y(n1442) );
  OAI21X1 U179 ( .A(n326), .B(n1441), .C(n1440), .Y(n1129) );
  NAND2X1 U180 ( .A(R_ENABLE), .B(n327), .Y(n1440) );
  AOI21X1 U181 ( .A(fr_enable), .B(n1439), .C(n1438), .Y(n1441) );
  OAI21X1 U182 ( .A(n318), .B(n1437), .C(n1436), .Y(n1128) );
  NAND2X1 U183 ( .A(W_ENABLE), .B(n326), .Y(n1436) );
  AOI21X1 U184 ( .A(fw_enable), .B(n1435), .C(n1434), .Y(n1437) );
  OAI21X1 U185 ( .A(n318), .B(n518), .C(n1433), .Y(n1127) );
  OAI21X1 U186 ( .A(n318), .B(n1439), .C(fr_enable), .Y(n1433) );
  NAND3X1 U187 ( .A(n1432), .B(n1431), .C(n1430), .Y(n1439) );
  NOR2X1 U188 ( .A(n606), .B(n1429), .Y(n1430) );
  NAND2X1 U189 ( .A(n247), .B(n44), .Y(n1429) );
  NAND2X1 U191 ( .A(n610), .B(n624), .Y(n1523) );
  OAI21X1 U192 ( .A(n318), .B(n528), .C(n1428), .Y(n1126) );
  OAI21X1 U193 ( .A(n318), .B(n1435), .C(fw_enable), .Y(n1428) );
  NAND3X1 U195 ( .A(n247), .B(n44), .C(n1427), .Y(n1434) );
  NOR2X1 U196 ( .A(n1599), .B(n604), .Y(n1427) );
  OAI22X1 U197 ( .A(n343), .B(n983), .C(n317), .D(n415), .Y(n1125) );
  OAI22X1 U200 ( .A(n343), .B(n982), .C(n311), .D(n462), .Y(n1124) );
  OAI22X1 U203 ( .A(n343), .B(n981), .C(n317), .D(n459), .Y(n1123) );
  OAI22X1 U206 ( .A(n343), .B(n980), .C(n311), .D(n458), .Y(n1122) );
  OAI22X1 U209 ( .A(n345), .B(n979), .C(n317), .D(n455), .Y(n1121) );
  OAI22X1 U212 ( .A(n341), .B(n978), .C(n311), .D(n453), .Y(n1120) );
  OAI22X1 U215 ( .A(n341), .B(n977), .C(n317), .D(n451), .Y(n1119) );
  OAI22X1 U218 ( .A(n341), .B(n976), .C(n311), .D(n449), .Y(n1118) );
  OAI21X1 U221 ( .A(n318), .B(n417), .C(n1426), .Y(n1117) );
  NAND2X1 U222 ( .A(ADDR[0]), .B(n326), .Y(n1426) );
  OAI22X1 U223 ( .A(n337), .B(n975), .C(n311), .D(n417), .Y(n1116) );
  OAI21X1 U226 ( .A(n318), .B(n501), .C(n1425), .Y(n1115) );
  NAND2X1 U227 ( .A(ADDR[1]), .B(n327), .Y(n1425) );
  OAI22X1 U228 ( .A(n347), .B(n974), .C(n311), .D(n501), .Y(n1114) );
  OAI21X1 U231 ( .A(n318), .B(n503), .C(n1424), .Y(n1113) );
  NAND2X1 U232 ( .A(ADDR[2]), .B(n326), .Y(n1424) );
  OAI22X1 U233 ( .A(n349), .B(n973), .C(n311), .D(n503), .Y(n1112) );
  OAI21X1 U236 ( .A(n318), .B(n504), .C(n1423), .Y(n1111) );
  NAND2X1 U237 ( .A(ADDR[3]), .B(n327), .Y(n1423) );
  OAI22X1 U238 ( .A(n339), .B(n972), .C(n311), .D(n504), .Y(n1110) );
  OAI21X1 U241 ( .A(n318), .B(n505), .C(n1422), .Y(n1109) );
  NAND2X1 U242 ( .A(ADDR[4]), .B(n327), .Y(n1422) );
  OAI22X1 U243 ( .A(n329), .B(n971), .C(n311), .D(n505), .Y(n1108) );
  OAI21X1 U246 ( .A(n318), .B(n506), .C(n1421), .Y(n1107) );
  NAND2X1 U247 ( .A(ADDR[5]), .B(n327), .Y(n1421) );
  OAI22X1 U248 ( .A(n335), .B(n970), .C(n311), .D(n506), .Y(n1106) );
  OAI21X1 U251 ( .A(n317), .B(n507), .C(n1420), .Y(n1105) );
  NAND2X1 U252 ( .A(ADDR[6]), .B(n327), .Y(n1420) );
  OAI22X1 U253 ( .A(n333), .B(n969), .C(n311), .D(n507), .Y(n1104) );
  OAI21X1 U256 ( .A(n317), .B(n509), .C(n1419), .Y(n1103) );
  NAND2X1 U257 ( .A(ADDR[7]), .B(n327), .Y(n1419) );
  OAI22X1 U258 ( .A(n331), .B(n968), .C(n311), .D(n509), .Y(n1102) );
  OAI21X1 U261 ( .A(n317), .B(n381), .C(n1418), .Y(n1101) );
  NAND2X1 U262 ( .A(PROCESSED_DATA[7]), .B(n327), .Y(n1418) );
  OAI21X1 U264 ( .A(n512), .B(n967), .C(n1417), .Y(nextProcessedData[7]) );
  AOI22X1 U265 ( .A(n37), .B(n1415), .C(BYTE[7]), .D(n605), .Y(n1417) );
  XOR2X1 U266 ( .A(temp[7]), .B(delaydata[7]), .Y(n1415) );
  OAI21X1 U268 ( .A(n317), .B(n385), .C(n1414), .Y(n1100) );
  NAND2X1 U269 ( .A(PROCESSED_DATA[6]), .B(n327), .Y(n1414) );
  OAI21X1 U271 ( .A(n512), .B(n966), .C(n1413), .Y(nextProcessedData[6]) );
  AOI22X1 U272 ( .A(n37), .B(n1412), .C(BYTE[6]), .D(n605), .Y(n1413) );
  XOR2X1 U273 ( .A(temp[6]), .B(delaydata[6]), .Y(n1412) );
  OAI21X1 U275 ( .A(n317), .B(n389), .C(n1411), .Y(n1099) );
  NAND2X1 U276 ( .A(PROCESSED_DATA[5]), .B(n327), .Y(n1411) );
  OAI21X1 U278 ( .A(n512), .B(n965), .C(n1410), .Y(nextProcessedData[5]) );
  AOI22X1 U279 ( .A(n37), .B(n1409), .C(BYTE[5]), .D(n605), .Y(n1410) );
  XOR2X1 U280 ( .A(temp[5]), .B(delaydata[5]), .Y(n1409) );
  OAI21X1 U282 ( .A(n317), .B(n393), .C(n1408), .Y(n1098) );
  NAND2X1 U283 ( .A(PROCESSED_DATA[4]), .B(n327), .Y(n1408) );
  OAI21X1 U285 ( .A(n512), .B(n964), .C(n1407), .Y(nextProcessedData[4]) );
  AOI22X1 U286 ( .A(n37), .B(n1406), .C(BYTE[4]), .D(n605), .Y(n1407) );
  XOR2X1 U287 ( .A(temp[4]), .B(delaydata[4]), .Y(n1406) );
  OAI21X1 U289 ( .A(n318), .B(n397), .C(n1405), .Y(n1097) );
  NAND2X1 U290 ( .A(PROCESSED_DATA[3]), .B(n327), .Y(n1405) );
  OAI21X1 U292 ( .A(n512), .B(n963), .C(n1404), .Y(nextProcessedData[3]) );
  AOI22X1 U293 ( .A(n37), .B(n1403), .C(BYTE[3]), .D(n605), .Y(n1404) );
  XOR2X1 U294 ( .A(temp[3]), .B(delaydata[3]), .Y(n1403) );
  OAI21X1 U296 ( .A(n317), .B(n401), .C(n1402), .Y(n1096) );
  NAND2X1 U297 ( .A(PROCESSED_DATA[2]), .B(n327), .Y(n1402) );
  OAI21X1 U299 ( .A(n512), .B(n962), .C(n1401), .Y(nextProcessedData[2]) );
  AOI22X1 U300 ( .A(n37), .B(n1400), .C(BYTE[2]), .D(n605), .Y(n1401) );
  XOR2X1 U301 ( .A(temp[2]), .B(delaydata[2]), .Y(n1400) );
  OAI21X1 U303 ( .A(n317), .B(n405), .C(n1399), .Y(n1095) );
  NAND2X1 U304 ( .A(PROCESSED_DATA[1]), .B(RST), .Y(n1399) );
  OAI21X1 U306 ( .A(n512), .B(n961), .C(n1398), .Y(nextProcessedData[1]) );
  AOI22X1 U307 ( .A(n37), .B(n1397), .C(BYTE[1]), .D(n605), .Y(n1398) );
  XOR2X1 U308 ( .A(temp[1]), .B(delaydata[1]), .Y(n1397) );
  OAI21X1 U310 ( .A(n317), .B(n409), .C(n1396), .Y(n1094) );
  NAND2X1 U311 ( .A(PROCESSED_DATA[0]), .B(RST), .Y(n1396) );
  OAI21X1 U313 ( .A(n512), .B(n960), .C(n1395), .Y(nextProcessedData[0]) );
  AOI22X1 U314 ( .A(n37), .B(n1394), .C(BYTE[0]), .D(n605), .Y(n1395) );
  XOR2X1 U315 ( .A(temp[0]), .B(delaydata[0]), .Y(n1394) );
  NAND3X1 U318 ( .A(n285), .B(n520), .C(n1392), .Y(n1393) );
  NOR2X1 U319 ( .A(n1391), .B(n1390), .Y(n1392) );
  AOI22X1 U322 ( .A(BYTE[7]), .B(n241), .C(n302), .D(delaydata[7]), .Y(n1388)
         );
  AOI22X1 U324 ( .A(BYTE[0]), .B(n241), .C(n302), .D(delaydata[0]), .Y(n1387)
         );
  AOI22X1 U326 ( .A(BYTE[1]), .B(n241), .C(n302), .D(delaydata[1]), .Y(n1386)
         );
  AOI22X1 U328 ( .A(BYTE[2]), .B(n241), .C(n302), .D(delaydata[2]), .Y(n1385)
         );
  AOI22X1 U330 ( .A(BYTE[3]), .B(n241), .C(n302), .D(delaydata[3]), .Y(n1384)
         );
  AOI22X1 U332 ( .A(BYTE[4]), .B(n241), .C(n302), .D(delaydata[4]), .Y(n1383)
         );
  AOI22X1 U334 ( .A(BYTE[5]), .B(n241), .C(n302), .D(delaydata[5]), .Y(n1382)
         );
  AOI22X1 U336 ( .A(BYTE[6]), .B(n241), .C(n302), .D(delaydata[6]), .Y(n1381)
         );
  OAI21X1 U339 ( .A(n20), .B(n637), .C(n1379), .Y(n1093) );
  NAND2X1 U340 ( .A(KEY[56]), .B(n7), .Y(n1379) );
  OAI21X1 U342 ( .A(n12), .B(n638), .C(n1378), .Y(n1092) );
  NAND2X1 U343 ( .A(KEY[57]), .B(n15), .Y(n1378) );
  OAI21X1 U345 ( .A(n10), .B(n648), .C(n1377), .Y(n1091) );
  NAND2X1 U346 ( .A(KEY[58]), .B(n16), .Y(n1377) );
  OAI21X1 U348 ( .A(n9), .B(n649), .C(n1376), .Y(n1090) );
  NAND2X1 U349 ( .A(KEY[59]), .B(n20), .Y(n1376) );
  OAI21X1 U351 ( .A(n8), .B(n650), .C(n1375), .Y(n1089) );
  NAND2X1 U352 ( .A(KEY[60]), .B(n17), .Y(n1375) );
  OAI21X1 U354 ( .A(n7), .B(n651), .C(n1374), .Y(n1088) );
  NAND2X1 U355 ( .A(KEY[61]), .B(n10), .Y(n1374) );
  OAI21X1 U357 ( .A(n12), .B(n692), .C(n1373), .Y(n1087) );
  NAND2X1 U358 ( .A(KEY[62]), .B(n14), .Y(n1373) );
  OAI21X1 U360 ( .A(n10), .B(n701), .C(n1372), .Y(n1086) );
  NAND2X1 U361 ( .A(KEY[63]), .B(n12), .Y(n1372) );
  OAI21X1 U363 ( .A(n9), .B(n746), .C(n1371), .Y(n1085) );
  NAND2X1 U364 ( .A(KEY[48]), .B(n14), .Y(n1371) );
  OAI21X1 U366 ( .A(n8), .B(n748), .C(n1370), .Y(n1084) );
  NAND2X1 U367 ( .A(KEY[49]), .B(n15), .Y(n1370) );
  OAI21X1 U369 ( .A(n9), .B(n750), .C(n1369), .Y(n1083) );
  NAND2X1 U370 ( .A(KEY[50]), .B(n12), .Y(n1369) );
  OAI21X1 U372 ( .A(n8), .B(n752), .C(n1368), .Y(n1082) );
  NAND2X1 U373 ( .A(KEY[51]), .B(n20), .Y(n1368) );
  OAI21X1 U375 ( .A(n7), .B(n754), .C(n1367), .Y(n1081) );
  NAND2X1 U376 ( .A(KEY[52]), .B(n24), .Y(n1367) );
  OAI21X1 U378 ( .A(n6), .B(n756), .C(n1366), .Y(n1080) );
  NAND2X1 U379 ( .A(KEY[53]), .B(n16), .Y(n1366) );
  OAI21X1 U381 ( .A(n20), .B(n758), .C(n1365), .Y(n1079) );
  NAND2X1 U382 ( .A(KEY[54]), .B(n29), .Y(n1365) );
  OAI21X1 U384 ( .A(n17), .B(n760), .C(n1364), .Y(n1078) );
  NAND2X1 U385 ( .A(KEY[55]), .B(n9), .Y(n1364) );
  OAI21X1 U387 ( .A(n16), .B(n761), .C(n1363), .Y(n1077) );
  NAND2X1 U388 ( .A(KEY[40]), .B(n22), .Y(n1363) );
  OAI21X1 U390 ( .A(n17), .B(n762), .C(n1362), .Y(n1076) );
  NAND2X1 U391 ( .A(KEY[41]), .B(n27), .Y(n1362) );
  OAI21X1 U393 ( .A(n16), .B(n763), .C(n1361), .Y(n1075) );
  NAND2X1 U394 ( .A(KEY[42]), .B(n12), .Y(n1361) );
  OAI21X1 U396 ( .A(n15), .B(n764), .C(n1360), .Y(n1074) );
  NAND2X1 U397 ( .A(KEY[43]), .B(n6), .Y(n1360) );
  OAI21X1 U399 ( .A(n14), .B(n765), .C(n1359), .Y(n1073) );
  NAND2X1 U400 ( .A(KEY[44]), .B(n14), .Y(n1359) );
  OAI21X1 U402 ( .A(n15), .B(n766), .C(n1358), .Y(n1072) );
  NAND2X1 U403 ( .A(KEY[45]), .B(n15), .Y(n1358) );
  OAI21X1 U405 ( .A(n14), .B(n767), .C(n1357), .Y(n1071) );
  NAND2X1 U406 ( .A(KEY[46]), .B(n10), .Y(n1357) );
  OAI21X1 U408 ( .A(n12), .B(n768), .C(n1356), .Y(n1070) );
  NAND2X1 U409 ( .A(KEY[47]), .B(n17), .Y(n1356) );
  OAI21X1 U411 ( .A(n10), .B(n769), .C(n1355), .Y(n1069) );
  NAND2X1 U412 ( .A(KEY[32]), .B(n9), .Y(n1355) );
  OAI21X1 U414 ( .A(n15), .B(n770), .C(n1354), .Y(n1068) );
  NAND2X1 U415 ( .A(KEY[33]), .B(n10), .Y(n1354) );
  OAI21X1 U417 ( .A(n14), .B(n771), .C(n1353), .Y(n1067) );
  NAND2X1 U418 ( .A(KEY[34]), .B(n27), .Y(n1353) );
  OAI21X1 U420 ( .A(n6), .B(n772), .C(n1352), .Y(n1066) );
  NAND2X1 U421 ( .A(KEY[35]), .B(n6), .Y(n1352) );
  OAI21X1 U423 ( .A(n29), .B(n773), .C(n1351), .Y(n1065) );
  NAND2X1 U424 ( .A(KEY[36]), .B(n16), .Y(n1351) );
  OAI21X1 U426 ( .A(n27), .B(n774), .C(n1350), .Y(n1064) );
  NAND2X1 U427 ( .A(KEY[37]), .B(n8), .Y(n1350) );
  OAI21X1 U429 ( .A(n24), .B(n775), .C(n1349), .Y(n1063) );
  NAND2X1 U430 ( .A(KEY[38]), .B(n6), .Y(n1349) );
  OAI21X1 U432 ( .A(n22), .B(n776), .C(n1348), .Y(n1062) );
  NAND2X1 U433 ( .A(KEY[39]), .B(n9), .Y(n1348) );
  OAI21X1 U435 ( .A(n15), .B(n777), .C(n1347), .Y(n1061) );
  NAND2X1 U436 ( .A(KEY[24]), .B(n6), .Y(n1347) );
  OAI21X1 U437 ( .A(n17), .B(n778), .C(n1346), .Y(n1060) );
  NAND2X1 U438 ( .A(KEY[25]), .B(n7), .Y(n1346) );
  OAI21X1 U439 ( .A(n7), .B(n779), .C(n1345), .Y(n1059) );
  NAND2X1 U440 ( .A(KEY[26]), .B(n29), .Y(n1345) );
  OAI21X1 U441 ( .A(n6), .B(n780), .C(n1344), .Y(n1058) );
  NAND2X1 U442 ( .A(KEY[27]), .B(n8), .Y(n1344) );
  OAI21X1 U443 ( .A(n29), .B(n781), .C(n1343), .Y(n1057) );
  NAND2X1 U444 ( .A(KEY[28]), .B(n7), .Y(n1343) );
  OAI21X1 U445 ( .A(n27), .B(n782), .C(n1342), .Y(n1056) );
  NAND2X1 U446 ( .A(KEY[29]), .B(n29), .Y(n1342) );
  OAI21X1 U447 ( .A(n29), .B(n783), .C(n1341), .Y(n1055) );
  NAND2X1 U448 ( .A(KEY[30]), .B(n7), .Y(n1341) );
  OAI21X1 U449 ( .A(n27), .B(n784), .C(n1340), .Y(n1054) );
  NAND2X1 U450 ( .A(KEY[31]), .B(n8), .Y(n1340) );
  OAI21X1 U451 ( .A(n24), .B(n785), .C(n1339), .Y(n1053) );
  NAND2X1 U452 ( .A(KEY[16]), .B(n24), .Y(n1339) );
  OAI21X1 U453 ( .A(n22), .B(n786), .C(n1338), .Y(n1052) );
  NAND2X1 U454 ( .A(KEY[17]), .B(n16), .Y(n1338) );
  OAI21X1 U455 ( .A(n16), .B(n787), .C(n1337), .Y(n1051) );
  NAND2X1 U456 ( .A(KEY[18]), .B(n22), .Y(n1337) );
  OAI21X1 U457 ( .A(n12), .B(n788), .C(n1336), .Y(n1050) );
  NAND2X1 U458 ( .A(KEY[19]), .B(n27), .Y(n1336) );
  OAI21X1 U459 ( .A(n10), .B(n789), .C(n1335), .Y(n1049) );
  NAND2X1 U460 ( .A(KEY[20]), .B(n24), .Y(n1335) );
  OAI21X1 U461 ( .A(n20), .B(n790), .C(n1334), .Y(n1048) );
  NAND2X1 U462 ( .A(KEY[21]), .B(n20), .Y(n1334) );
  OAI21X1 U463 ( .A(n14), .B(n791), .C(n1333), .Y(n1047) );
  NAND2X1 U464 ( .A(KEY[22]), .B(n29), .Y(n1333) );
  OAI21X1 U465 ( .A(n9), .B(n864), .C(n1332), .Y(n1046) );
  NAND2X1 U466 ( .A(KEY[23]), .B(n27), .Y(n1332) );
  OAI21X1 U467 ( .A(n9), .B(n865), .C(n1331), .Y(n1045) );
  NAND2X1 U468 ( .A(KEY[8]), .B(n6), .Y(n1331) );
  OAI21X1 U469 ( .A(n8), .B(n866), .C(n1330), .Y(n1044) );
  NAND2X1 U470 ( .A(KEY[9]), .B(n12), .Y(n1330) );
  OAI21X1 U471 ( .A(n22), .B(n867), .C(n1329), .Y(n1043) );
  NAND2X1 U472 ( .A(KEY[10]), .B(n20), .Y(n1329) );
  OAI21X1 U473 ( .A(n7), .B(n868), .C(n1328), .Y(n1042) );
  NAND2X1 U474 ( .A(KEY[11]), .B(n14), .Y(n1328) );
  OAI21X1 U475 ( .A(n6), .B(n869), .C(n1327), .Y(n1041) );
  NAND2X1 U476 ( .A(KEY[12]), .B(n15), .Y(n1327) );
  OAI21X1 U477 ( .A(n8), .B(n870), .C(n1326), .Y(n1040) );
  NAND2X1 U478 ( .A(KEY[13]), .B(n24), .Y(n1326) );
  OAI21X1 U479 ( .A(n24), .B(n871), .C(n1325), .Y(n1039) );
  NAND2X1 U480 ( .A(KEY[14]), .B(n22), .Y(n1325) );
  OAI21X1 U481 ( .A(n24), .B(n883), .C(n1324), .Y(n1038) );
  NAND2X1 U482 ( .A(KEY[6]), .B(n10), .Y(n1324) );
  OAI21X1 U483 ( .A(n17), .B(n884), .C(n1323), .Y(n1037) );
  NAND2X1 U484 ( .A(KEY[5]), .B(n17), .Y(n1323) );
  OAI21X1 U485 ( .A(n15), .B(n885), .C(n1322), .Y(n1036) );
  NAND2X1 U486 ( .A(KEY[4]), .B(n8), .Y(n1322) );
  OAI21X1 U487 ( .A(n14), .B(n886), .C(n1321), .Y(n1035) );
  NAND2X1 U488 ( .A(KEY[3]), .B(n9), .Y(n1321) );
  OAI21X1 U489 ( .A(n27), .B(n887), .C(n1320), .Y(n1034) );
  NAND2X1 U490 ( .A(KEY[2]), .B(n7), .Y(n1320) );
  OAI21X1 U491 ( .A(n29), .B(n888), .C(n1319), .Y(n1033) );
  NAND2X1 U492 ( .A(KEY[1]), .B(n22), .Y(n1319) );
  OAI21X1 U493 ( .A(n12), .B(n889), .C(n1318), .Y(n1032) );
  NAND2X1 U494 ( .A(KEY[0]), .B(n20), .Y(n1318) );
  OAI21X1 U495 ( .A(n22), .B(n890), .C(n1317), .Y(n1031) );
  NAND2X1 U496 ( .A(KEY[15]), .B(n17), .Y(n1317) );
  OAI21X1 U497 ( .A(n10), .B(n916), .C(n1316), .Y(n1030) );
  NAND2X1 U498 ( .A(KEY[7]), .B(n16), .Y(n1316) );
  NOR2X1 U499 ( .A(n1315), .B(n1391), .Y(n1380) );
  OAI21X1 U500 ( .A(n500), .B(n924), .C(n1314), .Y(n1029) );
  AOI22X1 U501 ( .A(N527), .B(n1313), .C(n237), .D(DATA_IN[7]), .Y(n1314) );
  OAI21X1 U503 ( .A(n500), .B(n931), .C(n1312), .Y(n1028) );
  AOI22X1 U504 ( .A(N526), .B(n1313), .C(n237), .D(DATA_IN[6]), .Y(n1312) );
  OAI21X1 U506 ( .A(n500), .B(n930), .C(n1311), .Y(n1027) );
  AOI22X1 U507 ( .A(N525), .B(n1313), .C(n237), .D(DATA_IN[5]), .Y(n1311) );
  OAI21X1 U509 ( .A(n500), .B(n929), .C(n1310), .Y(n1026) );
  AOI22X1 U510 ( .A(N524), .B(n1313), .C(n237), .D(DATA_IN[4]), .Y(n1310) );
  OAI21X1 U512 ( .A(n500), .B(n928), .C(n1309), .Y(n1025) );
  AOI22X1 U513 ( .A(N523), .B(n1313), .C(n237), .D(DATA_IN[3]), .Y(n1309) );
  OAI21X1 U515 ( .A(n500), .B(n927), .C(n1308), .Y(n1024) );
  AOI22X1 U516 ( .A(N522), .B(n1313), .C(n237), .D(DATA_IN[2]), .Y(n1308) );
  OAI21X1 U518 ( .A(n500), .B(n926), .C(n1307), .Y(n1023) );
  AOI22X1 U519 ( .A(N521), .B(n1313), .C(n237), .D(DATA_IN[1]), .Y(n1307) );
  OAI21X1 U521 ( .A(n500), .B(n925), .C(n1306), .Y(n1022) );
  AOI22X1 U522 ( .A(N520), .B(n1313), .C(n237), .D(DATA_IN[0]), .Y(n1306) );
  NAND3X1 U527 ( .A(n1303), .B(n522), .C(n1302), .Y(n1305) );
  NOR2X1 U528 ( .A(n1389), .B(n300), .Y(n1302) );
  NAND2X1 U529 ( .A(n1431), .B(n545), .Y(n1566) );
  NAND3X1 U530 ( .A(n1301), .B(n247), .C(n1300), .Y(n1389) );
  NOR2X1 U532 ( .A(n326), .B(n1475), .Y(n1303) );
  AOI22X1 U534 ( .A(n295), .B(extratemp[0]), .C(DATA_IN[0]), .D(n292), .Y(
        n1298) );
  AOI22X1 U536 ( .A(n295), .B(extratemp[1]), .C(DATA_IN[1]), .D(n292), .Y(
        n1296) );
  AOI22X1 U538 ( .A(n295), .B(extratemp[2]), .C(DATA_IN[2]), .D(n292), .Y(
        n1295) );
  AOI22X1 U540 ( .A(n295), .B(extratemp[3]), .C(DATA_IN[3]), .D(n292), .Y(
        n1294) );
  AOI22X1 U542 ( .A(n295), .B(extratemp[4]), .C(DATA_IN[4]), .D(n292), .Y(
        n1293) );
  AOI22X1 U544 ( .A(n295), .B(extratemp[5]), .C(DATA_IN[5]), .D(n292), .Y(
        n1292) );
  AOI22X1 U546 ( .A(n295), .B(extratemp[6]), .C(DATA_IN[6]), .D(n292), .Y(
        n1291) );
  AOI22X1 U548 ( .A(n295), .B(extratemp[7]), .C(DATA_IN[7]), .D(n292), .Y(
        n1290) );
  NAND3X1 U550 ( .A(n1504), .B(n247), .C(n1289), .Y(n1297) );
  NOR2X1 U551 ( .A(n1288), .B(n1577), .Y(n1289) );
  NAND3X1 U552 ( .A(n498), .B(n545), .C(n1432), .Y(n1577) );
  NAND2X1 U553 ( .A(n610), .B(n1501), .Y(n1504) );
  OAI22X1 U555 ( .A(n441), .B(n932), .C(n1286), .D(n959), .Y(n1021) );
  OAI22X1 U556 ( .A(n441), .B(n369), .C(n1286), .D(n259), .Y(n1020) );
  OAI22X1 U557 ( .A(n441), .B(n933), .C(n1286), .D(n953), .Y(n1019) );
  NOR2X1 U559 ( .A(n1285), .B(n1391), .Y(n1286) );
  OAI21X1 U560 ( .A(n240), .B(n938), .C(n1284), .Y(n1018) );
  NAND2X1 U561 ( .A(N519), .B(n1283), .Y(n1284) );
  OAI21X1 U563 ( .A(n240), .B(n945), .C(n1282), .Y(n1017) );
  NAND2X1 U564 ( .A(N518), .B(n1283), .Y(n1282) );
  OAI21X1 U566 ( .A(n240), .B(n944), .C(n1281), .Y(n1016) );
  NAND2X1 U567 ( .A(N517), .B(n1283), .Y(n1281) );
  OAI21X1 U569 ( .A(n240), .B(n943), .C(n1280), .Y(n1015) );
  NAND2X1 U570 ( .A(N516), .B(n1283), .Y(n1280) );
  OAI21X1 U572 ( .A(n240), .B(n942), .C(n1279), .Y(n1014) );
  NAND2X1 U573 ( .A(N515), .B(n1283), .Y(n1279) );
  OAI21X1 U575 ( .A(n240), .B(n941), .C(n1278), .Y(n1013) );
  NAND2X1 U576 ( .A(N514), .B(n1283), .Y(n1278) );
  OAI21X1 U578 ( .A(n240), .B(n940), .C(n1277), .Y(n1012) );
  NAND2X1 U579 ( .A(N513), .B(n1283), .Y(n1277) );
  OAI21X1 U581 ( .A(n240), .B(n939), .C(n1276), .Y(n1011) );
  NAND2X1 U582 ( .A(N512), .B(n1283), .Y(n1276) );
  NOR2X1 U583 ( .A(n1492), .B(n1275), .Y(n1283) );
  NAND3X1 U586 ( .A(n1274), .B(n551), .C(n1273), .Y(n1275) );
  NOR2X1 U587 ( .A(n326), .B(n616), .Y(n1273) );
  AOI22X1 U589 ( .A(n290), .B(inti[7]), .C(N503), .D(n255), .Y(n1272) );
  AOI22X1 U591 ( .A(n290), .B(inti[6]), .C(N502), .D(n255), .Y(n1269) );
  AOI22X1 U593 ( .A(n290), .B(inti[5]), .C(N501), .D(n255), .Y(n1268) );
  AOI22X1 U595 ( .A(n290), .B(inti[4]), .C(N500), .D(n255), .Y(n1267) );
  AOI22X1 U597 ( .A(n290), .B(inti[3]), .C(N499), .D(n253), .Y(n1266) );
  AOI22X1 U599 ( .A(n290), .B(inti[2]), .C(N498), .D(n253), .Y(n1265) );
  AOI22X1 U601 ( .A(n290), .B(inti[1]), .C(N497), .D(n253), .Y(n1264) );
  AOI22X1 U603 ( .A(n290), .B(inti[0]), .C(N496), .D(n253), .Y(n1263) );
  NOR2X1 U604 ( .A(n290), .B(n249), .Y(n1270) );
  NAND3X1 U605 ( .A(n581), .B(n545), .C(n443), .Y(n1271) );
  OAI21X1 U606 ( .A(n419), .B(n256), .C(n1262), .Y(n1010) );
  NAND2X1 U607 ( .A(N480), .B(n616), .Y(n1262) );
  OAI21X1 U609 ( .A(n419), .B(n952), .C(n1261), .Y(n1009) );
  NAND2X1 U610 ( .A(N481), .B(n616), .Y(n1261) );
  OAI21X1 U612 ( .A(n419), .B(n951), .C(n1260), .Y(n1008) );
  NAND2X1 U613 ( .A(N482), .B(n616), .Y(n1260) );
  OAI21X1 U615 ( .A(n419), .B(n950), .C(n1259), .Y(n1007) );
  NAND2X1 U616 ( .A(N483), .B(n616), .Y(n1259) );
  OAI21X1 U618 ( .A(n419), .B(n949), .C(n1258), .Y(n1006) );
  NAND2X1 U619 ( .A(N484), .B(n616), .Y(n1258) );
  OAI21X1 U621 ( .A(n419), .B(n948), .C(n1257), .Y(n1005) );
  NAND2X1 U622 ( .A(N485), .B(n616), .Y(n1257) );
  OAI21X1 U624 ( .A(n419), .B(n947), .C(n1256), .Y(n1004) );
  NAND2X1 U625 ( .A(N486), .B(n616), .Y(n1256) );
  NAND2X1 U628 ( .A(N487), .B(n616), .Y(n1255) );
  NAND3X1 U631 ( .A(n551), .B(n1492), .C(n1274), .Y(n1254) );
  NOR2X1 U632 ( .A(n1253), .B(n1252), .Y(n1274) );
  NAND3X1 U633 ( .A(n1432), .B(n581), .C(n447), .Y(n1252) );
  NAND3X1 U634 ( .A(n612), .B(n545), .C(n1251), .Y(n1253) );
  OAI21X1 U637 ( .A(n581), .B(n1249), .C(n1248), .Y(n1002) );
  OAI21X1 U638 ( .A(n1247), .B(n1285), .C(permuteComplete), .Y(n1248) );
  NAND2X1 U639 ( .A(n1246), .B(n439), .Y(n1249) );
  NAND3X1 U641 ( .A(n543), .B(n249), .C(n443), .Y(n1285) );
  NAND3X1 U643 ( .A(n285), .B(n341), .C(n447), .Y(n1245) );
  OAI21X1 U646 ( .A(n445), .B(n937), .C(n1244), .Y(n1001) );
  NAND2X1 U647 ( .A(N431), .B(n1243), .Y(n1244) );
  OAI21X1 U649 ( .A(n445), .B(n936), .C(n1242), .Y(n1000) );
  NAND2X1 U650 ( .A(N430), .B(n1243), .Y(n1242) );
  OAI21X1 U652 ( .A(n445), .B(n935), .C(n1241), .Y(n999) );
  NAND2X1 U653 ( .A(N429), .B(n1243), .Y(n1241) );
  OAI21X1 U654 ( .A(n445), .B(n934), .C(n1240), .Y(n998) );
  NAND2X1 U655 ( .A(N428), .B(n1243), .Y(n1240) );
  OAI21X1 U656 ( .A(n445), .B(n367), .C(n1239), .Y(n997) );
  NAND2X1 U657 ( .A(N427), .B(n1243), .Y(n1239) );
  OAI21X1 U659 ( .A(n445), .B(n933), .C(n1238), .Y(n996) );
  NAND2X1 U660 ( .A(N426), .B(n1243), .Y(n1238) );
  OAI21X1 U662 ( .A(n445), .B(n369), .C(n1237), .Y(n995) );
  NAND2X1 U663 ( .A(N425), .B(n1243), .Y(n1237) );
  OAI21X1 U664 ( .A(n445), .B(n932), .C(n1236), .Y(n994) );
  NAND2X1 U665 ( .A(N424), .B(n1243), .Y(n1236) );
  NOR2X1 U666 ( .A(n581), .B(n1246), .Y(n1243) );
  NOR2X1 U667 ( .A(n1235), .B(n1234), .Y(n1246) );
  NAND3X1 U668 ( .A(si[7]), .B(si[6]), .C(n1233), .Y(n1234) );
  NOR2X1 U669 ( .A(n934), .B(n935), .Y(n1233) );
  NAND3X1 U672 ( .A(si[3]), .B(si[2]), .C(n1232), .Y(n1235) );
  NOR2X1 U673 ( .A(n932), .B(n369), .Y(n1232) );
  NAND3X1 U677 ( .A(n447), .B(n285), .C(n1230), .Y(n1231) );
  NOR2X1 U678 ( .A(n268), .B(n1391), .Y(n1230) );
  NOR2X1 U679 ( .A(n1453), .B(n1519), .Y(n1391) );
  OAI21X1 U681 ( .A(n252), .B(n1287), .C(n549), .Y(n1229) );
  NAND3X1 U684 ( .A(n1515), .B(n1300), .C(n1226), .Y(n1227) );
  NOR2X1 U685 ( .A(n1225), .B(n1224), .Y(n1226) );
  OAI21X1 U686 ( .A(n252), .B(n220), .C(n1503), .Y(n1224) );
  OAI21X1 U690 ( .A(n1524), .B(n34), .C(n44), .Y(n1571) );
  OAI21X1 U693 ( .A(n488), .B(n923), .C(n1220), .Y(n993) );
  NAND2X1 U694 ( .A(N413), .B(n1219), .Y(n1220) );
  OAI21X1 U696 ( .A(n488), .B(n922), .C(n1218), .Y(n992) );
  NAND2X1 U697 ( .A(N412), .B(n1219), .Y(n1218) );
  OAI21X1 U699 ( .A(n488), .B(n921), .C(n1217), .Y(n991) );
  NAND2X1 U700 ( .A(N411), .B(n1219), .Y(n1217) );
  OAI21X1 U702 ( .A(n488), .B(n920), .C(n1216), .Y(n990) );
  NAND2X1 U703 ( .A(N410), .B(n1219), .Y(n1216) );
  OAI21X1 U705 ( .A(n488), .B(n919), .C(n1215), .Y(n989) );
  NAND2X1 U706 ( .A(N409), .B(n1219), .Y(n1215) );
  OAI21X1 U708 ( .A(n488), .B(n918), .C(n1214), .Y(n988) );
  NAND2X1 U709 ( .A(N408), .B(n1219), .Y(n1214) );
  OAI21X1 U711 ( .A(n488), .B(n917), .C(n1213), .Y(n987) );
  NAND2X1 U712 ( .A(N414), .B(n1219), .Y(n1213) );
  OAI21X1 U714 ( .A(n488), .B(n413), .C(n1212), .Y(n986) );
  NAND2X1 U715 ( .A(N407), .B(n1219), .Y(n1212) );
  NOR2X1 U716 ( .A(n1315), .B(n247), .Y(n1219) );
  NAND3X1 U721 ( .A(n498), .B(n1457), .C(n1211), .Y(n1315) );
  NOR2X1 U722 ( .A(n216), .B(n1288), .Y(n1211) );
  NAND3X1 U723 ( .A(n270), .B(n612), .C(n1210), .Y(n1288) );
  NOR2X1 U724 ( .A(n326), .B(n271), .Y(n1210) );
  NOR2X1 U727 ( .A(n1519), .B(n1287), .Y(n1475) );
  NOR2X1 U732 ( .A(n1467), .B(n1525), .Y(n1484) );
  OAI21X1 U733 ( .A(n1519), .B(n1208), .C(n524), .Y(n1299) );
  OAI21X1 U735 ( .A(n1476), .B(n626), .C(n592), .Y(n1207) );
  NOR2X1 U737 ( .A(n1524), .B(n626), .Y(n1494) );
  NAND3X1 U738 ( .A(n1206), .B(n624), .C(n614), .Y(n1457) );
  XOR2X1 U739 ( .A(n42), .B(n252), .Y(n1206) );
  NAND3X1 U741 ( .A(n1304), .B(n1431), .C(n518), .Y(n1435) );
  NAND2X1 U743 ( .A(n1301), .B(n540), .Y(n1438) );
  OAI21X1 U745 ( .A(n1524), .B(n34), .C(n1223), .Y(n1205) );
  NAND2X1 U746 ( .A(n629), .B(n541), .Y(n1223) );
  NOR2X1 U748 ( .A(n1225), .B(n268), .Y(n1301) );
  OAI21X1 U750 ( .A(n1525), .B(n1524), .C(n1204), .Y(n1225) );
  NOR2X1 U751 ( .A(n618), .B(n1518), .Y(n1204) );
  NOR2X1 U752 ( .A(n1467), .B(n1519), .Y(n1518) );
  NAND2X1 U754 ( .A(n39), .B(n42), .Y(n1456) );
  NOR2X1 U755 ( .A(n1390), .B(n553), .Y(n1431) );
  NOR2X1 U757 ( .A(n37), .B(n605), .Y(n1503) );
  NAND3X1 U759 ( .A(n1501), .B(n614), .C(n42), .Y(n1203) );
  NOR2X1 U760 ( .A(n1209), .B(n626), .Y(n1416) );
  OAI21X1 U762 ( .A(n220), .B(n1525), .C(n581), .Y(n1202) );
  NOR2X1 U764 ( .A(n1524), .B(n1519), .Y(n1247) );
  NAND2X1 U765 ( .A(n600), .B(n630), .Y(n1524) );
  NAND2X1 U766 ( .A(state[0]), .B(n547), .Y(n1476) );
  NAND2X1 U767 ( .A(n542), .B(n514), .Y(n1502) );
  AOI21X1 U769 ( .A(n1467), .B(n1208), .C(n626), .Y(n1488) );
  NOR2X1 U771 ( .A(n636), .B(state[2]), .Y(n1501) );
  NAND3X1 U772 ( .A(n42), .B(n579), .C(state[0]), .Y(n1467) );
  NAND2X1 U774 ( .A(n543), .B(n1221), .Y(n1487) );
  NAND2X1 U778 ( .A(n547), .B(n632), .Y(n1453) );
  NAND2X1 U780 ( .A(n579), .B(n630), .Y(n1495) );
  NOR2X1 U781 ( .A(n1228), .B(n616), .Y(n1304) );
  NAND2X1 U783 ( .A(n39), .B(n630), .Y(n1455) );
  NOR2X1 U784 ( .A(n1525), .B(n1520), .Y(n1568) );
  NAND3X1 U785 ( .A(n1492), .B(n1250), .C(n551), .Y(n1228) );
  NOR2X1 U787 ( .A(n1519), .B(n1209), .Y(n1450) );
  NAND3X1 U788 ( .A(n632), .B(n579), .C(n42), .Y(n1209) );
  NAND2X1 U790 ( .A(n624), .B(n636), .Y(n1519) );
  NAND2X1 U792 ( .A(n594), .B(n629), .Y(n1250) );
  NAND2X1 U794 ( .A(state[2]), .B(n636), .Y(n1525) );
  NAND2X1 U797 ( .A(n600), .B(n42), .Y(n1208) );
  NAND2X1 U799 ( .A(state[0]), .B(state[1]), .Y(n1491) );
  NAND2X1 U801 ( .A(n614), .B(n630), .Y(n1287) );
  NAND2X1 U804 ( .A(state[1]), .B(n632), .Y(n1520) );
  NAND2X1 U806 ( .A(state[2]), .B(n252), .Y(n1222) );
  NAND3X1 U807 ( .A(n1199), .B(n1201), .C(n1200), .Y(N479) );
  NOR2X1 U808 ( .A(n1198), .B(n1197), .Y(n1199) );
  OAI22X1 U809 ( .A(n865), .B(n1196), .C(n889), .D(n250), .Y(n1197) );
  OAI22X1 U812 ( .A(n777), .B(n1194), .C(n785), .D(n1193), .Y(n1198) );
  AOI22X1 U815 ( .A(n955), .B(\keyTable[5][0] ), .C(n954), .D(\keyTable[4][0] ), .Y(n1200) );
  AOI22X1 U816 ( .A(n957), .B(\keyTable[7][0] ), .C(\keyTable[6][0] ), .D(n956), .Y(n1201) );
  NAND3X1 U817 ( .A(n1192), .B(n1191), .C(n1190), .Y(N478) );
  NOR2X1 U818 ( .A(n1189), .B(n1188), .Y(n1190) );
  OAI22X1 U819 ( .A(n866), .B(n1196), .C(n888), .D(n250), .Y(n1188) );
  OAI22X1 U822 ( .A(n778), .B(n1194), .C(n786), .D(n1193), .Y(n1189) );
  AOI22X1 U825 ( .A(n955), .B(\keyTable[5][1] ), .C(n954), .D(\keyTable[4][1] ), .Y(n1191) );
  AOI22X1 U826 ( .A(n957), .B(\keyTable[7][1] ), .C(n956), .D(\keyTable[6][1] ), .Y(n1192) );
  NAND3X1 U827 ( .A(n1187), .B(n1186), .C(n1185), .Y(N477) );
  NOR2X1 U828 ( .A(n1184), .B(n1183), .Y(n1185) );
  OAI22X1 U829 ( .A(n867), .B(n1196), .C(n887), .D(n250), .Y(n1183) );
  OAI22X1 U832 ( .A(n779), .B(n1194), .C(n787), .D(n264), .Y(n1184) );
  AOI22X1 U835 ( .A(n955), .B(\keyTable[5][2] ), .C(n954), .D(\keyTable[4][2] ), .Y(n1186) );
  AOI22X1 U836 ( .A(n957), .B(\keyTable[7][2] ), .C(n956), .D(\keyTable[6][2] ), .Y(n1187) );
  NAND3X1 U837 ( .A(n1182), .B(n1181), .C(n1180), .Y(N476) );
  NOR2X1 U838 ( .A(n1179), .B(n1178), .Y(n1180) );
  OAI22X1 U839 ( .A(n868), .B(n1196), .C(n886), .D(n250), .Y(n1178) );
  OAI22X1 U842 ( .A(n780), .B(n1194), .C(n788), .D(n264), .Y(n1179) );
  AOI22X1 U845 ( .A(n955), .B(\keyTable[5][3] ), .C(n954), .D(\keyTable[4][3] ), .Y(n1181) );
  AOI22X1 U846 ( .A(n957), .B(\keyTable[7][3] ), .C(n956), .D(\keyTable[6][3] ), .Y(n1182) );
  NAND3X1 U847 ( .A(n1177), .B(n1176), .C(n1175), .Y(N475) );
  NOR2X1 U848 ( .A(n1174), .B(n1173), .Y(n1175) );
  OAI22X1 U849 ( .A(n869), .B(n1196), .C(n885), .D(n250), .Y(n1173) );
  OAI22X1 U852 ( .A(n781), .B(n1194), .C(n789), .D(n264), .Y(n1174) );
  AOI22X1 U855 ( .A(n955), .B(\keyTable[5][4] ), .C(n954), .D(\keyTable[4][4] ), .Y(n1176) );
  AOI22X1 U856 ( .A(n957), .B(\keyTable[7][4] ), .C(n956), .D(\keyTable[6][4] ), .Y(n1177) );
  NAND3X1 U857 ( .A(n1172), .B(n1171), .C(n1170), .Y(N474) );
  NOR2X1 U858 ( .A(n1169), .B(n1168), .Y(n1170) );
  OAI22X1 U859 ( .A(n870), .B(n1196), .C(n884), .D(n250), .Y(n1168) );
  OAI22X1 U862 ( .A(n782), .B(n1194), .C(n790), .D(n264), .Y(n1169) );
  AOI22X1 U865 ( .A(n955), .B(\keyTable[5][5] ), .C(n954), .D(\keyTable[4][5] ), .Y(n1171) );
  AOI22X1 U866 ( .A(n957), .B(\keyTable[7][5] ), .C(n956), .D(\keyTable[6][5] ), .Y(n1172) );
  NAND3X1 U867 ( .A(n1167), .B(n1166), .C(n1165), .Y(N473) );
  NOR2X1 U868 ( .A(n1164), .B(n1163), .Y(n1165) );
  OAI22X1 U869 ( .A(n871), .B(n1196), .C(n883), .D(n250), .Y(n1163) );
  OAI22X1 U872 ( .A(n783), .B(n1194), .C(n791), .D(n264), .Y(n1164) );
  AOI22X1 U875 ( .A(n955), .B(\keyTable[5][6] ), .C(n954), .D(\keyTable[4][6] ), .Y(n1166) );
  AOI22X1 U876 ( .A(n957), .B(\keyTable[7][6] ), .C(n956), .D(\keyTable[6][6] ), .Y(n1167) );
  NAND3X1 U877 ( .A(n1162), .B(n1161), .C(n1160), .Y(N472) );
  NOR2X1 U878 ( .A(n1159), .B(n1158), .Y(n1160) );
  OAI22X1 U879 ( .A(n890), .B(n1196), .C(n916), .D(n250), .Y(n1158) );
  NAND3X1 U880 ( .A(n953), .B(n958), .C(n959), .Y(n1195) );
  NAND3X1 U882 ( .A(n958), .B(keyi[0]), .C(n953), .Y(n1196) );
  OAI22X1 U884 ( .A(n784), .B(n1194), .C(n864), .D(n264), .Y(n1159) );
  NAND3X1 U885 ( .A(n959), .B(n953), .C(n265), .Y(n1193) );
  NAND3X1 U887 ( .A(keyi[1]), .B(keyi[0]), .C(n953), .Y(n1194) );
  AOI22X1 U890 ( .A(n955), .B(\keyTable[5][7] ), .C(n954), .D(\keyTable[4][7] ), .Y(n1161) );
  NAND3X1 U892 ( .A(n959), .B(n259), .C(n261), .Y(n1157) );
  NAND3X1 U894 ( .A(n259), .B(n258), .C(n261), .Y(n1156) );
  AOI22X1 U896 ( .A(n957), .B(\keyTable[7][7] ), .C(n956), .D(\keyTable[6][7] ), .Y(n1162) );
  NAND3X1 U898 ( .A(keyi[1]), .B(n959), .C(n261), .Y(n1155) );
  NAND3X1 U901 ( .A(n265), .B(n258), .C(n261), .Y(n1154) );
  OR2X2 U105 ( .A(n1517), .B(n1516), .Y(nextState[4]) );
  OR2X2 U134 ( .A(n1484), .B(n605), .Y(n1480) );
  AND2X2 U142 ( .A(n1509), .B(n1465), .Y(n1485) );
  AND2X2 U524 ( .A(n1484), .B(n500), .Y(n1313) );
  AND2X2 U635 ( .A(n249), .B(n1250), .Y(n1251) );
  AND2X2 U692 ( .A(n1221), .B(n514), .Y(n1515) );
  OR2X2 U761 ( .A(n1502), .B(n1202), .Y(n1390) );
  OR2X2 U775 ( .A(n34), .B(n1209), .Y(n1221) );
  OR2X2 U800 ( .A(n34), .B(n1287), .Y(n1492) );
  KSA_0_DW01_add_0 add_377 ( .A(temp), .B(extratemp), .CI(1'b0), .SUM({N527, 
        N526, N525, N524, N523, N522, N521, N520}) );
  KSA_0_DW01_add_1 add_337 ( .A(intj), .B(DATA_IN), .CI(1'b0), .SUM({N519, 
        N518, N517, N516, N515, N514, N513, N512}) );
  KSA_0_DW01_inc_0 add_289 ( .A(si), .SUM({N431, N430, N429, N428, N427, N426, 
        N425, N424}) );
  KSA_0_DW01_inc_1 add_263 ( .A(prefillCounter), .SUM({N414, N413, N412, N411, 
        N410, N409, N408, N407}) );
  KSA_0_DW01_inc_2 r126 ( .A(inti), .SUM({N503, N502, N501, N500, N499, N498, 
        N497, N496}) );
  KSA_0_DW01_add_3 add_1_root_add_0_root_add_302_2 ( .A(DATA_IN), .B(sj), .CI(
        1'b0), .SUM({N456, N455, N454, N453, N452, N451, N450, N449}) );
  KSA_0_DW01_add_2 add_0_root_add_0_root_add_302_2 ( .A({N472, N473, N474, 
        N475, N476, N477, N478, N479}), .B({N456, N455, N454, N453, N452, N451, 
        N450, N449}), .CI(1'b0), .SUM({N487, N486, N485, N484, N483, N482, 
        N481, N480}) );
  TBUFX1 \nfaddr_tri[5]  ( .A(n1143), .EN(n285), .Y(nfaddr[5]) );
  TBUFX1 \nfaddr_tri[0]  ( .A(n1138), .EN(n285), .Y(nfaddr[0]) );
  TBUFX1 \nfaddr_tri[1]  ( .A(n1139), .EN(n285), .Y(nfaddr[1]) );
  TBUFX1 \nfaddr_tri[2]  ( .A(n1140), .EN(n285), .Y(nfaddr[2]) );
  TBUFX1 \nfaddr_tri[3]  ( .A(n1141), .EN(n285), .Y(nfaddr[3]) );
  TBUFX1 \nfaddr_tri[4]  ( .A(n1142), .EN(n285), .Y(nfaddr[4]) );
  TBUFX1 \nfaddr_tri[6]  ( .A(n1144), .EN(n285), .Y(nfaddr[6]) );
  TBUFX1 \nfaddr_tri[7]  ( .A(n1145), .EN(n285), .Y(nfaddr[7]) );
  TBUFX1 \nfdata_tri[0]  ( .A(n1146), .EN(n612), .Y(nfdata[0]) );
  TBUFX1 \nfdata_tri[1]  ( .A(n1147), .EN(n612), .Y(nfdata[1]) );
  TBUFX1 \nfdata_tri[2]  ( .A(n1148), .EN(n612), .Y(nfdata[2]) );
  TBUFX1 \nfdata_tri[3]  ( .A(n1149), .EN(n612), .Y(nfdata[3]) );
  TBUFX1 \nfdata_tri[4]  ( .A(n1150), .EN(n612), .Y(nfdata[4]) );
  TBUFX1 \nfdata_tri[5]  ( .A(n1151), .EN(n612), .Y(nfdata[5]) );
  TBUFX1 \nfdata_tri[6]  ( .A(n1152), .EN(n612), .Y(nfdata[6]) );
  TBUFX1 \nfdata_tri[7]  ( .A(n1153), .EN(n612), .Y(nfdata[7]) );
  DFFSR PDATA_READY_reg ( .D(n553), .CLK(CLK), .R(n307), .S(1'b1), .Q(
        PDATA_READY) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n307), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[3]  ( .D(nextState[3]), .CLK(CLK), .R(n307), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[4]  ( .D(nextState[4]), .CLK(CLK), .R(n307), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n307), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n307), .S(1'b1), .Q(
        state[0]) );
  DFFSR \si_reg[7]  ( .D(n1001), .CLK(CLK), .R(n307), .S(1'b1), .Q(si[7]) );
  DFFSR \si_reg[6]  ( .D(n1000), .CLK(CLK), .R(n307), .S(1'b1), .Q(si[6]) );
  DFFSR \si_reg[5]  ( .D(n999), .CLK(CLK), .R(n307), .S(1'b1), .Q(si[5]) );
  DFFSR \si_reg[4]  ( .D(n998), .CLK(CLK), .R(n307), .S(1'b1), .Q(si[4]) );
  DFFSR \si_reg[3]  ( .D(n997), .CLK(CLK), .R(n307), .S(1'b1), .Q(si[3]) );
  DFFSR \si_reg[2]  ( .D(n996), .CLK(CLK), .R(n307), .S(1'b1), .Q(si[2]) );
  DFFSR \si_reg[1]  ( .D(n995), .CLK(CLK), .R(n307), .S(1'b1), .Q(si[1]) );
  DFFSR \si_reg[0]  ( .D(n994), .CLK(CLK), .R(n307), .S(1'b1), .Q(si[0]) );
  DFFSR \currentProcessedData_reg[7]  ( .D(nextProcessedData[7]), .CLK(CLK), 
        .R(n307), .S(1'b1), .Q(currentProcessedData[7]) );
  DFFSR \currentProcessedData_reg[6]  ( .D(nextProcessedData[6]), .CLK(CLK), 
        .R(n307), .S(1'b1), .Q(currentProcessedData[6]) );
  DFFSR \currentProcessedData_reg[5]  ( .D(nextProcessedData[5]), .CLK(CLK), 
        .R(n307), .S(1'b1), .Q(currentProcessedData[5]) );
  DFFSR \currentProcessedData_reg[4]  ( .D(nextProcessedData[4]), .CLK(CLK), 
        .R(n307), .S(1'b1), .Q(currentProcessedData[4]) );
  DFFSR \currentProcessedData_reg[3]  ( .D(nextProcessedData[3]), .CLK(CLK), 
        .R(n307), .S(1'b1), .Q(currentProcessedData[3]) );
  DFFSR \currentProcessedData_reg[2]  ( .D(nextProcessedData[2]), .CLK(CLK), 
        .R(n307), .S(1'b1), .Q(currentProcessedData[2]) );
  DFFSR \currentProcessedData_reg[1]  ( .D(nextProcessedData[1]), .CLK(CLK), 
        .R(n307), .S(1'b1), .Q(currentProcessedData[1]) );
  DFFSR \currentProcessedData_reg[0]  ( .D(nextProcessedData[0]), .CLK(CLK), 
        .R(n307), .S(1'b1), .Q(currentProcessedData[0]) );
  DFFSR \sj_reg[5]  ( .D(n1005), .CLK(CLK), .R(n307), .S(1'b1), .Q(sj[5]) );
  DFFSR \sj_reg[4]  ( .D(n1006), .CLK(CLK), .R(n307), .S(1'b1), .Q(sj[4]) );
  DFFSR \sj_reg[3]  ( .D(n1007), .CLK(CLK), .R(n307), .S(1'b1), .Q(sj[3]) );
  DFFSR \sj_reg[2]  ( .D(n1008), .CLK(CLK), .R(n307), .S(1'b1), .Q(sj[2]) );
  DFFSR \sj_reg[1]  ( .D(n1009), .CLK(CLK), .R(n307), .S(1'b1), .Q(sj[1]) );
  DFFSR \sj_reg[0]  ( .D(n1010), .CLK(CLK), .R(n307), .S(1'b1), .Q(sj[0]) );
  DFFSR \sj_reg[6]  ( .D(n1004), .CLK(CLK), .R(n307), .S(1'b1), .Q(sj[6]) );
  DFFSR \sj_reg[7]  ( .D(n1003), .CLK(CLK), .R(n307), .S(1'b1), .Q(sj[7]) );
  BUFX4 U4 ( .A(n1195), .Y(n250) );
  INVX4 U11 ( .A(n1157), .Y(n954) );
  BUFX2 U16 ( .A(n1380), .Y(n3) );
  BUFX2 U21 ( .A(n1380), .Y(n4) );
  BUFX2 U26 ( .A(n1380), .Y(n5) );
  BUFX2 U31 ( .A(n3), .Y(n6) );
  BUFX2 U36 ( .A(n3), .Y(n7) );
  BUFX2 U41 ( .A(n3), .Y(n8) );
  BUFX2 U45 ( .A(n3), .Y(n9) );
  BUFX2 U103 ( .A(n3), .Y(n10) );
  BUFX2 U107 ( .A(n4), .Y(n12) );
  BUFX2 U136 ( .A(n4), .Y(n14) );
  BUFX2 U141 ( .A(n4), .Y(n15) );
  BUFX2 U144 ( .A(n4), .Y(n16) );
  BUFX2 U155 ( .A(n4), .Y(n17) );
  BUFX2 U157 ( .A(n5), .Y(n20) );
  BUFX2 U190 ( .A(n5), .Y(n22) );
  BUFX2 U194 ( .A(n5), .Y(n24) );
  BUFX2 U198 ( .A(n5), .Y(n27) );
  BUFX2 U199 ( .A(n5), .Y(n29) );
  INVX4 U201 ( .A(n297), .Y(n300) );
  INVX2 U202 ( .A(n1222), .Y(n32) );
  INVX4 U204 ( .A(n32), .Y(n34) );
  BUFX2 U205 ( .A(n1416), .Y(n37) );
  BUFX4 U207 ( .A(state[3]), .Y(n252) );
  INVX2 U208 ( .A(n1155), .Y(n956) );
  BUFX2 U210 ( .A(state[4]), .Y(n42) );
  INVX2 U211 ( .A(n287), .Y(n290) );
  INVX2 U213 ( .A(n241), .Y(n302) );
  INVX2 U214 ( .A(n1305), .Y(n500) );
  INVX4 U216 ( .A(n1156), .Y(n955) );
  BUFX4 U217 ( .A(n1568), .Y(n39) );
  INVX2 U219 ( .A(n44), .Y(n271) );
  INVX1 U220 ( .A(sj[0]), .Y(n256) );
  INVX2 U224 ( .A(keyi[0]), .Y(n959) );
  INVX1 U225 ( .A(keyi[1]), .Y(n259) );
  OR2X2 U229 ( .A(n1525), .B(n1209), .Y(n44) );
  INVX2 U230 ( .A(n292), .Y(n295) );
  INVX2 U234 ( .A(n249), .Y(n268) );
  OR2X2 U235 ( .A(n34), .B(n1476), .Y(n249) );
  BUFX2 U239 ( .A(keyi[0]), .Y(n258) );
  AND2X2 U240 ( .A(n270), .B(n1223), .Y(n47) );
  INVX4 U244 ( .A(RST), .Y(n307) );
  OR2X2 U331 ( .A(n1299), .B(n1484), .Y(n216) );
  INVX2 U333 ( .A(n216), .Y(n1432) );
  INVX2 U335 ( .A(n42), .Y(n630) );
  INVX1 U337 ( .A(n1476), .Y(n218) );
  INVX2 U338 ( .A(n218), .Y(n220) );
  BUFX2 U341 ( .A(n244), .Y(n237) );
  INVX2 U344 ( .A(n1501), .Y(n626) );
  INVX2 U347 ( .A(n34), .Y(n230) );
  NOR2X1 U350 ( .A(n1495), .B(n235), .Y(n1511) );
  NAND2X1 U353 ( .A(n632), .B(n230), .Y(n235) );
  INVX1 U356 ( .A(n1503), .Y(n553) );
  INVX2 U359 ( .A(n238), .Y(n1300) );
  INVX2 U362 ( .A(n277), .Y(n280) );
  INVX1 U365 ( .A(state[2]), .Y(n624) );
  NAND3X1 U368 ( .A(n277), .B(n1457), .C(n47), .Y(n238) );
  INVX1 U371 ( .A(n47), .Y(n282) );
  NOR2X1 U374 ( .A(n1495), .B(n239), .Y(n1599) );
  NAND2X1 U377 ( .A(n632), .B(n1501), .Y(n239) );
  INVX2 U380 ( .A(n1275), .Y(n240) );
  INVX2 U383 ( .A(n1275), .Y(n421) );
  INVX2 U386 ( .A(n337), .Y(n317) );
  INVX2 U389 ( .A(n335), .Y(n318) );
  INVX2 U392 ( .A(n331), .Y(n327) );
  INVX2 U395 ( .A(n333), .Y(n326) );
  INVX2 U398 ( .A(n339), .Y(n311) );
  BUFX2 U401 ( .A(n345), .Y(n341) );
  BUFX2 U404 ( .A(n347), .Y(n339) );
  BUFX2 U407 ( .A(n329), .Y(n337) );
  BUFX2 U410 ( .A(n347), .Y(n335) );
  BUFX2 U413 ( .A(n329), .Y(n333) );
  BUFX2 U416 ( .A(n349), .Y(n331) );
  BUFX2 U419 ( .A(n349), .Y(n329) );
  BUFX2 U422 ( .A(n345), .Y(n343) );
  INVX2 U425 ( .A(n1475), .Y(n612) );
  AND2X2 U428 ( .A(n421), .B(n543), .Y(n241) );
  INVX2 U431 ( .A(n1271), .Y(n287) );
  NOR2X1 U434 ( .A(n1305), .B(n1304), .Y(n244) );
  INVX2 U502 ( .A(n1566), .Y(n297) );
  INVX2 U505 ( .A(n305), .Y(n347) );
  INVX2 U508 ( .A(n305), .Y(n345) );
  INVX2 U511 ( .A(n305), .Y(n349) );
  INVX1 U514 ( .A(n1193), .Y(n262) );
  INVX2 U517 ( .A(n1455), .Y(n616) );
  INVX2 U520 ( .A(n1254), .Y(n419) );
  INVX2 U523 ( .A(n1599), .Y(n270) );
  INVX2 U525 ( .A(n1297), .Y(n292) );
  INVX2 U526 ( .A(n247), .Y(n275) );
  INVX2 U531 ( .A(n246), .Y(n285) );
  INVX2 U533 ( .A(n307), .Y(n305) );
  INVX2 U535 ( .A(n1457), .Y(n604) );
  OR2X2 U537 ( .A(n216), .B(n1229), .Y(n246) );
  OR2X2 U539 ( .A(n220), .B(n1519), .Y(n247) );
  INVX2 U541 ( .A(n1571), .Y(n277) );
  INVX2 U543 ( .A(n1203), .Y(n605) );
  INVX2 U545 ( .A(keyi[1]), .Y(n958) );
  BUFX2 U547 ( .A(n1270), .Y(n253) );
  BUFX2 U549 ( .A(n1270), .Y(n255) );
  INVX2 U554 ( .A(keyi[2]), .Y(n953) );
  BUFX2 U558 ( .A(keyi[2]), .Y(n261) );
  INVX2 U562 ( .A(n262), .Y(n264) );
  INVX4 U565 ( .A(n1154), .Y(n957) );
  BUFX2 U568 ( .A(keyi[1]), .Y(n265) );
  INVX1 U571 ( .A(n1315), .Y(n488) );
  INVX1 U574 ( .A(n1453), .Y(n541) );
  OR2X2 U577 ( .A(n419), .B(n946), .Y(n267) );
  NAND2X1 U580 ( .A(n267), .B(n1255), .Y(n1003) );
  NAND2X1 U584 ( .A(n369), .B(n932), .Y(n351) );
  OAI21X1 U585 ( .A(n932), .B(n369), .C(n351), .Y(N442) );
  NOR2X1 U588 ( .A(n351), .B(si[2]), .Y(n355) );
  AOI21X1 U590 ( .A(n351), .B(si[2]), .C(n355), .Y(n353) );
  NAND2X1 U592 ( .A(n355), .B(n367), .Y(n357) );
  OAI21X1 U594 ( .A(n355), .B(n367), .C(n357), .Y(N444) );
  NOR2X1 U596 ( .A(n357), .B(si[4]), .Y(n361) );
  AOI21X1 U598 ( .A(n357), .B(si[4]), .C(n361), .Y(n359) );
  NAND2X1 U600 ( .A(n361), .B(n935), .Y(n363) );
  OAI21X1 U602 ( .A(n361), .B(n935), .C(n363), .Y(N446) );
  XNOR2X1 U608 ( .A(si[6]), .B(n363), .Y(N447) );
  NOR2X1 U611 ( .A(si[6]), .B(n363), .Y(n365) );
  XOR2X1 U614 ( .A(si[7]), .B(n365), .Y(N448) );
  INVX2 U617 ( .A(si[3]), .Y(n367) );
  INVX2 U620 ( .A(si[1]), .Y(n369) );
  INVX2 U623 ( .A(n359), .Y(N445) );
  INVX2 U626 ( .A(n353), .Y(N443) );
  INVX2 U627 ( .A(KEY_ERROR), .Y(n371) );
  INVX2 U629 ( .A(BYTE_READY), .Y(n373) );
  INVX2 U630 ( .A(n1509), .Y(n375) );
  INVX2 U636 ( .A(OPCODE[1]), .Y(n377) );
  INVX2 U640 ( .A(OPCODE[0]), .Y(n379) );
  INVX2 U642 ( .A(nextProcessedData[7]), .Y(n381) );
  INVX2 U644 ( .A(n1388), .Y(n383) );
  INVX2 U645 ( .A(nextProcessedData[6]), .Y(n385) );
  INVX2 U648 ( .A(n1381), .Y(n387) );
  INVX2 U651 ( .A(nextProcessedData[5]), .Y(n389) );
  INVX2 U658 ( .A(n1382), .Y(n391) );
  INVX2 U661 ( .A(nextProcessedData[4]), .Y(n393) );
  INVX2 U670 ( .A(n1383), .Y(n395) );
  INVX2 U671 ( .A(nextProcessedData[3]), .Y(n397) );
  INVX2 U674 ( .A(n1384), .Y(n399) );
  INVX2 U675 ( .A(nextProcessedData[2]), .Y(n401) );
  INVX2 U676 ( .A(n1385), .Y(n403) );
  INVX2 U680 ( .A(nextProcessedData[1]), .Y(n405) );
  INVX2 U682 ( .A(n1386), .Y(n407) );
  INVX2 U683 ( .A(nextProcessedData[0]), .Y(n409) );
  INVX2 U687 ( .A(n1387), .Y(n411) );
  INVX2 U688 ( .A(prefillCounter[0]), .Y(n413) );
  INVX2 U689 ( .A(nfdata[0]), .Y(n415) );
  INVX2 U691 ( .A(nfaddr[0]), .Y(n417) );
  INVX2 U695 ( .A(n1263), .Y(n423) );
  INVX2 U698 ( .A(n1264), .Y(n425) );
  INVX2 U701 ( .A(n1265), .Y(n427) );
  INVX2 U704 ( .A(n1266), .Y(n429) );
  INVX2 U707 ( .A(n1267), .Y(n431) );
  INVX2 U710 ( .A(n1268), .Y(n433) );
  INVX2 U713 ( .A(n1269), .Y(n435) );
  INVX2 U717 ( .A(n1272), .Y(n437) );
  INVX2 U718 ( .A(n1285), .Y(n439) );
  INVX2 U719 ( .A(n1286), .Y(n441) );
  INVX2 U720 ( .A(n1245), .Y(n443) );
  INVX2 U725 ( .A(n1231), .Y(n445) );
  INVX2 U726 ( .A(n1227), .Y(n447) );
  INVX2 U728 ( .A(nfdata[7]), .Y(n449) );
  INVX2 U729 ( .A(nfdata[6]), .Y(n451) );
  INVX2 U730 ( .A(nfdata[5]), .Y(n453) );
  INVX2 U731 ( .A(nfdata[4]), .Y(n455) );
  INVX2 U734 ( .A(nfdata[3]), .Y(n458) );
  INVX2 U736 ( .A(nfdata[2]), .Y(n459) );
  INVX2 U740 ( .A(nfdata[1]), .Y(n462) );
  INVX2 U742 ( .A(n1577), .Y(n463) );
  INVX2 U744 ( .A(n1298), .Y(n465) );
  INVX2 U747 ( .A(n1296), .Y(n467) );
  INVX2 U749 ( .A(n1295), .Y(n469) );
  INVX2 U753 ( .A(n1294), .Y(n471) );
  INVX2 U756 ( .A(n1293), .Y(n473) );
  INVX2 U758 ( .A(n1292), .Y(n475) );
  INVX2 U763 ( .A(n1291), .Y(n480) );
  INVX2 U768 ( .A(n1290), .Y(n482) );
  INVX2 U770 ( .A(n1435), .Y(n498) );
  INVX2 U773 ( .A(nfaddr[1]), .Y(n501) );
  INVX2 U776 ( .A(nfaddr[2]), .Y(n503) );
  INVX2 U777 ( .A(nfaddr[3]), .Y(n504) );
  INVX2 U779 ( .A(nfaddr[4]), .Y(n505) );
  INVX2 U782 ( .A(nfaddr[5]), .Y(n506) );
  INVX2 U786 ( .A(nfaddr[6]), .Y(n507) );
  INVX2 U789 ( .A(nfaddr[7]), .Y(n509) );
  INVX2 U791 ( .A(n1393), .Y(n512) );
  INVX2 U793 ( .A(n1488), .Y(n514) );
  INVX2 U795 ( .A(n1518), .Y(n516) );
  INVX2 U796 ( .A(n1438), .Y(n518) );
  INVX2 U798 ( .A(n1389), .Y(n520) );
  INVX2 U802 ( .A(n1299), .Y(n522) );
  INVX2 U803 ( .A(n1207), .Y(n524) );
  INVX2 U805 ( .A(n1434), .Y(n528) );
  INVX2 U810 ( .A(n1205), .Y(n540) );
  INVX2 U811 ( .A(n1487), .Y(n542) );
  INVX2 U813 ( .A(n1511), .Y(n543) );
  INVX2 U814 ( .A(n1391), .Y(n545) );
  INVX2 U820 ( .A(n1495), .Y(n547) );
  INVX2 U821 ( .A(n1228), .Y(n549) );
  INVX2 U823 ( .A(n1450), .Y(n551) );
  INVX2 U824 ( .A(n1579), .Y(n555) );
  INVX2 U830 ( .A(n1582), .Y(n557) );
  INVX2 U831 ( .A(n1585), .Y(n562) );
  INVX2 U833 ( .A(n1588), .Y(n569) );
  INVX2 U834 ( .A(n1591), .Y(n571) );
  INVX2 U840 ( .A(n1594), .Y(n572) );
  INVX2 U841 ( .A(n1597), .Y(n575) );
  INVX2 U843 ( .A(n1601), .Y(n577) );
  INVX2 U844 ( .A(state[1]), .Y(n579) );
  INVX2 U850 ( .A(n1247), .Y(n581) );
  INVX2 U851 ( .A(n1494), .Y(n592) );
  INVX2 U853 ( .A(n1208), .Y(n594) );
  INVX2 U854 ( .A(n1491), .Y(n600) );
  INVX2 U860 ( .A(n1523), .Y(n606) );
  INVX2 U861 ( .A(n1287), .Y(n610) );
  INVX2 U863 ( .A(n1520), .Y(n614) );
  INVX2 U864 ( .A(n1456), .Y(n618) );
  INVX2 U870 ( .A(n1525), .Y(n629) );
  INVX2 U871 ( .A(state[0]), .Y(n632) );
  INVX2 U873 ( .A(state[3]), .Y(n636) );
  INVX2 U874 ( .A(\keyTable[7][0] ), .Y(n637) );
  INVX2 U881 ( .A(\keyTable[7][1] ), .Y(n638) );
  INVX2 U883 ( .A(\keyTable[7][2] ), .Y(n648) );
  INVX2 U886 ( .A(\keyTable[7][3] ), .Y(n649) );
  INVX2 U888 ( .A(\keyTable[7][4] ), .Y(n650) );
  INVX2 U889 ( .A(\keyTable[7][5] ), .Y(n651) );
  INVX2 U891 ( .A(\keyTable[7][6] ), .Y(n692) );
  INVX2 U893 ( .A(\keyTable[7][7] ), .Y(n701) );
  INVX2 U895 ( .A(\keyTable[6][0] ), .Y(n746) );
  INVX2 U897 ( .A(\keyTable[6][1] ), .Y(n748) );
  INVX2 U899 ( .A(\keyTable[6][2] ), .Y(n750) );
  INVX2 U900 ( .A(\keyTable[6][3] ), .Y(n752) );
  INVX2 U902 ( .A(\keyTable[6][4] ), .Y(n754) );
  INVX2 U903 ( .A(\keyTable[6][5] ), .Y(n756) );
  INVX2 U904 ( .A(\keyTable[6][6] ), .Y(n758) );
  INVX2 U905 ( .A(\keyTable[6][7] ), .Y(n760) );
  INVX2 U906 ( .A(\keyTable[5][0] ), .Y(n761) );
  INVX2 U907 ( .A(\keyTable[5][1] ), .Y(n762) );
  INVX2 U908 ( .A(\keyTable[5][2] ), .Y(n763) );
  INVX2 U909 ( .A(\keyTable[5][3] ), .Y(n764) );
  INVX2 U910 ( .A(\keyTable[5][4] ), .Y(n765) );
  INVX2 U911 ( .A(\keyTable[5][5] ), .Y(n766) );
  INVX2 U912 ( .A(\keyTable[5][6] ), .Y(n767) );
  INVX2 U913 ( .A(\keyTable[5][7] ), .Y(n768) );
  INVX2 U914 ( .A(\keyTable[4][0] ), .Y(n769) );
  INVX2 U915 ( .A(\keyTable[4][1] ), .Y(n770) );
  INVX2 U916 ( .A(\keyTable[4][2] ), .Y(n771) );
  INVX2 U917 ( .A(\keyTable[4][3] ), .Y(n772) );
  INVX2 U918 ( .A(\keyTable[4][4] ), .Y(n773) );
  INVX2 U919 ( .A(\keyTable[4][5] ), .Y(n774) );
  INVX2 U920 ( .A(\keyTable[4][6] ), .Y(n775) );
  INVX2 U921 ( .A(\keyTable[4][7] ), .Y(n776) );
  INVX2 U922 ( .A(\keyTable[3][0] ), .Y(n777) );
  INVX2 U923 ( .A(\keyTable[3][1] ), .Y(n778) );
  INVX2 U924 ( .A(\keyTable[3][2] ), .Y(n779) );
  INVX2 U925 ( .A(\keyTable[3][3] ), .Y(n780) );
  INVX2 U926 ( .A(\keyTable[3][4] ), .Y(n781) );
  INVX2 U927 ( .A(\keyTable[3][5] ), .Y(n782) );
  INVX2 U928 ( .A(\keyTable[3][6] ), .Y(n783) );
  INVX2 U929 ( .A(\keyTable[3][7] ), .Y(n784) );
  INVX2 U930 ( .A(\keyTable[2][0] ), .Y(n785) );
  INVX2 U931 ( .A(\keyTable[2][1] ), .Y(n786) );
  INVX2 U932 ( .A(\keyTable[2][2] ), .Y(n787) );
  INVX2 U933 ( .A(\keyTable[2][3] ), .Y(n788) );
  INVX2 U934 ( .A(\keyTable[2][4] ), .Y(n789) );
  INVX2 U935 ( .A(\keyTable[2][5] ), .Y(n790) );
  INVX2 U936 ( .A(\keyTable[2][6] ), .Y(n791) );
  INVX2 U937 ( .A(\keyTable[2][7] ), .Y(n864) );
  INVX2 U938 ( .A(\keyTable[1][0] ), .Y(n865) );
  INVX2 U939 ( .A(\keyTable[1][1] ), .Y(n866) );
  INVX2 U940 ( .A(\keyTable[1][2] ), .Y(n867) );
  INVX2 U941 ( .A(\keyTable[1][3] ), .Y(n868) );
  INVX2 U942 ( .A(\keyTable[1][4] ), .Y(n869) );
  INVX2 U943 ( .A(\keyTable[1][5] ), .Y(n870) );
  INVX2 U944 ( .A(\keyTable[1][6] ), .Y(n871) );
  INVX2 U945 ( .A(\keyTable[0][6] ), .Y(n883) );
  INVX2 U946 ( .A(\keyTable[0][5] ), .Y(n884) );
  INVX2 U947 ( .A(\keyTable[0][4] ), .Y(n885) );
  INVX2 U948 ( .A(\keyTable[0][3] ), .Y(n886) );
  INVX2 U949 ( .A(\keyTable[0][2] ), .Y(n887) );
  INVX2 U950 ( .A(\keyTable[0][1] ), .Y(n888) );
  INVX2 U951 ( .A(\keyTable[0][0] ), .Y(n889) );
  INVX2 U952 ( .A(\keyTable[1][7] ), .Y(n890) );
  INVX2 U953 ( .A(\keyTable[0][7] ), .Y(n916) );
  INVX2 U954 ( .A(prefillCounter[7]), .Y(n917) );
  INVX2 U955 ( .A(prefillCounter[1]), .Y(n918) );
  INVX2 U956 ( .A(prefillCounter[2]), .Y(n919) );
  INVX2 U957 ( .A(prefillCounter[3]), .Y(n920) );
  INVX2 U958 ( .A(prefillCounter[4]), .Y(n921) );
  INVX2 U959 ( .A(prefillCounter[5]), .Y(n922) );
  INVX2 U960 ( .A(prefillCounter[6]), .Y(n923) );
  INVX2 U961 ( .A(temp[7]), .Y(n924) );
  INVX2 U962 ( .A(temp[0]), .Y(n925) );
  INVX2 U963 ( .A(temp[1]), .Y(n926) );
  INVX2 U964 ( .A(temp[2]), .Y(n927) );
  INVX2 U965 ( .A(temp[3]), .Y(n928) );
  INVX2 U966 ( .A(temp[4]), .Y(n929) );
  INVX2 U967 ( .A(temp[5]), .Y(n930) );
  INVX2 U968 ( .A(temp[6]), .Y(n931) );
  INVX2 U969 ( .A(si[0]), .Y(n932) );
  INVX2 U970 ( .A(si[2]), .Y(n933) );
  INVX2 U971 ( .A(si[4]), .Y(n934) );
  INVX2 U972 ( .A(si[5]), .Y(n935) );
  INVX2 U973 ( .A(si[6]), .Y(n936) );
  INVX2 U974 ( .A(si[7]), .Y(n937) );
  INVX2 U975 ( .A(intj[7]), .Y(n938) );
  INVX2 U976 ( .A(intj[0]), .Y(n939) );
  INVX2 U977 ( .A(intj[1]), .Y(n940) );
  INVX2 U978 ( .A(intj[2]), .Y(n941) );
  INVX2 U979 ( .A(intj[3]), .Y(n942) );
  INVX2 U980 ( .A(intj[4]), .Y(n943) );
  INVX2 U981 ( .A(intj[5]), .Y(n944) );
  INVX2 U982 ( .A(intj[6]), .Y(n945) );
  INVX2 U983 ( .A(sj[7]), .Y(n946) );
  INVX2 U984 ( .A(sj[6]), .Y(n947) );
  INVX2 U985 ( .A(sj[5]), .Y(n948) );
  INVX2 U986 ( .A(sj[4]), .Y(n949) );
  INVX2 U987 ( .A(sj[3]), .Y(n950) );
  INVX2 U988 ( .A(sj[2]), .Y(n951) );
  INVX2 U989 ( .A(sj[1]), .Y(n952) );
  INVX2 U990 ( .A(currentProcessedData[0]), .Y(n960) );
  INVX2 U991 ( .A(currentProcessedData[1]), .Y(n961) );
  INVX2 U992 ( .A(currentProcessedData[2]), .Y(n962) );
  INVX2 U993 ( .A(currentProcessedData[3]), .Y(n963) );
  INVX2 U994 ( .A(currentProcessedData[4]), .Y(n964) );
  INVX2 U995 ( .A(currentProcessedData[5]), .Y(n965) );
  INVX2 U996 ( .A(currentProcessedData[6]), .Y(n966) );
  INVX2 U997 ( .A(currentProcessedData[7]), .Y(n967) );
  INVX2 U998 ( .A(faddr[7]), .Y(n968) );
  INVX2 U999 ( .A(faddr[6]), .Y(n969) );
  INVX2 U1000 ( .A(faddr[5]), .Y(n970) );
  INVX2 U1001 ( .A(faddr[4]), .Y(n971) );
  INVX2 U1002 ( .A(faddr[3]), .Y(n972) );
  INVX2 U1003 ( .A(faddr[2]), .Y(n973) );
  INVX2 U1004 ( .A(faddr[1]), .Y(n974) );
  INVX2 U1005 ( .A(faddr[0]), .Y(n975) );
  INVX2 U1006 ( .A(fdata[7]), .Y(n976) );
  INVX2 U1007 ( .A(fdata[6]), .Y(n977) );
  INVX2 U1008 ( .A(fdata[5]), .Y(n978) );
  INVX2 U1009 ( .A(fdata[4]), .Y(n979) );
  INVX2 U1010 ( .A(fdata[3]), .Y(n980) );
  INVX2 U1011 ( .A(fdata[2]), .Y(n981) );
  INVX2 U1012 ( .A(fdata[1]), .Y(n982) );
  INVX2 U1013 ( .A(fdata[0]), .Y(n983) );
endmodule


module uart_edge_detector_0 ( CLK, RST, SERIAL_IN, START_BIT );
  input CLK, RST, SERIAL_IN;
  output START_BIT;
  wire   Q_int, Q_int2, n2, n4;

  DFFSR Q_int_reg ( .D(SERIAL_IN), .CLK(CLK), .R(n2), .S(1'b1), .Q(Q_int) );
  NOR2X1 U7 ( .A(Q_int), .B(n4), .Y(START_BIT) );
  DFFSR Q_int2_reg ( .D(Q_int), .CLK(CLK), .R(n2), .S(1'b1), .Q(Q_int2) );
  INVX2 U4 ( .A(RST), .Y(n2) );
  INVX2 U6 ( .A(Q_int2), .Y(n4) );
endmodule


module uart_error_0 ( RST, CLK, RBUF_FULL, CHK_ERROR, OE );
  input RST, CLK, RBUF_FULL, CHK_ERROR;
  output OE;
  wire   OE_prime, n2;

  AND2X2 U5 ( .A(RBUF_FULL), .B(CHK_ERROR), .Y(OE_prime) );
  DFFSR OE_reg ( .D(OE_prime), .CLK(CLK), .R(n2), .S(1'b1), .Q(OE) );
  INVX2 U4 ( .A(RST), .Y(n2) );
endmodule


module uart_rcu_0 ( CLK, RST, START_BIT, STOP_RCVING, SB_DETECT, RBUF_LOAD, 
        TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR );
  input CLK, RST, START_BIT, STOP_RCVING, SB_DETECT;
  output RBUF_LOAD, TIMER_TRIG, CHK_ERROR, SET_RBUF_FULL, SBC_EN, SBC_CLR;
  wire   timerRunning, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N99, \add_46/carry[7] , \add_46/carry[6] ,
         \add_46/carry[5] , \add_46/carry[4] , \add_46/carry[3] , n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113;
  wire   [2:0] state;
  wire   [7:0] count;
  wire   [7:0] nextCount;
  wire   [2:0] nextState;

  DFFSR \nextCount_reg[0]  ( .D(N31), .CLK(CLK), .R(1'b1), .S(n27), .Q(
        nextCount[0]) );
  AND2X2 U33 ( .A(N30), .B(timerRunning), .Y(N38) );
  AND2X2 U34 ( .A(N29), .B(timerRunning), .Y(N37) );
  AND2X2 U35 ( .A(N28), .B(timerRunning), .Y(N36) );
  AND2X2 U36 ( .A(N27), .B(timerRunning), .Y(N35) );
  AND2X2 U37 ( .A(N26), .B(timerRunning), .Y(N34) );
  AND2X2 U38 ( .A(N25), .B(timerRunning), .Y(N33) );
  AND2X2 U39 ( .A(N24), .B(timerRunning), .Y(N32) );
  OAI21X1 U54 ( .A(n112), .B(n43), .C(n111), .Y(n113) );
  OAI21X1 U55 ( .A(n44), .B(n42), .C(n43), .Y(n111) );
  NAND2X1 U56 ( .A(n110), .B(n109), .Y(n87) );
  OAI21X1 U57 ( .A(n108), .B(n107), .C(timerRunning), .Y(n109) );
  NAND2X1 U58 ( .A(n106), .B(n105), .Y(n107) );
  NAND2X1 U59 ( .A(n104), .B(n105), .Y(n86) );
  NAND3X1 U60 ( .A(n35), .B(n110), .C(CHK_ERROR), .Y(n104) );
  OAI21X1 U61 ( .A(n103), .B(n47), .C(n102), .Y(n85) );
  NAND2X1 U62 ( .A(n105), .B(n101), .Y(n103) );
  NAND2X1 U63 ( .A(n100), .B(n38), .Y(n105) );
  NAND3X1 U64 ( .A(n99), .B(n98), .C(n97), .Y(n84) );
  NAND3X1 U65 ( .A(n34), .B(n110), .C(SET_RBUF_FULL), .Y(n97) );
  NAND2X1 U66 ( .A(n101), .B(n98), .Y(n108) );
  NAND3X1 U67 ( .A(nextState[0]), .B(nextState[1]), .C(n100), .Y(n98) );
  NAND3X1 U68 ( .A(n36), .B(n38), .C(n100), .Y(n99) );
  OAI21X1 U69 ( .A(n96), .B(n45), .C(n110), .Y(n83) );
  OAI21X1 U70 ( .A(n96), .B(n46), .C(n110), .Y(n82) );
  NAND2X1 U71 ( .A(n101), .B(n102), .Y(n96) );
  NAND3X1 U72 ( .A(nextState[1]), .B(n36), .C(n39), .Y(n102) );
  NAND2X1 U73 ( .A(n95), .B(n106), .Y(n81) );
  NAND3X1 U74 ( .A(nextState[1]), .B(n36), .C(n100), .Y(n106) );
  NAND3X1 U75 ( .A(n101), .B(n110), .C(RBUF_LOAD), .Y(n95) );
  NAND3X1 U76 ( .A(nextState[0]), .B(n38), .C(n39), .Y(n110) );
  NAND3X1 U77 ( .A(n36), .B(n38), .C(n39), .Y(n101) );
  OAI21X1 U78 ( .A(n40), .B(n43), .C(n94), .Y(n100) );
  NAND3X1 U79 ( .A(state[0]), .B(n43), .C(state[1]), .Y(n94) );
  NAND2X1 U80 ( .A(n93), .B(n92), .Y(n112) );
  OAI21X1 U81 ( .A(n91), .B(n92), .C(n93), .Y(nextState[1]) );
  NOR2X1 U82 ( .A(N99), .B(state[2]), .Y(n91) );
  OAI21X1 U83 ( .A(state[2]), .B(n90), .C(n93), .Y(nextState[0]) );
  NAND2X1 U84 ( .A(state[1]), .B(n44), .Y(n93) );
  AOI21X1 U85 ( .A(START_BIT), .B(n44), .C(n89), .Y(n90) );
  OAI21X1 U86 ( .A(N99), .B(n92), .C(n88), .Y(n89) );
  NAND2X1 U87 ( .A(SB_DETECT), .B(state[1]), .Y(n88) );
  NAND2X1 U88 ( .A(state[0]), .B(n42), .Y(n92) );
  NAND2X1 U89 ( .A(n37), .B(timerRunning), .Y(N31) );
  DFFSR \count_reg[7]  ( .D(nextCount[7]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[7]) );
  DFFSR \count_reg[6]  ( .D(nextCount[6]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[6]) );
  DFFSR \count_reg[5]  ( .D(nextCount[5]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[5]) );
  DFFSR \count_reg[4]  ( .D(nextCount[4]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[4]) );
  DFFSR \count_reg[3]  ( .D(nextCount[3]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[3]) );
  DFFSR \count_reg[2]  ( .D(nextCount[2]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[1]  ( .D(nextCount[1]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[1]) );
  DFFSR \count_reg[0]  ( .D(nextCount[0]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        count[0]) );
  DFFSR \nextCount_reg[2]  ( .D(N33), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[2]) );
  DFFSR \nextCount_reg[1]  ( .D(N32), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[1]) );
  DFFSR \state_reg[2]  ( .D(n41), .CLK(CLK), .R(n27), .S(1'b1), .Q(state[2])
         );
  DFFSR \nextCount_reg[3]  ( .D(N34), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[3]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        state[1]) );
  DFFSR \nextCount_reg[4]  ( .D(N35), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[4]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        state[0]) );
  DFFSR \nextCount_reg[5]  ( .D(N36), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[5]) );
  DFFSR \nextCount_reg[6]  ( .D(N37), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[6]) );
  DFFSR RBUF_LOAD_reg ( .D(n81), .CLK(CLK), .R(n27), .S(1'b1), .Q(RBUF_LOAD)
         );
  DFFSR timerRunning_reg ( .D(n87), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        timerRunning) );
  DFFSR TIMER_TRIG_reg ( .D(n82), .CLK(CLK), .R(n27), .S(1'b1), .Q(TIMER_TRIG)
         );
  DFFSR SBC_CLR_reg ( .D(n83), .CLK(CLK), .R(n27), .S(1'b1), .Q(SBC_CLR) );
  DFFSR SBC_EN_reg ( .D(n85), .CLK(CLK), .R(n27), .S(1'b1), .Q(SBC_EN) );
  DFFSR \nextCount_reg[7]  ( .D(N38), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        nextCount[7]) );
  DFFSR SET_RBUF_FULL_reg ( .D(n84), .CLK(CLK), .R(n27), .S(1'b1), .Q(
        SET_RBUF_FULL) );
  DFFSR CHK_ERROR_reg ( .D(n86), .CLK(CLK), .R(n27), .S(1'b1), .Q(CHK_ERROR)
         );
  INVX4 U3 ( .A(RST), .Y(n27) );
  XOR2X1 U30 ( .A(count[7]), .B(\add_46/carry[7] ), .Y(N30) );
  AND2X1 U31 ( .A(count[6]), .B(\add_46/carry[6] ), .Y(\add_46/carry[7] ) );
  XOR2X1 U32 ( .A(\add_46/carry[6] ), .B(count[6]), .Y(N29) );
  AND2X1 U40 ( .A(count[5]), .B(\add_46/carry[5] ), .Y(\add_46/carry[6] ) );
  XOR2X1 U41 ( .A(\add_46/carry[5] ), .B(count[5]), .Y(N28) );
  AND2X1 U42 ( .A(count[4]), .B(\add_46/carry[4] ), .Y(\add_46/carry[5] ) );
  XOR2X1 U43 ( .A(\add_46/carry[4] ), .B(count[4]), .Y(N27) );
  AND2X1 U44 ( .A(count[3]), .B(\add_46/carry[3] ), .Y(\add_46/carry[4] ) );
  XOR2X1 U45 ( .A(\add_46/carry[3] ), .B(count[3]), .Y(N26) );
  AND2X1 U46 ( .A(count[2]), .B(count[1]), .Y(\add_46/carry[3] ) );
  XOR2X1 U47 ( .A(count[1]), .B(count[2]), .Y(N25) );
  INVX2 U48 ( .A(count[1]), .Y(N24) );
  OAI21X1 U49 ( .A(count[0]), .B(count[1]), .C(count[2]), .Y(n28) );
  NOR2X1 U50 ( .A(n33), .B(n28), .Y(n29) );
  OAI21X1 U51 ( .A(n29), .B(count[4]), .C(count[6]), .Y(n30) );
  OAI21X1 U52 ( .A(n32), .B(n30), .C(n31), .Y(N99) );
  INVX2 U53 ( .A(count[7]), .Y(n31) );
  INVX2 U90 ( .A(count[5]), .Y(n32) );
  INVX2 U91 ( .A(count[3]), .Y(n33) );
  INVX2 U92 ( .A(n108), .Y(n34) );
  INVX2 U93 ( .A(n103), .Y(n35) );
  INVX2 U94 ( .A(nextState[0]), .Y(n36) );
  INVX2 U95 ( .A(count[0]), .Y(n37) );
  INVX2 U96 ( .A(nextState[1]), .Y(n38) );
  INVX2 U97 ( .A(n100), .Y(n39) );
  INVX2 U98 ( .A(n112), .Y(n40) );
  INVX2 U99 ( .A(n113), .Y(n41) );
  INVX2 U100 ( .A(state[1]), .Y(n42) );
  INVX2 U101 ( .A(state[2]), .Y(n43) );
  INVX2 U102 ( .A(state[0]), .Y(n44) );
  INVX2 U103 ( .A(SBC_CLR), .Y(n45) );
  INVX2 U104 ( .A(TIMER_TRIG), .Y(n46) );
  INVX2 U105 ( .A(SBC_EN), .Y(n47) );
endmodule


module uart_rcv_buf_0 ( CLK, RST, LOAD_RBUF, LOAD_DATA, RCV_DATA );
  input [7:0] LOAD_DATA;
  output [7:0] RCV_DATA;
  input CLK, RST, LOAD_RBUF;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;

  AOI22X1 U3 ( .A(n17), .B(LOAD_DATA[0]), .C(RCV_DATA[0]), .D(n27), .Y(n35) );
  AOI22X1 U5 ( .A(LOAD_DATA[1]), .B(n17), .C(RCV_DATA[1]), .D(n27), .Y(n34) );
  AOI22X1 U7 ( .A(LOAD_DATA[2]), .B(n17), .C(RCV_DATA[2]), .D(n27), .Y(n33) );
  AOI22X1 U9 ( .A(LOAD_DATA[3]), .B(n17), .C(RCV_DATA[3]), .D(n27), .Y(n32) );
  AOI22X1 U11 ( .A(LOAD_DATA[4]), .B(n17), .C(RCV_DATA[4]), .D(n27), .Y(n31)
         );
  AOI22X1 U13 ( .A(LOAD_DATA[5]), .B(n17), .C(RCV_DATA[5]), .D(n27), .Y(n30)
         );
  AOI22X1 U15 ( .A(LOAD_DATA[6]), .B(n17), .C(RCV_DATA[6]), .D(n27), .Y(n29)
         );
  AOI22X1 U18 ( .A(LOAD_DATA[7]), .B(n17), .C(RCV_DATA[7]), .D(n27), .Y(n28)
         );
  DFFSR \Q_int_reg[0]  ( .D(n26), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[0]) );
  DFFSR \Q_int_reg[7]  ( .D(n19), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[7]) );
  DFFSR \Q_int_reg[6]  ( .D(n20), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[6]) );
  DFFSR \Q_int_reg[5]  ( .D(n21), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[5]) );
  DFFSR \Q_int_reg[4]  ( .D(n22), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[4]) );
  DFFSR \Q_int_reg[1]  ( .D(n25), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[1]) );
  DFFSR \Q_int_reg[2]  ( .D(n24), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[2]) );
  DFFSR \Q_int_reg[3]  ( .D(n23), .CLK(CLK), .R(n18), .S(1'b1), .Q(RCV_DATA[3]) );
  INVX2 U17 ( .A(RST), .Y(n18) );
  BUFX2 U19 ( .A(LOAD_RBUF), .Y(n17) );
  INVX2 U20 ( .A(n28), .Y(n19) );
  INVX2 U21 ( .A(n29), .Y(n20) );
  INVX2 U22 ( .A(n30), .Y(n21) );
  INVX2 U23 ( .A(n31), .Y(n22) );
  INVX2 U24 ( .A(n32), .Y(n23) );
  INVX2 U25 ( .A(n33), .Y(n24) );
  INVX2 U26 ( .A(n34), .Y(n25) );
  INVX2 U27 ( .A(n35), .Y(n26) );
  INVX2 U28 ( .A(n17), .Y(n27) );
endmodule


module uart_rcv_buf_full_0 ( CLK, RST, CLR_RBUF, SET_RBUF_FULL, RBUF_FULL );
  input CLK, RST, CLR_RBUF, SET_RBUF_FULL;
  output RBUF_FULL;
  wire   n4, n5;

  NOR2X1 U3 ( .A(RST), .B(CLR_RBUF), .Y(n5) );
  OR2X2 U4 ( .A(RBUF_FULL), .B(SET_RBUF_FULL), .Y(n4) );
  DFFSR Q_int_reg ( .D(n4), .CLK(CLK), .R(n5), .S(1'b1), .Q(RBUF_FULL) );
endmodule


module uart_sb_check_0 ( RST, CLK, SBC_CLR, SBC_EN, STOP_DATA, SB_DETECT, SBE
 );
  input [1:0] STOP_DATA;
  input RST, CLK, SBC_CLR, SBC_EN;
  output SB_DETECT, SBE;
  wire   SBE_prime, sb_detect_flag, n3, n4, n5, n6, n10, n11, n12;

  OR2X2 U6 ( .A(SBC_CLR), .B(STOP_DATA[0]), .Y(n12) );
  NOR2X1 U10 ( .A(n12), .B(n11), .Y(sb_detect_flag) );
  NAND2X1 U11 ( .A(STOP_DATA[1]), .B(SBC_EN), .Y(n11) );
  NOR2X1 U12 ( .A(n6), .B(n10), .Y(SBE_prime) );
  OAI21X1 U13 ( .A(STOP_DATA[0]), .B(n4), .C(n5), .Y(n10) );
  DFFSR SBE_reg ( .D(SBE_prime), .CLK(CLK), .R(n3), .S(1'b1), .Q(SBE) );
  DFFSR SB_DETECT_reg ( .D(sb_detect_flag), .CLK(CLK), .R(n3), .S(1'b1), .Q(
        SB_DETECT) );
  INVX2 U5 ( .A(RST), .Y(n3) );
  INVX2 U7 ( .A(STOP_DATA[1]), .Y(n4) );
  INVX2 U8 ( .A(SBC_CLR), .Y(n5) );
  INVX2 U9 ( .A(SBC_EN), .Y(n6) );
endmodule


module uart_sr_10bit_0 ( CLK, RST, SHIFT_STROBE, SERIAL_IN, LOAD_DATA, 
        STOP_DATA );
  output [7:0] LOAD_DATA;
  output [1:0] STOP_DATA;
  input CLK, RST, SHIFT_STROBE, SERIAL_IN;
  wire   n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, n32, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45;

  OAI21X1 U2 ( .A(n32), .B(n13), .C(n45), .Y(n43) );
  NAND2X1 U3 ( .A(LOAD_DATA[0]), .B(n13), .Y(n45) );
  OAI22X1 U4 ( .A(n13), .B(n31), .C(SHIFT_STROBE), .D(n32), .Y(n42) );
  OAI22X1 U6 ( .A(n13), .B(n29), .C(SHIFT_STROBE), .D(n31), .Y(n41) );
  OAI22X1 U8 ( .A(n13), .B(n27), .C(SHIFT_STROBE), .D(n29), .Y(n40) );
  OAI22X1 U10 ( .A(n13), .B(n25), .C(SHIFT_STROBE), .D(n27), .Y(n39) );
  OAI22X1 U12 ( .A(n13), .B(n23), .C(SHIFT_STROBE), .D(n25), .Y(n38) );
  OAI22X1 U14 ( .A(n13), .B(n21), .C(SHIFT_STROBE), .D(n23), .Y(n37) );
  OAI22X1 U16 ( .A(n13), .B(n19), .C(SHIFT_STROBE), .D(n21), .Y(n36) );
  OAI22X1 U18 ( .A(n13), .B(n17), .C(SHIFT_STROBE), .D(n19), .Y(n35) );
  OAI21X1 U22 ( .A(SHIFT_STROBE), .B(n17), .C(n44), .Y(n34) );
  NAND2X1 U23 ( .A(SERIAL_IN), .B(SHIFT_STROBE), .Y(n44) );
  DFFSR \present_val_reg[9]  ( .D(n34), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        STOP_DATA[1]) );
  DFFSR \present_val_reg[8]  ( .D(n35), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        STOP_DATA[0]) );
  DFFSR \present_val_reg[7]  ( .D(n36), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[7]) );
  DFFSR \present_val_reg[6]  ( .D(n37), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[6]) );
  DFFSR \present_val_reg[5]  ( .D(n38), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[5]) );
  DFFSR \present_val_reg[4]  ( .D(n39), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[4]) );
  DFFSR \present_val_reg[3]  ( .D(n40), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[3]) );
  DFFSR \present_val_reg[2]  ( .D(n41), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[2]) );
  DFFSR \present_val_reg[1]  ( .D(n42), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[1]) );
  DFFSR \present_val_reg[0]  ( .D(n43), .CLK(CLK), .R(n15), .S(1'b1), .Q(
        LOAD_DATA[0]) );
  INVX2 U24 ( .A(RST), .Y(n15) );
  INVX2 U25 ( .A(SHIFT_STROBE), .Y(n13) );
  INVX2 U26 ( .A(STOP_DATA[1]), .Y(n17) );
  INVX2 U27 ( .A(STOP_DATA[0]), .Y(n19) );
  INVX2 U28 ( .A(LOAD_DATA[7]), .Y(n21) );
  INVX2 U29 ( .A(LOAD_DATA[6]), .Y(n23) );
  INVX2 U30 ( .A(LOAD_DATA[5]), .Y(n25) );
  INVX2 U31 ( .A(LOAD_DATA[4]), .Y(n27) );
  INVX2 U32 ( .A(LOAD_DATA[3]), .Y(n29) );
  INVX2 U33 ( .A(LOAD_DATA[2]), .Y(n31) );
  INVX2 U34 ( .A(LOAD_DATA[1]), .Y(n32) );
endmodule


module keyreg_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module keyreg_0 ( CLK, RST, SBE, OE, RBUF_FULL, RCV_DATA, PLAINKEY, KEY_ERROR, 
        PROG_ERROR, CLR_RBUFF, PARITY_ERROR );
  input [7:0] RCV_DATA;
  output [63:0] PLAINKEY;
  input CLK, RST, SBE, OE, RBUF_FULL;
  output KEY_ERROR, PROG_ERROR, CLR_RBUFF, PARITY_ERROR;
  wire   parityError, nextParityError, N694, N1792, N1793, N1794, N1795, N1796,
         N1797, N1798, N1799, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n14,
         n16, n17, n19, n20, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39,
         n41, n43, n45, n47, n49, n51, n53, n55, n57, n71, n73, n75, n77, n79,
         n81, n83, n85, n87, n89, n91, n93, n95, n97, n99, n101, n103, n105,
         n107, n109, n111, n113, n115, n117, n119, n121, n123, n125, n127,
         n129, n131, n133, n135, n137, n139, n141, n143, n145, n147, n149,
         n150, n151, n153, n154, n156, n158, n160, n161, n165, n166, n168,
         n172, n173, n175, n177, n178, n180, n181, n183, n184, n185, n186,
         n187, n188, n189, n192, n193, n195, n197, n203, n205, n206, n207,
         n208, n209, n210, n217, n219, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n240, n241, n242,
         n243, n244, n245, n247, n248, n249, n250, n255, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n275, n277, n278, n279, n280, n281, n282, n284, n285, n286,
         n287, n289, n291, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n311, n312, n313, n314, n315, n316, n317, n319,
         n320, n321, n322, n324, n326, n327, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n343, n344, n345, n346, n347,
         n348, n350, n351, n352, n353, n355, n357, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n373, n374, n375, n376,
         n377, n378, n380, n381, n382, n383, n385, n387, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n404, n405, n406,
         n407, n408, n409, n411, n412, n413, n414, n416, n418, n419, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n435,
         n436, n437, n438, n439, n440, n441, n443, n444, n445, n446, n448,
         n450, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n465, n466, n467, n468, n469, n471, n472, n473, n474, n476,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n492, n493, n494, n495, n496, n498, n499, n500, n501, n503, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n519,
         n520, n521, n522, n523, n525, n526, n527, n528, n530, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n547, n548,
         n549, n550, n551, n552, n554, n555, n556, n557, n559, n561, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n576,
         n577, n578, n579, n580, n582, n583, n584, n585, n587, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n603, n604,
         n605, n606, n607, n609, n610, n611, n612, n614, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n630, n631, n632,
         n633, n634, n636, n637, n638, n639, n641, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n657, n658, n659, n660,
         n661, n662, n663, n665, n666, n667, n668, n670, n672, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n687, n688,
         n689, n690, n691, n693, n694, n695, n696, n698, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n714, n715, n716,
         n717, n718, n720, n721, n722, n723, n725, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n741, n742, n743, n744,
         n745, n747, n748, n749, n750, n752, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n769, n770, n771, n772, n773,
         n774, n776, n777, n778, n779, n781, n783, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n798, n799, n800, n801,
         n802, n804, n805, n806, n807, n809, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n825, n826, n827, n828, n829,
         n831, n832, n833, n834, n836, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n852, n853, n854, n855, n856, n858,
         n859, n860, n861, n863, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n879, n880, n881, n882, n883, n884, n885,
         n887, n888, n889, n890, n892, n894, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n909, n910, n911, n912, n913,
         n915, n916, n917, n918, n920, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n936, n937, n938, n939, n940, n942,
         n943, n944, n945, n947, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n963, n964, n965, n966, n967, n969, n970,
         n971, n972, n974, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1003, n1005, n1007, n1008, n1009, n1010, n1012,
         n1013, n1014, n1015, n1016, n1017, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1032, n1035, n1036, n1037,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1102, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037;
  wire   [3:0] state;
  wire   [3:0] keyCount;
  wire   [7:0] address;
  wire   [63:0] currentPlainKey;
  wire   [7:0] parityAccumulator;

  DFFPOSX1 \keyCount_reg[0]  ( .D(n1577), .CLK(CLK), .Q(keyCount[0]) );
  DFFPOSX1 \keyCount_reg[2]  ( .D(n1584), .CLK(CLK), .Q(keyCount[2]) );
  DFFPOSX1 \keyCount_reg[3]  ( .D(n1578), .CLK(CLK), .Q(keyCount[3]) );
  DFFPOSX1 \parityAccumulator_reg[0]  ( .D(n1585), .CLK(CLK), .Q(
        parityAccumulator[0]) );
  DFFPOSX1 \parityAccumulator_reg[1]  ( .D(n1586), .CLK(CLK), .Q(
        parityAccumulator[1]) );
  DFFPOSX1 \parityAccumulator_reg[2]  ( .D(n1587), .CLK(CLK), .Q(
        parityAccumulator[2]) );
  DFFPOSX1 \parityAccumulator_reg[3]  ( .D(n1588), .CLK(CLK), .Q(
        parityAccumulator[3]) );
  DFFPOSX1 \parityAccumulator_reg[4]  ( .D(n1589), .CLK(CLK), .Q(
        parityAccumulator[4]) );
  DFFPOSX1 \parityAccumulator_reg[5]  ( .D(n1590), .CLK(CLK), .Q(
        parityAccumulator[5]) );
  DFFPOSX1 \parityAccumulator_reg[6]  ( .D(n1591), .CLK(CLK), .Q(
        parityAccumulator[6]) );
  DFFPOSX1 \parityAccumulator_reg[7]  ( .D(n1592), .CLK(CLK), .Q(
        parityAccumulator[7]) );
  DFFPOSX1 \keyCount_reg[1]  ( .D(n1583), .CLK(CLK), .Q(keyCount[1]) );
  DFFPOSX1 \address_reg[7]  ( .D(n1593), .CLK(CLK), .Q(address[7]) );
  DFFPOSX1 \address_reg[6]  ( .D(n1594), .CLK(CLK), .Q(address[6]) );
  DFFPOSX1 \address_reg[5]  ( .D(n1595), .CLK(CLK), .Q(address[5]) );
  DFFPOSX1 \address_reg[4]  ( .D(n1596), .CLK(CLK), .Q(address[4]) );
  DFFPOSX1 \address_reg[3]  ( .D(n1597), .CLK(CLK), .Q(address[3]) );
  DFFPOSX1 \address_reg[2]  ( .D(n1598), .CLK(CLK), .Q(address[2]) );
  DFFPOSX1 \address_reg[1]  ( .D(n1599), .CLK(CLK), .Q(address[1]) );
  DFFPOSX1 \address_reg[0]  ( .D(n1600), .CLK(CLK), .Q(address[0]) );
  DFFPOSX1 \currentPlainKey_reg[63]  ( .D(n1664), .CLK(CLK), .Q(
        currentPlainKey[63]) );
  DFFPOSX1 \currentPlainKey_reg[62]  ( .D(n1663), .CLK(CLK), .Q(
        currentPlainKey[62]) );
  DFFPOSX1 \currentPlainKey_reg[61]  ( .D(n1662), .CLK(CLK), .Q(
        currentPlainKey[61]) );
  DFFPOSX1 \currentPlainKey_reg[60]  ( .D(n1661), .CLK(CLK), .Q(
        currentPlainKey[60]) );
  DFFPOSX1 \currentPlainKey_reg[59]  ( .D(n1660), .CLK(CLK), .Q(
        currentPlainKey[59]) );
  DFFPOSX1 \currentPlainKey_reg[58]  ( .D(n1659), .CLK(CLK), .Q(
        currentPlainKey[58]) );
  DFFPOSX1 \currentPlainKey_reg[57]  ( .D(n1658), .CLK(CLK), .Q(
        currentPlainKey[57]) );
  DFFPOSX1 \currentPlainKey_reg[56]  ( .D(n1657), .CLK(CLK), .Q(
        currentPlainKey[56]) );
  DFFPOSX1 \currentPlainKey_reg[55]  ( .D(n1656), .CLK(CLK), .Q(
        currentPlainKey[55]) );
  DFFPOSX1 \currentPlainKey_reg[54]  ( .D(n1655), .CLK(CLK), .Q(
        currentPlainKey[54]) );
  DFFPOSX1 \currentPlainKey_reg[53]  ( .D(n1654), .CLK(CLK), .Q(
        currentPlainKey[53]) );
  DFFPOSX1 \currentPlainKey_reg[52]  ( .D(n1653), .CLK(CLK), .Q(
        currentPlainKey[52]) );
  DFFPOSX1 \currentPlainKey_reg[51]  ( .D(n1652), .CLK(CLK), .Q(
        currentPlainKey[51]) );
  DFFPOSX1 \currentPlainKey_reg[50]  ( .D(n1651), .CLK(CLK), .Q(
        currentPlainKey[50]) );
  DFFPOSX1 \currentPlainKey_reg[49]  ( .D(n1650), .CLK(CLK), .Q(
        currentPlainKey[49]) );
  DFFPOSX1 \currentPlainKey_reg[48]  ( .D(n1649), .CLK(CLK), .Q(
        currentPlainKey[48]) );
  DFFPOSX1 \currentPlainKey_reg[47]  ( .D(n1648), .CLK(CLK), .Q(
        currentPlainKey[47]) );
  DFFPOSX1 \currentPlainKey_reg[46]  ( .D(n1647), .CLK(CLK), .Q(
        currentPlainKey[46]) );
  DFFPOSX1 \currentPlainKey_reg[45]  ( .D(n1646), .CLK(CLK), .Q(
        currentPlainKey[45]) );
  DFFPOSX1 \currentPlainKey_reg[44]  ( .D(n1645), .CLK(CLK), .Q(
        currentPlainKey[44]) );
  DFFPOSX1 \currentPlainKey_reg[43]  ( .D(n1644), .CLK(CLK), .Q(
        currentPlainKey[43]) );
  DFFPOSX1 \currentPlainKey_reg[42]  ( .D(n1643), .CLK(CLK), .Q(
        currentPlainKey[42]) );
  DFFPOSX1 \currentPlainKey_reg[41]  ( .D(n1642), .CLK(CLK), .Q(
        currentPlainKey[41]) );
  DFFPOSX1 \currentPlainKey_reg[40]  ( .D(n1641), .CLK(CLK), .Q(
        currentPlainKey[40]) );
  DFFPOSX1 \currentPlainKey_reg[39]  ( .D(n1640), .CLK(CLK), .Q(
        currentPlainKey[39]) );
  DFFPOSX1 \currentPlainKey_reg[38]  ( .D(n1639), .CLK(CLK), .Q(
        currentPlainKey[38]) );
  DFFPOSX1 \currentPlainKey_reg[37]  ( .D(n1638), .CLK(CLK), .Q(
        currentPlainKey[37]) );
  DFFPOSX1 \currentPlainKey_reg[36]  ( .D(n1637), .CLK(CLK), .Q(
        currentPlainKey[36]) );
  DFFPOSX1 \currentPlainKey_reg[35]  ( .D(n1636), .CLK(CLK), .Q(
        currentPlainKey[35]) );
  DFFPOSX1 \currentPlainKey_reg[34]  ( .D(n1635), .CLK(CLK), .Q(
        currentPlainKey[34]) );
  DFFPOSX1 \currentPlainKey_reg[33]  ( .D(n1634), .CLK(CLK), .Q(
        currentPlainKey[33]) );
  DFFPOSX1 \currentPlainKey_reg[32]  ( .D(n1633), .CLK(CLK), .Q(
        currentPlainKey[32]) );
  DFFPOSX1 \currentPlainKey_reg[31]  ( .D(n1632), .CLK(CLK), .Q(
        currentPlainKey[31]) );
  DFFPOSX1 \currentPlainKey_reg[30]  ( .D(n1631), .CLK(CLK), .Q(
        currentPlainKey[30]) );
  DFFPOSX1 \currentPlainKey_reg[29]  ( .D(n1630), .CLK(CLK), .Q(
        currentPlainKey[29]) );
  DFFPOSX1 \currentPlainKey_reg[28]  ( .D(n1629), .CLK(CLK), .Q(
        currentPlainKey[28]) );
  DFFPOSX1 \currentPlainKey_reg[27]  ( .D(n1628), .CLK(CLK), .Q(
        currentPlainKey[27]) );
  DFFPOSX1 \currentPlainKey_reg[26]  ( .D(n1627), .CLK(CLK), .Q(
        currentPlainKey[26]) );
  DFFPOSX1 \currentPlainKey_reg[25]  ( .D(n1626), .CLK(CLK), .Q(
        currentPlainKey[25]) );
  DFFPOSX1 \currentPlainKey_reg[24]  ( .D(n1625), .CLK(CLK), .Q(
        currentPlainKey[24]) );
  DFFPOSX1 \currentPlainKey_reg[23]  ( .D(n1624), .CLK(CLK), .Q(
        currentPlainKey[23]) );
  DFFPOSX1 \currentPlainKey_reg[22]  ( .D(n1623), .CLK(CLK), .Q(
        currentPlainKey[22]) );
  DFFPOSX1 \currentPlainKey_reg[21]  ( .D(n1622), .CLK(CLK), .Q(
        currentPlainKey[21]) );
  DFFPOSX1 \currentPlainKey_reg[20]  ( .D(n1621), .CLK(CLK), .Q(
        currentPlainKey[20]) );
  DFFPOSX1 \currentPlainKey_reg[19]  ( .D(n1620), .CLK(CLK), .Q(
        currentPlainKey[19]) );
  DFFPOSX1 \currentPlainKey_reg[18]  ( .D(n1619), .CLK(CLK), .Q(
        currentPlainKey[18]) );
  DFFPOSX1 \currentPlainKey_reg[17]  ( .D(n1618), .CLK(CLK), .Q(
        currentPlainKey[17]) );
  DFFPOSX1 \currentPlainKey_reg[16]  ( .D(n1617), .CLK(CLK), .Q(
        currentPlainKey[16]) );
  DFFPOSX1 \currentPlainKey_reg[15]  ( .D(n1616), .CLK(CLK), .Q(
        currentPlainKey[15]) );
  DFFPOSX1 \currentPlainKey_reg[14]  ( .D(n1615), .CLK(CLK), .Q(
        currentPlainKey[14]) );
  DFFPOSX1 \currentPlainKey_reg[13]  ( .D(n1614), .CLK(CLK), .Q(
        currentPlainKey[13]) );
  DFFPOSX1 \currentPlainKey_reg[12]  ( .D(n1613), .CLK(CLK), .Q(
        currentPlainKey[12]) );
  DFFPOSX1 \currentPlainKey_reg[11]  ( .D(n1612), .CLK(CLK), .Q(
        currentPlainKey[11]) );
  DFFPOSX1 \currentPlainKey_reg[10]  ( .D(n1611), .CLK(CLK), .Q(
        currentPlainKey[10]) );
  DFFPOSX1 \currentPlainKey_reg[9]  ( .D(n1610), .CLK(CLK), .Q(
        currentPlainKey[9]) );
  DFFPOSX1 \currentPlainKey_reg[8]  ( .D(n1609), .CLK(CLK), .Q(
        currentPlainKey[8]) );
  DFFPOSX1 \currentPlainKey_reg[7]  ( .D(n1608), .CLK(CLK), .Q(
        currentPlainKey[7]) );
  DFFPOSX1 \currentPlainKey_reg[6]  ( .D(n1607), .CLK(CLK), .Q(
        currentPlainKey[6]) );
  DFFPOSX1 \currentPlainKey_reg[5]  ( .D(n1606), .CLK(CLK), .Q(
        currentPlainKey[5]) );
  DFFPOSX1 \currentPlainKey_reg[4]  ( .D(n1605), .CLK(CLK), .Q(
        currentPlainKey[4]) );
  DFFPOSX1 \currentPlainKey_reg[3]  ( .D(n1604), .CLK(CLK), .Q(
        currentPlainKey[3]) );
  DFFPOSX1 \currentPlainKey_reg[2]  ( .D(n1603), .CLK(CLK), .Q(
        currentPlainKey[2]) );
  DFFPOSX1 \currentPlainKey_reg[1]  ( .D(n1602), .CLK(CLK), .Q(
        currentPlainKey[1]) );
  DFFPOSX1 \currentPlainKey_reg[0]  ( .D(n1601), .CLK(CLK), .Q(
        currentPlainKey[0]) );
  DFFPOSX1 \PLAINKEY_reg[63]  ( .D(n1665), .CLK(CLK), .Q(PLAINKEY[63]) );
  DFFPOSX1 \PLAINKEY_reg[62]  ( .D(n1666), .CLK(CLK), .Q(PLAINKEY[62]) );
  DFFPOSX1 \PLAINKEY_reg[61]  ( .D(n1667), .CLK(CLK), .Q(PLAINKEY[61]) );
  DFFPOSX1 \PLAINKEY_reg[60]  ( .D(n1668), .CLK(CLK), .Q(PLAINKEY[60]) );
  DFFPOSX1 \PLAINKEY_reg[59]  ( .D(n1669), .CLK(CLK), .Q(PLAINKEY[59]) );
  DFFPOSX1 \PLAINKEY_reg[58]  ( .D(n1670), .CLK(CLK), .Q(PLAINKEY[58]) );
  DFFPOSX1 \PLAINKEY_reg[57]  ( .D(n1671), .CLK(CLK), .Q(PLAINKEY[57]) );
  DFFPOSX1 \PLAINKEY_reg[56]  ( .D(n1672), .CLK(CLK), .Q(PLAINKEY[56]) );
  DFFPOSX1 \PLAINKEY_reg[55]  ( .D(n1673), .CLK(CLK), .Q(PLAINKEY[55]) );
  DFFPOSX1 \PLAINKEY_reg[54]  ( .D(n1674), .CLK(CLK), .Q(PLAINKEY[54]) );
  DFFPOSX1 \PLAINKEY_reg[53]  ( .D(n1675), .CLK(CLK), .Q(PLAINKEY[53]) );
  DFFPOSX1 \PLAINKEY_reg[52]  ( .D(n1676), .CLK(CLK), .Q(PLAINKEY[52]) );
  DFFPOSX1 \PLAINKEY_reg[51]  ( .D(n1677), .CLK(CLK), .Q(PLAINKEY[51]) );
  DFFPOSX1 \PLAINKEY_reg[50]  ( .D(n1678), .CLK(CLK), .Q(PLAINKEY[50]) );
  DFFPOSX1 \PLAINKEY_reg[49]  ( .D(n1679), .CLK(CLK), .Q(PLAINKEY[49]) );
  DFFPOSX1 \PLAINKEY_reg[48]  ( .D(n1680), .CLK(CLK), .Q(PLAINKEY[48]) );
  DFFPOSX1 \PLAINKEY_reg[47]  ( .D(n1681), .CLK(CLK), .Q(PLAINKEY[47]) );
  DFFPOSX1 \PLAINKEY_reg[46]  ( .D(n1682), .CLK(CLK), .Q(PLAINKEY[46]) );
  DFFPOSX1 \PLAINKEY_reg[45]  ( .D(n1683), .CLK(CLK), .Q(PLAINKEY[45]) );
  DFFPOSX1 \PLAINKEY_reg[44]  ( .D(n1684), .CLK(CLK), .Q(PLAINKEY[44]) );
  DFFPOSX1 \PLAINKEY_reg[43]  ( .D(n1685), .CLK(CLK), .Q(PLAINKEY[43]) );
  DFFPOSX1 \PLAINKEY_reg[42]  ( .D(n1686), .CLK(CLK), .Q(PLAINKEY[42]) );
  DFFPOSX1 \PLAINKEY_reg[41]  ( .D(n1687), .CLK(CLK), .Q(PLAINKEY[41]) );
  DFFPOSX1 \PLAINKEY_reg[40]  ( .D(n1688), .CLK(CLK), .Q(PLAINKEY[40]) );
  DFFPOSX1 \PLAINKEY_reg[39]  ( .D(n1689), .CLK(CLK), .Q(PLAINKEY[39]) );
  DFFPOSX1 \PLAINKEY_reg[38]  ( .D(n1690), .CLK(CLK), .Q(PLAINKEY[38]) );
  DFFPOSX1 \PLAINKEY_reg[37]  ( .D(n1691), .CLK(CLK), .Q(PLAINKEY[37]) );
  DFFPOSX1 \PLAINKEY_reg[36]  ( .D(n1692), .CLK(CLK), .Q(PLAINKEY[36]) );
  DFFPOSX1 \PLAINKEY_reg[35]  ( .D(n1693), .CLK(CLK), .Q(PLAINKEY[35]) );
  DFFPOSX1 \PLAINKEY_reg[34]  ( .D(n1694), .CLK(CLK), .Q(PLAINKEY[34]) );
  DFFPOSX1 \PLAINKEY_reg[33]  ( .D(n1695), .CLK(CLK), .Q(PLAINKEY[33]) );
  DFFPOSX1 \PLAINKEY_reg[32]  ( .D(n1696), .CLK(CLK), .Q(PLAINKEY[32]) );
  DFFPOSX1 \PLAINKEY_reg[31]  ( .D(n1697), .CLK(CLK), .Q(PLAINKEY[31]) );
  DFFPOSX1 \PLAINKEY_reg[30]  ( .D(n1698), .CLK(CLK), .Q(PLAINKEY[30]) );
  DFFPOSX1 \PLAINKEY_reg[29]  ( .D(n1699), .CLK(CLK), .Q(PLAINKEY[29]) );
  DFFPOSX1 \PLAINKEY_reg[28]  ( .D(n1700), .CLK(CLK), .Q(PLAINKEY[28]) );
  DFFPOSX1 \PLAINKEY_reg[27]  ( .D(n1701), .CLK(CLK), .Q(PLAINKEY[27]) );
  DFFPOSX1 \PLAINKEY_reg[26]  ( .D(n1702), .CLK(CLK), .Q(PLAINKEY[26]) );
  DFFPOSX1 \PLAINKEY_reg[25]  ( .D(n1703), .CLK(CLK), .Q(PLAINKEY[25]) );
  DFFPOSX1 \PLAINKEY_reg[24]  ( .D(n1704), .CLK(CLK), .Q(PLAINKEY[24]) );
  DFFPOSX1 \PLAINKEY_reg[23]  ( .D(n1705), .CLK(CLK), .Q(PLAINKEY[23]) );
  DFFPOSX1 \PLAINKEY_reg[22]  ( .D(n1706), .CLK(CLK), .Q(PLAINKEY[22]) );
  DFFPOSX1 \PLAINKEY_reg[21]  ( .D(n1707), .CLK(CLK), .Q(PLAINKEY[21]) );
  DFFPOSX1 \PLAINKEY_reg[20]  ( .D(n1708), .CLK(CLK), .Q(PLAINKEY[20]) );
  DFFPOSX1 \PLAINKEY_reg[19]  ( .D(n1709), .CLK(CLK), .Q(PLAINKEY[19]) );
  DFFPOSX1 \PLAINKEY_reg[18]  ( .D(n1710), .CLK(CLK), .Q(PLAINKEY[18]) );
  DFFPOSX1 \PLAINKEY_reg[17]  ( .D(n1711), .CLK(CLK), .Q(PLAINKEY[17]) );
  DFFPOSX1 \PLAINKEY_reg[16]  ( .D(n1712), .CLK(CLK), .Q(PLAINKEY[16]) );
  DFFPOSX1 \PLAINKEY_reg[15]  ( .D(n1713), .CLK(CLK), .Q(PLAINKEY[15]) );
  DFFPOSX1 \PLAINKEY_reg[14]  ( .D(n1714), .CLK(CLK), .Q(PLAINKEY[14]) );
  DFFPOSX1 \PLAINKEY_reg[13]  ( .D(n1715), .CLK(CLK), .Q(PLAINKEY[13]) );
  DFFPOSX1 \PLAINKEY_reg[12]  ( .D(n1716), .CLK(CLK), .Q(PLAINKEY[12]) );
  DFFPOSX1 \PLAINKEY_reg[11]  ( .D(n1717), .CLK(CLK), .Q(PLAINKEY[11]) );
  DFFPOSX1 \PLAINKEY_reg[10]  ( .D(n1718), .CLK(CLK), .Q(PLAINKEY[10]) );
  DFFPOSX1 \PLAINKEY_reg[9]  ( .D(n1719), .CLK(CLK), .Q(PLAINKEY[9]) );
  DFFPOSX1 \PLAINKEY_reg[8]  ( .D(n1720), .CLK(CLK), .Q(PLAINKEY[8]) );
  DFFPOSX1 \PLAINKEY_reg[7]  ( .D(n1721), .CLK(CLK), .Q(PLAINKEY[7]) );
  DFFPOSX1 \PLAINKEY_reg[6]  ( .D(n1722), .CLK(CLK), .Q(PLAINKEY[6]) );
  DFFPOSX1 \PLAINKEY_reg[5]  ( .D(n1723), .CLK(CLK), .Q(PLAINKEY[5]) );
  DFFPOSX1 \PLAINKEY_reg[4]  ( .D(n1724), .CLK(CLK), .Q(PLAINKEY[4]) );
  DFFPOSX1 \PLAINKEY_reg[3]  ( .D(n1725), .CLK(CLK), .Q(PLAINKEY[3]) );
  DFFPOSX1 \PLAINKEY_reg[2]  ( .D(n1726), .CLK(CLK), .Q(PLAINKEY[2]) );
  DFFPOSX1 \PLAINKEY_reg[1]  ( .D(n1727), .CLK(CLK), .Q(PLAINKEY[1]) );
  DFFPOSX1 \PLAINKEY_reg[0]  ( .D(n1728), .CLK(CLK), .Q(PLAINKEY[0]) );
  NAND3X1 U9 ( .A(parityAccumulator[7]), .B(parityAccumulator[6]), .C(n2035), 
        .Y(n2036) );
  NOR2X1 U10 ( .A(n1486), .B(n1487), .Y(n2035) );
  NAND3X1 U11 ( .A(parityAccumulator[3]), .B(parityAccumulator[2]), .C(n2034), 
        .Y(n2037) );
  NOR2X1 U12 ( .A(n1482), .B(n1483), .Y(n2034) );
  OAI21X1 U13 ( .A(n223), .B(n1569), .C(n2033), .Y(n1728) );
  NAND2X1 U14 ( .A(PLAINKEY[0]), .B(n227), .Y(n2033) );
  OAI21X1 U15 ( .A(n223), .B(n1568), .C(n2032), .Y(n1727) );
  NAND2X1 U16 ( .A(PLAINKEY[1]), .B(RST), .Y(n2032) );
  OAI21X1 U17 ( .A(n223), .B(n1567), .C(n2031), .Y(n1726) );
  NAND2X1 U18 ( .A(PLAINKEY[2]), .B(RST), .Y(n2031) );
  OAI21X1 U19 ( .A(n223), .B(n1566), .C(n2030), .Y(n1725) );
  NAND2X1 U20 ( .A(PLAINKEY[3]), .B(RST), .Y(n2030) );
  OAI21X1 U21 ( .A(n223), .B(n1565), .C(n2029), .Y(n1724) );
  NAND2X1 U22 ( .A(PLAINKEY[4]), .B(n227), .Y(n2029) );
  OAI21X1 U24 ( .A(n223), .B(n1564), .C(n2028), .Y(n1723) );
  NAND2X1 U25 ( .A(PLAINKEY[5]), .B(n228), .Y(n2028) );
  OAI21X1 U27 ( .A(n223), .B(n1563), .C(n2027), .Y(n1722) );
  NAND2X1 U28 ( .A(PLAINKEY[6]), .B(n229), .Y(n2027) );
  OAI21X1 U30 ( .A(n223), .B(n1562), .C(n2026), .Y(n1721) );
  NAND2X1 U31 ( .A(PLAINKEY[7]), .B(RST), .Y(n2026) );
  OAI21X1 U33 ( .A(n223), .B(n1561), .C(n2025), .Y(n1720) );
  NAND2X1 U34 ( .A(PLAINKEY[8]), .B(n227), .Y(n2025) );
  OAI21X1 U36 ( .A(n224), .B(n1560), .C(n2024), .Y(n1719) );
  NAND2X1 U37 ( .A(PLAINKEY[9]), .B(n228), .Y(n2024) );
  OAI21X1 U39 ( .A(n224), .B(n1559), .C(n2023), .Y(n1718) );
  NAND2X1 U40 ( .A(PLAINKEY[10]), .B(n229), .Y(n2023) );
  OAI21X1 U42 ( .A(n224), .B(n1558), .C(n2022), .Y(n1717) );
  NAND2X1 U43 ( .A(PLAINKEY[11]), .B(n229), .Y(n2022) );
  OAI21X1 U45 ( .A(n224), .B(n1557), .C(n2021), .Y(n1716) );
  NAND2X1 U46 ( .A(PLAINKEY[12]), .B(n229), .Y(n2021) );
  OAI21X1 U48 ( .A(n224), .B(n1556), .C(n2020), .Y(n1715) );
  NAND2X1 U49 ( .A(PLAINKEY[13]), .B(n229), .Y(n2020) );
  OAI21X1 U51 ( .A(n224), .B(n1555), .C(n2019), .Y(n1714) );
  NAND2X1 U52 ( .A(PLAINKEY[14]), .B(n229), .Y(n2019) );
  OAI21X1 U54 ( .A(n224), .B(n1554), .C(n2018), .Y(n1713) );
  NAND2X1 U55 ( .A(PLAINKEY[15]), .B(n229), .Y(n2018) );
  OAI21X1 U57 ( .A(n225), .B(n1553), .C(n2017), .Y(n1712) );
  NAND2X1 U58 ( .A(PLAINKEY[16]), .B(n229), .Y(n2017) );
  OAI21X1 U60 ( .A(n225), .B(n1552), .C(n2016), .Y(n1711) );
  NAND2X1 U61 ( .A(PLAINKEY[17]), .B(n229), .Y(n2016) );
  OAI21X1 U63 ( .A(n225), .B(n1551), .C(n2015), .Y(n1710) );
  NAND2X1 U64 ( .A(PLAINKEY[18]), .B(n229), .Y(n2015) );
  OAI21X1 U66 ( .A(n225), .B(n1550), .C(n2014), .Y(n1709) );
  NAND2X1 U67 ( .A(PLAINKEY[19]), .B(n229), .Y(n2014) );
  OAI21X1 U69 ( .A(n225), .B(n1549), .C(n2013), .Y(n1708) );
  NAND2X1 U70 ( .A(PLAINKEY[20]), .B(n229), .Y(n2013) );
  OAI21X1 U72 ( .A(n225), .B(n1548), .C(n2012), .Y(n1707) );
  NAND2X1 U73 ( .A(PLAINKEY[21]), .B(n229), .Y(n2012) );
  OAI21X1 U75 ( .A(n225), .B(n1547), .C(n2011), .Y(n1706) );
  NAND2X1 U76 ( .A(PLAINKEY[22]), .B(n229), .Y(n2011) );
  OAI21X1 U78 ( .A(n226), .B(n1546), .C(n2010), .Y(n1705) );
  NAND2X1 U79 ( .A(PLAINKEY[23]), .B(n229), .Y(n2010) );
  OAI21X1 U81 ( .A(n225), .B(n1545), .C(n2009), .Y(n1704) );
  NAND2X1 U82 ( .A(PLAINKEY[24]), .B(n229), .Y(n2009) );
  OAI21X1 U84 ( .A(n224), .B(n1544), .C(n2008), .Y(n1703) );
  NAND2X1 U85 ( .A(PLAINKEY[25]), .B(n229), .Y(n2008) );
  OAI21X1 U87 ( .A(n226), .B(n1543), .C(n2007), .Y(n1702) );
  NAND2X1 U88 ( .A(PLAINKEY[26]), .B(n229), .Y(n2007) );
  OAI21X1 U90 ( .A(n226), .B(n1542), .C(n2006), .Y(n1701) );
  NAND2X1 U91 ( .A(PLAINKEY[27]), .B(n229), .Y(n2006) );
  OAI21X1 U93 ( .A(n225), .B(n1541), .C(n2005), .Y(n1700) );
  NAND2X1 U94 ( .A(PLAINKEY[28]), .B(n229), .Y(n2005) );
  OAI21X1 U96 ( .A(n226), .B(n1540), .C(n2004), .Y(n1699) );
  NAND2X1 U97 ( .A(PLAINKEY[29]), .B(n228), .Y(n2004) );
  OAI21X1 U99 ( .A(n226), .B(n1539), .C(n2003), .Y(n1698) );
  NAND2X1 U100 ( .A(PLAINKEY[30]), .B(n228), .Y(n2003) );
  OAI21X1 U102 ( .A(n225), .B(n1538), .C(n2002), .Y(n1697) );
  NAND2X1 U103 ( .A(PLAINKEY[31]), .B(n228), .Y(n2002) );
  OAI21X1 U105 ( .A(RST), .B(n1537), .C(n2001), .Y(n1696) );
  NAND2X1 U106 ( .A(PLAINKEY[32]), .B(n228), .Y(n2001) );
  OAI21X1 U108 ( .A(n226), .B(n1536), .C(n2000), .Y(n1695) );
  NAND2X1 U109 ( .A(PLAINKEY[33]), .B(n228), .Y(n2000) );
  OAI21X1 U111 ( .A(n229), .B(n1535), .C(n1999), .Y(n1694) );
  NAND2X1 U112 ( .A(PLAINKEY[34]), .B(n228), .Y(n1999) );
  OAI21X1 U114 ( .A(n226), .B(n1534), .C(n1998), .Y(n1693) );
  NAND2X1 U115 ( .A(PLAINKEY[35]), .B(n228), .Y(n1998) );
  OAI21X1 U117 ( .A(n226), .B(n1533), .C(n1997), .Y(n1692) );
  NAND2X1 U118 ( .A(PLAINKEY[36]), .B(n228), .Y(n1997) );
  OAI21X1 U120 ( .A(n227), .B(n1532), .C(n1996), .Y(n1691) );
  NAND2X1 U121 ( .A(PLAINKEY[37]), .B(n228), .Y(n1996) );
  OAI21X1 U123 ( .A(n223), .B(n1531), .C(n1995), .Y(n1690) );
  NAND2X1 U124 ( .A(PLAINKEY[38]), .B(n228), .Y(n1995) );
  OAI21X1 U126 ( .A(n226), .B(n1530), .C(n1994), .Y(n1689) );
  NAND2X1 U127 ( .A(PLAINKEY[39]), .B(n228), .Y(n1994) );
  OAI21X1 U129 ( .A(n225), .B(n1529), .C(n1993), .Y(n1688) );
  NAND2X1 U130 ( .A(PLAINKEY[40]), .B(n228), .Y(n1993) );
  OAI21X1 U132 ( .A(n226), .B(n1528), .C(n1992), .Y(n1687) );
  NAND2X1 U133 ( .A(PLAINKEY[41]), .B(n228), .Y(n1992) );
  OAI21X1 U135 ( .A(n226), .B(n1527), .C(n1991), .Y(n1686) );
  NAND2X1 U136 ( .A(PLAINKEY[42]), .B(n228), .Y(n1991) );
  OAI21X1 U138 ( .A(RST), .B(n1526), .C(n1990), .Y(n1685) );
  NAND2X1 U139 ( .A(PLAINKEY[43]), .B(n228), .Y(n1990) );
  OAI21X1 U141 ( .A(n224), .B(n1525), .C(n1989), .Y(n1684) );
  NAND2X1 U142 ( .A(PLAINKEY[44]), .B(n227), .Y(n1989) );
  OAI21X1 U144 ( .A(n224), .B(n1524), .C(n1988), .Y(n1683) );
  NAND2X1 U145 ( .A(PLAINKEY[45]), .B(n227), .Y(n1988) );
  OAI21X1 U147 ( .A(n228), .B(n1523), .C(n1987), .Y(n1682) );
  NAND2X1 U148 ( .A(PLAINKEY[46]), .B(n228), .Y(n1987) );
  OAI21X1 U150 ( .A(n224), .B(n1522), .C(n1986), .Y(n1681) );
  NAND2X1 U151 ( .A(PLAINKEY[47]), .B(n227), .Y(n1986) );
  OAI21X1 U153 ( .A(n226), .B(n1521), .C(n1985), .Y(n1680) );
  NAND2X1 U154 ( .A(PLAINKEY[48]), .B(n227), .Y(n1985) );
  OAI21X1 U156 ( .A(n226), .B(n1520), .C(n1984), .Y(n1679) );
  NAND2X1 U157 ( .A(PLAINKEY[49]), .B(n227), .Y(n1984) );
  OAI21X1 U159 ( .A(n226), .B(n1519), .C(n1983), .Y(n1678) );
  NAND2X1 U160 ( .A(PLAINKEY[50]), .B(n227), .Y(n1983) );
  OAI21X1 U162 ( .A(n225), .B(n1518), .C(n1982), .Y(n1677) );
  NAND2X1 U163 ( .A(PLAINKEY[51]), .B(n227), .Y(n1982) );
  OAI21X1 U165 ( .A(n226), .B(n1517), .C(n1981), .Y(n1676) );
  NAND2X1 U166 ( .A(PLAINKEY[52]), .B(n227), .Y(n1981) );
  OAI21X1 U168 ( .A(n225), .B(n1516), .C(n1980), .Y(n1675) );
  NAND2X1 U169 ( .A(PLAINKEY[53]), .B(n227), .Y(n1980) );
  OAI21X1 U171 ( .A(n225), .B(n1515), .C(n1979), .Y(n1674) );
  NAND2X1 U172 ( .A(PLAINKEY[54]), .B(n227), .Y(n1979) );
  OAI21X1 U174 ( .A(n224), .B(n1514), .C(n1978), .Y(n1673) );
  NAND2X1 U175 ( .A(PLAINKEY[55]), .B(n228), .Y(n1978) );
  OAI21X1 U177 ( .A(n225), .B(n1513), .C(n1977), .Y(n1672) );
  NAND2X1 U178 ( .A(PLAINKEY[56]), .B(n227), .Y(n1977) );
  OAI21X1 U180 ( .A(n224), .B(n1512), .C(n1976), .Y(n1671) );
  NAND2X1 U181 ( .A(PLAINKEY[57]), .B(n227), .Y(n1976) );
  OAI21X1 U183 ( .A(n224), .B(n1511), .C(n1975), .Y(n1670) );
  NAND2X1 U184 ( .A(PLAINKEY[58]), .B(n227), .Y(n1975) );
  OAI21X1 U186 ( .A(n224), .B(n1510), .C(n1974), .Y(n1669) );
  NAND2X1 U187 ( .A(PLAINKEY[59]), .B(n227), .Y(n1974) );
  OAI21X1 U188 ( .A(n223), .B(n1509), .C(n1973), .Y(n1668) );
  NAND2X1 U189 ( .A(PLAINKEY[60]), .B(n227), .Y(n1973) );
  OAI21X1 U191 ( .A(n223), .B(n1508), .C(n1972), .Y(n1667) );
  NAND2X1 U192 ( .A(PLAINKEY[61]), .B(n227), .Y(n1972) );
  OAI21X1 U194 ( .A(n223), .B(n1507), .C(n1971), .Y(n1666) );
  NAND2X1 U195 ( .A(PLAINKEY[62]), .B(n227), .Y(n1971) );
  OAI21X1 U196 ( .A(n223), .B(n1506), .C(n1970), .Y(n1665) );
  NAND2X1 U197 ( .A(PLAINKEY[63]), .B(n228), .Y(n1970) );
  OAI21X1 U202 ( .A(n1445), .B(n1965), .C(n1967), .Y(n1968) );
  AOI22X1 U203 ( .A(n1964), .B(n1963), .C(n1494), .D(n1572), .Y(n1965) );
  OAI22X1 U205 ( .A(RCV_DATA[3]), .B(n1962), .C(n1495), .D(n1961), .Y(n1964)
         );
  AOI22X1 U206 ( .A(n1960), .B(n1959), .C(n1496), .D(n1574), .Y(n1961) );
  OAI22X1 U208 ( .A(n1958), .B(n1497), .C(n221), .D(n1957), .Y(n1960) );
  NAND2X1 U210 ( .A(n21), .B(n6), .Y(n1957) );
  AOI22X1 U211 ( .A(n1956), .B(n1575), .C(n1503), .D(n1506), .Y(n1958) );
  NOR2X1 U213 ( .A(n1955), .B(n127), .Y(n1956) );
  OAI22X1 U220 ( .A(n1967), .B(n1571), .C(n1966), .D(n1572), .Y(n1953) );
  OAI21X1 U221 ( .A(n1963), .B(n1573), .C(n1952), .Y(n1954) );
  AOI22X1 U222 ( .A(RCV_DATA[2]), .B(n1495), .C(n1492), .D(n1951), .Y(n1952)
         );
  OAI21X1 U223 ( .A(n1959), .B(n222), .C(n1950), .Y(n1951) );
  NAND2X1 U224 ( .A(n1949), .B(n1959), .Y(n1950) );
  OAI21X1 U225 ( .A(n1955), .B(n1948), .C(n1947), .Y(n1949) );
  OAI21X1 U226 ( .A(n1946), .B(n1955), .C(currentPlainKey[62]), .Y(n1947) );
  NAND2X1 U227 ( .A(n20), .B(n6), .Y(n1959) );
  OAI21X1 U233 ( .A(n1943), .B(n1942), .C(n1969), .Y(n1944) );
  OAI22X1 U234 ( .A(n1967), .B(n1572), .C(n1963), .D(n1574), .Y(n1942) );
  OAI21X1 U235 ( .A(n1941), .B(n1945), .C(n1940), .Y(n1943) );
  AOI22X1 U236 ( .A(n221), .B(n1495), .C(RCV_DATA[3]), .D(n1445), .Y(n1940) );
  NAND2X1 U238 ( .A(n1939), .B(n1962), .Y(n1945) );
  NAND2X1 U239 ( .A(n19), .B(n6), .Y(n1962) );
  AOI22X1 U240 ( .A(n1938), .B(n139), .C(currentPlainKey[61]), .D(n1502), .Y(
        n1941) );
  NOR2X1 U242 ( .A(n1955), .B(n1937), .Y(n1938) );
  OAI21X1 U252 ( .A(n1955), .B(n1935), .C(n1934), .Y(n1936) );
  OAI21X1 U253 ( .A(n1933), .B(n1955), .C(currentPlainKey[60]), .Y(n1934) );
  OAI21X1 U264 ( .A(n1967), .B(n1574), .C(n1929), .Y(n1930) );
  AOI22X1 U265 ( .A(n1932), .B(n1928), .C(n221), .D(n1445), .Y(n1929) );
  OAI22X1 U266 ( .A(n1927), .B(n1510), .C(n1575), .D(n1501), .Y(n1928) );
  NOR2X1 U270 ( .A(n1955), .B(n1926), .Y(n1927) );
  NOR2X1 U271 ( .A(n1445), .B(n1493), .Y(n1932) );
  OAI22X1 U284 ( .A(n1967), .B(n222), .C(n1493), .D(n1924), .Y(n1925) );
  AOI22X1 U285 ( .A(n1923), .B(n139), .C(currentPlainKey[58]), .D(n1500), .Y(
        n1924) );
  NOR2X1 U287 ( .A(n1955), .B(n1922), .Y(n1923) );
  AOI22X1 U300 ( .A(n1919), .B(n1969), .C(n221), .D(n1446), .Y(n1920) );
  OAI21X1 U303 ( .A(n1955), .B(n1918), .C(n1917), .Y(n1919) );
  OAI21X1 U304 ( .A(n1916), .B(n1955), .C(currentPlainKey[57]), .Y(n1917) );
  OAI21X1 U314 ( .A(n1955), .B(n1914), .C(n1913), .Y(n1915) );
  OAI21X1 U315 ( .A(n1912), .B(n1955), .C(currentPlainKey[56]), .Y(n1913) );
  NAND2X1 U316 ( .A(address[3]), .B(n1911), .Y(n1955) );
  AOI22X1 U330 ( .A(n1908), .B(n1931), .C(n1447), .D(n221), .Y(n1909) );
  OAI21X1 U333 ( .A(n151), .B(n1907), .C(n1906), .Y(n1908) );
  OAI21X1 U334 ( .A(n127), .B(n151), .C(currentPlainKey[55]), .Y(n1906) );
  OAI21X1 U344 ( .A(n1948), .B(n151), .C(n1904), .Y(n1905) );
  OAI21X1 U345 ( .A(n1946), .B(n151), .C(currentPlainKey[54]), .Y(n1904) );
  AOI22X1 U359 ( .A(n1901), .B(n1921), .C(n1448), .D(n221), .Y(n1902) );
  OAI21X1 U362 ( .A(n151), .B(n1900), .C(n1899), .Y(n1901) );
  OAI21X1 U363 ( .A(n1937), .B(n151), .C(currentPlainKey[53]), .Y(n1899) );
  OAI21X1 U373 ( .A(n1935), .B(n151), .C(n1897), .Y(n1898) );
  OAI21X1 U374 ( .A(n1933), .B(n151), .C(currentPlainKey[52]), .Y(n1897) );
  AOI22X1 U388 ( .A(n1894), .B(n1910), .C(n1449), .D(n221), .Y(n1895) );
  OAI21X1 U391 ( .A(n151), .B(n1893), .C(n1892), .Y(n1894) );
  OAI21X1 U392 ( .A(n1926), .B(n151), .C(currentPlainKey[51]), .Y(n1892) );
  OAI21X1 U402 ( .A(n151), .B(n1890), .C(n1889), .Y(n1891) );
  OAI21X1 U403 ( .A(n1922), .B(n151), .C(currentPlainKey[50]), .Y(n1889) );
  AOI22X1 U417 ( .A(n1886), .B(n1903), .C(n1450), .D(n221), .Y(n1887) );
  OAI21X1 U422 ( .A(n1918), .B(n151), .C(n1884), .Y(n1886) );
  OAI21X1 U423 ( .A(n1916), .B(n151), .C(currentPlainKey[49]), .Y(n1884) );
  OAI21X1 U433 ( .A(n1914), .B(n151), .C(n1882), .Y(n1883) );
  OAI21X1 U434 ( .A(n1912), .B(n151), .C(currentPlainKey[48]), .Y(n1882) );
  AOI22X1 U449 ( .A(n1879), .B(n1896), .C(n1451), .D(n221), .Y(n1880) );
  OAI21X1 U452 ( .A(n1907), .B(n150), .C(n1878), .Y(n1879) );
  OAI21X1 U453 ( .A(n127), .B(n150), .C(currentPlainKey[47]), .Y(n1878) );
  OAI21X1 U463 ( .A(n1948), .B(n150), .C(n1876), .Y(n1877) );
  OAI21X1 U464 ( .A(n1946), .B(n150), .C(currentPlainKey[46]), .Y(n1876) );
  AOI22X1 U478 ( .A(n1873), .B(n1888), .C(n1452), .D(n221), .Y(n1874) );
  OAI21X1 U481 ( .A(n1900), .B(n150), .C(n1872), .Y(n1873) );
  OAI21X1 U482 ( .A(n1937), .B(n150), .C(currentPlainKey[45]), .Y(n1872) );
  OAI21X1 U492 ( .A(n1935), .B(n150), .C(n1870), .Y(n1871) );
  OAI21X1 U493 ( .A(n1933), .B(n150), .C(currentPlainKey[44]), .Y(n1870) );
  AOI22X1 U507 ( .A(n1867), .B(n1881), .C(n1453), .D(n221), .Y(n1868) );
  OAI21X1 U510 ( .A(n1893), .B(n150), .C(n1866), .Y(n1867) );
  OAI21X1 U511 ( .A(n1926), .B(n150), .C(currentPlainKey[43]), .Y(n1866) );
  OAI21X1 U521 ( .A(n1890), .B(n150), .C(n1864), .Y(n1865) );
  OAI21X1 U522 ( .A(n1922), .B(n150), .C(currentPlainKey[42]), .Y(n1864) );
  AOI22X1 U536 ( .A(n1861), .B(n1875), .C(n1454), .D(n221), .Y(n1862) );
  OAI21X1 U539 ( .A(n1918), .B(n150), .C(n1860), .Y(n1861) );
  OAI21X1 U540 ( .A(n1916), .B(n150), .C(currentPlainKey[41]), .Y(n1860) );
  OAI21X1 U550 ( .A(n1914), .B(n150), .C(n1858), .Y(n1859) );
  OAI21X1 U551 ( .A(n1912), .B(n150), .C(currentPlainKey[40]), .Y(n1858) );
  AOI22X1 U566 ( .A(n1854), .B(n1869), .C(n1455), .D(n221), .Y(n1855) );
  OAI21X1 U569 ( .A(n1907), .B(n149), .C(n1853), .Y(n1854) );
  OAI21X1 U570 ( .A(n127), .B(n149), .C(currentPlainKey[39]), .Y(n1853) );
  OAI21X1 U580 ( .A(n1948), .B(n149), .C(n1851), .Y(n1852) );
  OAI21X1 U581 ( .A(n1946), .B(n149), .C(currentPlainKey[38]), .Y(n1851) );
  AOI22X1 U595 ( .A(n1848), .B(n1863), .C(n1456), .D(n221), .Y(n1849) );
  OAI21X1 U598 ( .A(n1900), .B(n149), .C(n1847), .Y(n1848) );
  OAI21X1 U599 ( .A(n1937), .B(n149), .C(currentPlainKey[37]), .Y(n1847) );
  OAI21X1 U609 ( .A(n1935), .B(n149), .C(n1845), .Y(n1846) );
  OAI21X1 U610 ( .A(n1933), .B(n149), .C(currentPlainKey[36]), .Y(n1845) );
  AOI22X1 U624 ( .A(n1842), .B(n1856), .C(n1457), .D(n221), .Y(n1843) );
  OAI21X1 U627 ( .A(n1893), .B(n149), .C(n1841), .Y(n1842) );
  OAI21X1 U628 ( .A(n1926), .B(n149), .C(currentPlainKey[35]), .Y(n1841) );
  OAI21X1 U638 ( .A(n1890), .B(n149), .C(n1839), .Y(n1840) );
  OAI21X1 U639 ( .A(n1922), .B(n149), .C(currentPlainKey[34]), .Y(n1839) );
  AOI22X1 U653 ( .A(n1836), .B(n1850), .C(n1458), .D(n221), .Y(n1837) );
  OAI21X1 U658 ( .A(n1918), .B(n149), .C(n1835), .Y(n1836) );
  OAI21X1 U659 ( .A(n1916), .B(n149), .C(currentPlainKey[33]), .Y(n1835) );
  OAI21X1 U669 ( .A(n1914), .B(n149), .C(n1833), .Y(n1834) );
  OAI21X1 U670 ( .A(n1912), .B(n149), .C(currentPlainKey[32]), .Y(n1833) );
  NOR2X1 U672 ( .A(n1504), .B(address[4]), .Y(n1857) );
  AOI22X1 U686 ( .A(n1830), .B(n1844), .C(n1459), .D(n221), .Y(n1831) );
  OAI21X1 U689 ( .A(n1907), .B(n147), .C(n1829), .Y(n1830) );
  OAI21X1 U690 ( .A(n127), .B(n147), .C(currentPlainKey[31]), .Y(n1829) );
  OAI21X1 U700 ( .A(n1948), .B(n147), .C(n1827), .Y(n1828) );
  OAI21X1 U701 ( .A(n1946), .B(n147), .C(currentPlainKey[30]), .Y(n1827) );
  AOI22X1 U715 ( .A(n1824), .B(n1838), .C(n1460), .D(n221), .Y(n1825) );
  OAI21X1 U718 ( .A(n1900), .B(n147), .C(n1823), .Y(n1824) );
  OAI21X1 U719 ( .A(n1937), .B(n147), .C(currentPlainKey[29]), .Y(n1823) );
  OAI21X1 U729 ( .A(n1935), .B(n147), .C(n1821), .Y(n1822) );
  OAI21X1 U730 ( .A(n1933), .B(n147), .C(currentPlainKey[28]), .Y(n1821) );
  AOI22X1 U744 ( .A(n1818), .B(n1832), .C(n1461), .D(n221), .Y(n1819) );
  OAI21X1 U747 ( .A(n1893), .B(n147), .C(n1817), .Y(n1818) );
  OAI21X1 U748 ( .A(n1926), .B(n147), .C(currentPlainKey[27]), .Y(n1817) );
  OAI21X1 U758 ( .A(n1890), .B(n147), .C(n1815), .Y(n1816) );
  OAI21X1 U759 ( .A(n1922), .B(n147), .C(currentPlainKey[26]), .Y(n1815) );
  AOI22X1 U773 ( .A(n1812), .B(n1826), .C(n1462), .D(n221), .Y(n1813) );
  OAI21X1 U776 ( .A(n1918), .B(n147), .C(n1811), .Y(n1812) );
  OAI21X1 U777 ( .A(n1916), .B(n147), .C(currentPlainKey[25]), .Y(n1811) );
  OAI21X1 U787 ( .A(n1914), .B(n147), .C(n1809), .Y(n1810) );
  OAI21X1 U788 ( .A(n1912), .B(n147), .C(currentPlainKey[24]), .Y(n1809) );
  AOI22X1 U803 ( .A(n1805), .B(n1820), .C(n1463), .D(n221), .Y(n1806) );
  OAI21X1 U806 ( .A(n1907), .B(n145), .C(n1804), .Y(n1805) );
  OAI21X1 U807 ( .A(n127), .B(n145), .C(currentPlainKey[23]), .Y(n1804) );
  OAI21X1 U817 ( .A(n1948), .B(n145), .C(n1802), .Y(n1803) );
  OAI21X1 U818 ( .A(n1946), .B(n145), .C(currentPlainKey[22]), .Y(n1802) );
  AOI22X1 U832 ( .A(n1799), .B(n1814), .C(n1464), .D(n221), .Y(n1800) );
  OAI21X1 U835 ( .A(n1900), .B(n145), .C(n1798), .Y(n1799) );
  OAI21X1 U836 ( .A(n1937), .B(n145), .C(currentPlainKey[21]), .Y(n1798) );
  OAI21X1 U846 ( .A(n1935), .B(n145), .C(n1796), .Y(n1797) );
  OAI21X1 U847 ( .A(n1933), .B(n145), .C(currentPlainKey[20]), .Y(n1796) );
  AOI22X1 U861 ( .A(n1793), .B(n1807), .C(n1465), .D(n221), .Y(n1794) );
  OAI21X1 U864 ( .A(n1893), .B(n145), .C(n1792), .Y(n1793) );
  OAI21X1 U865 ( .A(n1926), .B(n145), .C(currentPlainKey[19]), .Y(n1792) );
  OAI21X1 U875 ( .A(n1890), .B(n145), .C(n1790), .Y(n1791) );
  OAI21X1 U876 ( .A(n1922), .B(n145), .C(currentPlainKey[18]), .Y(n1790) );
  AOI22X1 U890 ( .A(n1787), .B(n1801), .C(n1466), .D(n221), .Y(n1788) );
  OAI21X1 U895 ( .A(n1918), .B(n145), .C(n1786), .Y(n1787) );
  OAI21X1 U896 ( .A(n1916), .B(n145), .C(currentPlainKey[17]), .Y(n1786) );
  OAI21X1 U906 ( .A(n1914), .B(n145), .C(n1784), .Y(n1785) );
  OAI21X1 U907 ( .A(n1912), .B(n145), .C(currentPlainKey[16]), .Y(n1784) );
  NOR2X1 U909 ( .A(n1505), .B(address[5]), .Y(n1808) );
  AOI22X1 U923 ( .A(n1781), .B(n1795), .C(n1467), .D(n221), .Y(n1782) );
  OAI21X1 U926 ( .A(n1907), .B(n143), .C(n1780), .Y(n1781) );
  OAI21X1 U927 ( .A(n127), .B(n143), .C(currentPlainKey[15]), .Y(n1780) );
  OAI21X1 U937 ( .A(n1948), .B(n143), .C(n1778), .Y(n1779) );
  OAI21X1 U938 ( .A(n1946), .B(n143), .C(currentPlainKey[14]), .Y(n1778) );
  AOI22X1 U952 ( .A(n1775), .B(n1789), .C(n1468), .D(n221), .Y(n1776) );
  OAI21X1 U955 ( .A(n1900), .B(n143), .C(n1774), .Y(n1775) );
  OAI21X1 U956 ( .A(n1937), .B(n143), .C(currentPlainKey[13]), .Y(n1774) );
  OAI21X1 U966 ( .A(n1935), .B(n143), .C(n1772), .Y(n1773) );
  OAI21X1 U967 ( .A(n1933), .B(n143), .C(currentPlainKey[12]), .Y(n1772) );
  AOI22X1 U981 ( .A(n1769), .B(n1783), .C(n1469), .D(n221), .Y(n1770) );
  OAI21X1 U984 ( .A(n1893), .B(n143), .C(n1768), .Y(n1769) );
  OAI21X1 U985 ( .A(n1926), .B(n143), .C(currentPlainKey[11]), .Y(n1768) );
  OAI21X1 U995 ( .A(n1890), .B(n143), .C(n1766), .Y(n1767) );
  OAI21X1 U996 ( .A(n1922), .B(n143), .C(currentPlainKey[10]), .Y(n1766) );
  AOI22X1 U1010 ( .A(n1763), .B(n1777), .C(n1470), .D(n221), .Y(n1764) );
  OAI21X1 U1014 ( .A(n1918), .B(n143), .C(n1762), .Y(n1763) );
  OAI21X1 U1015 ( .A(n1916), .B(n143), .C(currentPlainKey[9]), .Y(n1762) );
  OAI21X1 U1025 ( .A(n1914), .B(n143), .C(n1760), .Y(n1761) );
  OAI21X1 U1026 ( .A(n1912), .B(n143), .C(currentPlainKey[8]), .Y(n1760) );
  AOI22X1 U1041 ( .A(n1757), .B(n1771), .C(n1471), .D(n221), .Y(n1758) );
  OAI21X1 U1044 ( .A(n1907), .B(n141), .C(n1756), .Y(n1757) );
  OAI21X1 U1045 ( .A(n127), .B(n141), .C(currentPlainKey[7]), .Y(n1756) );
  NAND2X1 U1046 ( .A(n139), .B(n7), .Y(n1907) );
  OAI21X1 U1057 ( .A(n1948), .B(n141), .C(n1753), .Y(n1754) );
  OAI21X1 U1058 ( .A(n1946), .B(n141), .C(currentPlainKey[6]), .Y(n1753) );
  NAND2X1 U1059 ( .A(n139), .B(n125), .Y(n1948) );
  AOI22X1 U1074 ( .A(n1751), .B(n1765), .C(n1472), .D(n221), .Y(n1752) );
  OAI21X1 U1077 ( .A(n1900), .B(n141), .C(n1750), .Y(n1751) );
  OAI21X1 U1078 ( .A(n1937), .B(n141), .C(currentPlainKey[5]), .Y(n1750) );
  NAND2X1 U1079 ( .A(n139), .B(n1474), .Y(n1900) );
  OAI21X1 U1090 ( .A(n1935), .B(n141), .C(n1747), .Y(n1748) );
  OAI21X1 U1091 ( .A(n1933), .B(n141), .C(currentPlainKey[4]), .Y(n1747) );
  NAND2X1 U1092 ( .A(n139), .B(n129), .Y(n1935) );
  OAI21X1 U1111 ( .A(n1893), .B(n141), .C(n1745), .Y(n1746) );
  OAI21X1 U1112 ( .A(n1926), .B(n141), .C(currentPlainKey[3]), .Y(n1745) );
  NAND2X1 U1113 ( .A(n139), .B(n1477), .Y(n1893) );
  OAI21X1 U1126 ( .A(n1890), .B(n141), .C(n1743), .Y(n1744) );
  OAI21X1 U1127 ( .A(n1922), .B(n141), .C(currentPlainKey[2]), .Y(n1743) );
  NAND2X1 U1128 ( .A(n139), .B(n131), .Y(n1890) );
  NOR2X1 U1154 ( .A(address[6]), .B(address[7]), .Y(n1885) );
  OAI21X1 U1155 ( .A(n1918), .B(n141), .C(n1741), .Y(n1742) );
  OAI21X1 U1156 ( .A(n1916), .B(n141), .C(currentPlainKey[1]), .Y(n1741) );
  NAND2X1 U1157 ( .A(n139), .B(n119), .Y(n1918) );
  AOI22X1 U1182 ( .A(n9), .B(n1572), .C(n1739), .D(n1738), .Y(n1740) );
  AOI21X1 U1183 ( .A(n1737), .B(n1749), .C(n9), .Y(n1738) );
  OAI21X1 U1184 ( .A(n222), .B(n1755), .C(n1736), .Y(n1737) );
  NAND2X1 U1185 ( .A(n16), .B(n1735), .Y(n1736) );
  OAI21X1 U1186 ( .A(n1914), .B(n141), .C(n1734), .Y(n1735) );
  OAI21X1 U1187 ( .A(n1912), .B(n141), .C(currentPlainKey[0]), .Y(n1734) );
  NOR2X1 U1189 ( .A(address[4]), .B(address[5]), .Y(n1759) );
  NAND2X1 U1190 ( .A(n139), .B(n1473), .Y(n1914) );
  AOI22X1 U1199 ( .A(n1475), .B(RCV_DATA[2]), .C(n1498), .D(RCV_DATA[3]), .Y(
        n1739) );
  NOR2X1 U1220 ( .A(n1504), .B(n1505), .Y(n1911) );
  OAI21X1 U1273 ( .A(n1476), .B(n1480), .C(n1733), .Y(n1584) );
  NAND3X1 U1274 ( .A(keyCount[0]), .B(n1480), .C(n1732), .Y(n1733) );
  NAND2X1 U1305 ( .A(n1576), .B(n1570), .Y(n1730) );
  NAND3X1 U1314 ( .A(keyCount[2]), .B(keyCount[1]), .C(n1729), .Y(n1731) );
  NOR2X1 U1315 ( .A(keyCount[3]), .B(n1479), .Y(n1729) );
  AND2X2 U254 ( .A(n1932), .B(n1963), .Y(n1939) );
  keyreg_0_DW01_add_0 r577 ( .A(parityAccumulator), .B({RCV_DATA[7:2], n221, 
        n139}), .CI(1'b0), .SUM({N1799, N1798, N1797, N1796, N1795, N1794, 
        N1793, N1792}) );
  DFFSR \state_reg[0]  ( .D(n1580), .CLK(CLK), .R(n234), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[3]  ( .D(n1579), .CLK(CLK), .R(n234), .S(1'b1), .Q(state[3]) );
  DFFSR \state_reg[2]  ( .D(n1581), .CLK(CLK), .R(n234), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[1]  ( .D(n1582), .CLK(CLK), .R(n234), .S(1'b1), .Q(state[1]) );
  DFFSR parityError_reg ( .D(nextParityError), .CLK(CLK), .R(n234), .S(1'b1), 
        .Q(parityError) );
  DFFSR PARITY_ERROR_reg ( .D(nextParityError), .CLK(CLK), .R(n234), .S(1'b1), 
        .Q(PARITY_ERROR) );
  INVX8 U3 ( .A(n154), .Y(n153) );
  INVX2 U4 ( .A(n101), .Y(n103) );
  BUFX2 U5 ( .A(n1181), .Y(n181) );
  BUFX2 U7 ( .A(n75), .Y(n188) );
  BUFX2 U8 ( .A(n1364), .Y(n203) );
  INVX2 U23 ( .A(n123), .Y(n1391) );
  BUFX2 U26 ( .A(n1367), .Y(n219) );
  INVX1 U29 ( .A(n139), .Y(n1575) );
  AND2X2 U32 ( .A(n79), .B(n1478), .Y(n1) );
  AND2X2 U35 ( .A(n81), .B(n1478), .Y(n2) );
  AND2X2 U38 ( .A(n83), .B(n1478), .Y(n4) );
  AND2X2 U41 ( .A(n6), .B(n1478), .Y(n5) );
  AND2X2 U44 ( .A(n1911), .B(n1885), .Y(n6) );
  AND2X2 U47 ( .A(n53), .B(address[0]), .Y(n7) );
  INVX2 U50 ( .A(n11), .Y(n154) );
  AND2X2 U53 ( .A(n1477), .B(address[3]), .Y(n8) );
  AND2X2 U56 ( .A(n266), .B(n19), .Y(n9) );
  AND2X2 U59 ( .A(n266), .B(n8), .Y(n10) );
  INVX2 U62 ( .A(n121), .Y(n123) );
  INVX2 U65 ( .A(state[3]), .Y(n115) );
  AND2X2 U68 ( .A(n188), .B(n1420), .Y(n11) );
  AND2X2 U71 ( .A(n1432), .B(n103), .Y(n14) );
  AND2X2 U74 ( .A(n295), .B(n1755), .Y(n16) );
  AND2X2 U77 ( .A(n131), .B(address[3]), .Y(n17) );
  AND2X2 U80 ( .A(n129), .B(address[3]), .Y(n19) );
  AND2X2 U83 ( .A(n1474), .B(address[3]), .Y(n20) );
  AND2X2 U86 ( .A(n125), .B(address[3]), .Y(n21) );
  AND2X2 U89 ( .A(n7), .B(address[3]), .Y(n23) );
  AND2X2 U92 ( .A(n1473), .B(address[3]), .Y(n25) );
  AND2X2 U95 ( .A(n313), .B(n340), .Y(n27) );
  AND2X2 U98 ( .A(n1888), .B(n1010), .Y(n29) );
  AND2X2 U101 ( .A(n1875), .B(n950), .Y(n31) );
  AND2X2 U104 ( .A(n1777), .B(n455), .Y(n33) );
  AND2X2 U107 ( .A(n1789), .B(n515), .Y(n35) );
  AND2X2 U110 ( .A(n1826), .B(n702), .Y(n37) );
  AND2X2 U113 ( .A(n1838), .B(n762), .Y(n39) );
  AND2X2 U116 ( .A(n1765), .B(n392), .Y(n41) );
  AND2X2 U119 ( .A(n1801), .B(n578), .Y(n43) );
  AND2X2 U122 ( .A(n1814), .B(n639), .Y(n45) );
  AND2X2 U125 ( .A(n1850), .B(n825), .Y(n47) );
  AND2X2 U128 ( .A(n1863), .B(n885), .Y(n49) );
  AND2X2 U131 ( .A(n1903), .B(n1069), .Y(n51) );
  AND2X2 U134 ( .A(address[1]), .B(address[2]), .Y(n53) );
  AND2X2 U137 ( .A(n1939), .B(n1936), .Y(n55) );
  AND2X2 U140 ( .A(n266), .B(n17), .Y(n57) );
  INVX1 U161 ( .A(RCV_DATA[0]), .Y(n137) );
  INVX4 U164 ( .A(n133), .Y(n1132) );
  INVX1 U167 ( .A(state[1]), .Y(n244) );
  NAND2X1 U170 ( .A(n111), .B(n14), .Y(n1425) );
  AND2X1 U173 ( .A(n249), .B(n1425), .Y(n113) );
  INVX2 U176 ( .A(n91), .Y(n71) );
  INVX4 U179 ( .A(n166), .Y(n156) );
  AND2X1 U182 ( .A(n1098), .B(n221), .Y(n73) );
  INVX8 U185 ( .A(n222), .Y(n221) );
  INVX2 U190 ( .A(n137), .Y(n139) );
  INVX2 U193 ( .A(n231), .Y(n226) );
  INVX2 U198 ( .A(n231), .Y(n225) );
  INVX2 U199 ( .A(n230), .Y(n224) );
  INVX2 U200 ( .A(n230), .Y(n223) );
  INVX2 U201 ( .A(n232), .Y(n227) );
  INVX2 U204 ( .A(n232), .Y(n228) );
  INVX2 U207 ( .A(n233), .Y(n229) );
  INVX2 U209 ( .A(n188), .Y(n187) );
  BUFX2 U212 ( .A(n234), .Y(n232) );
  BUFX2 U214 ( .A(n232), .Y(n231) );
  BUFX2 U215 ( .A(n233), .Y(n230) );
  BUFX2 U216 ( .A(n234), .Y(n233) );
  INVX2 U217 ( .A(n73), .Y(n135) );
  INVX2 U218 ( .A(n73), .Y(n133) );
  INVX2 U219 ( .A(n189), .Y(n186) );
  INVX2 U228 ( .A(n189), .Y(n185) );
  INVX2 U229 ( .A(RST), .Y(n234) );
  BUFX2 U230 ( .A(n1360), .Y(n192) );
  BUFX2 U231 ( .A(n1360), .Y(n193) );
  BUFX2 U232 ( .A(n1360), .Y(n195) );
  BUFX2 U237 ( .A(n1360), .Y(n197) );
  BUFX2 U241 ( .A(n1364), .Y(n206) );
  INVX2 U243 ( .A(n165), .Y(n160) );
  BUFX2 U244 ( .A(n1364), .Y(n205) );
  BUFX2 U245 ( .A(n1181), .Y(n183) );
  BUFX2 U246 ( .A(n1181), .Y(n180) );
  BUFX2 U247 ( .A(n1181), .Y(n178) );
  INVX2 U248 ( .A(n165), .Y(n161) );
  INVX2 U249 ( .A(n166), .Y(n158) );
  AND2X2 U250 ( .A(n264), .B(n1414), .Y(n75) );
  BUFX2 U251 ( .A(n1181), .Y(n184) );
  BUFX2 U255 ( .A(n1364), .Y(n207) );
  INVX2 U256 ( .A(n77), .Y(n141) );
  INVX2 U257 ( .A(n85), .Y(n151) );
  INVX2 U258 ( .A(n87), .Y(n145) );
  INVX2 U259 ( .A(n89), .Y(n149) );
  INVX2 U260 ( .A(n177), .Y(n173) );
  INVX2 U261 ( .A(n177), .Y(n172) );
  INVX2 U262 ( .A(n175), .Y(n168) );
  INVX2 U263 ( .A(n1158), .Y(n165) );
  INVX2 U267 ( .A(n1158), .Y(n166) );
  AND2X2 U268 ( .A(n1759), .B(n1478), .Y(n77) );
  AND2X2 U269 ( .A(n1857), .B(n1885), .Y(n79) );
  AND2X2 U272 ( .A(n1759), .B(n1885), .Y(n81) );
  AND2X2 U273 ( .A(n1808), .B(n1885), .Y(n83) );
  INVX2 U274 ( .A(n1946), .Y(n125) );
  AND2X2 U275 ( .A(n1911), .B(n1478), .Y(n85) );
  AND2X2 U276 ( .A(n1808), .B(n1478), .Y(n87) );
  AND2X2 U277 ( .A(n1857), .B(n1478), .Y(n89) );
  INVX2 U278 ( .A(n93), .Y(n143) );
  INVX2 U279 ( .A(n95), .Y(n147) );
  INVX2 U280 ( .A(n97), .Y(n150) );
  INVX2 U281 ( .A(RCV_DATA[1]), .Y(n222) );
  AND2X2 U282 ( .A(n11), .B(RCV_DATA[2]), .Y(n91) );
  INVX2 U283 ( .A(n1916), .Y(n119) );
  INVX2 U286 ( .A(n1933), .Y(n129) );
  INVX2 U288 ( .A(n1922), .Y(n131) );
  INVX2 U289 ( .A(n7), .Y(n127) );
  AND2X2 U290 ( .A(n1759), .B(address[3]), .Y(n93) );
  AND2X2 U291 ( .A(n1808), .B(address[3]), .Y(n95) );
  AND2X2 U292 ( .A(n1857), .B(address[3]), .Y(n97) );
  NAND2X1 U293 ( .A(n188), .B(n1420), .Y(n99) );
  INVX2 U294 ( .A(state[2]), .Y(n101) );
  AND2X2 U295 ( .A(n109), .B(n1413), .Y(n117) );
  BUFX2 U296 ( .A(state[0]), .Y(n105) );
  INVX1 U297 ( .A(n115), .Y(n107) );
  INVX2 U298 ( .A(n1427), .Y(n1406) );
  INVX2 U299 ( .A(state[0]), .Y(n1432) );
  NOR2X1 U301 ( .A(state[1]), .B(state[0]), .Y(n109) );
  INVX1 U302 ( .A(n109), .Y(n1408) );
  AND2X2 U305 ( .A(state[1]), .B(n115), .Y(n111) );
  INVX1 U306 ( .A(n123), .Y(n1395) );
  INVX1 U307 ( .A(n123), .Y(n1393) );
  INVX1 U308 ( .A(n123), .Y(n1399) );
  BUFX2 U309 ( .A(n91), .Y(n177) );
  BUFX2 U310 ( .A(n91), .Y(n175) );
  INVX1 U311 ( .A(n117), .Y(n1424) );
  BUFX2 U312 ( .A(n75), .Y(n189) );
  INVX1 U313 ( .A(n1426), .Y(n1384) );
  INVX2 U317 ( .A(n1403), .Y(n121) );
  INVX1 U318 ( .A(n1361), .Y(n1098) );
  BUFX4 U319 ( .A(n1367), .Y(n208) );
  BUFX4 U320 ( .A(n1367), .Y(n209) );
  BUFX4 U321 ( .A(n1367), .Y(n210) );
  BUFX4 U322 ( .A(n1367), .Y(n217) );
  NAND2X1 U323 ( .A(address[0]), .B(address[1]), .Y(n240) );
  OR2X2 U324 ( .A(address[2]), .B(n240), .Y(n1926) );
  INVX2 U325 ( .A(n1926), .Y(n1477) );
  NAND2X1 U326 ( .A(n8), .B(n6), .Y(n1963) );
  INVX2 U327 ( .A(address[2]), .Y(n262) );
  INVX2 U328 ( .A(address[1]), .Y(n261) );
  NAND3X1 U329 ( .A(address[0]), .B(n262), .C(n261), .Y(n1916) );
  NAND2X1 U331 ( .A(n119), .B(address[3]), .Y(n269) );
  INVX2 U332 ( .A(n269), .Y(n917) );
  NAND2X1 U335 ( .A(n917), .B(n6), .Y(n1967) );
  INVX2 U336 ( .A(n103), .Y(n1413) );
  NAND3X1 U337 ( .A(n111), .B(n1432), .C(n1413), .Y(n1438) );
  NAND3X1 U338 ( .A(n103), .B(n105), .C(n111), .Y(n1411) );
  NAND2X1 U339 ( .A(n1438), .B(n1411), .Y(CLR_RBUFF) );
  NAND3X1 U340 ( .A(n109), .B(n103), .C(n115), .Y(n241) );
  INVX2 U341 ( .A(n241), .Y(PROG_ERROR) );
  NAND3X1 U342 ( .A(n111), .B(n105), .C(n1413), .Y(n1427) );
  OAI21X1 U343 ( .A(n107), .B(n1424), .C(n1427), .Y(n243) );
  NAND2X1 U346 ( .A(n1425), .B(n241), .Y(n242) );
  NOR3X1 U347 ( .A(CLR_RBUFF), .B(n243), .C(n242), .Y(n1371) );
  NAND2X1 U348 ( .A(n117), .B(n107), .Y(n1426) );
  NAND3X1 U349 ( .A(n105), .B(n244), .C(n115), .Y(n245) );
  INVX2 U350 ( .A(n245), .Y(n247) );
  NAND2X1 U351 ( .A(n247), .B(n103), .Y(n1414) );
  INVX2 U352 ( .A(n1414), .Y(n1435) );
  NAND2X1 U353 ( .A(n247), .B(n1413), .Y(n249) );
  INVX2 U354 ( .A(n249), .Y(n1383) );
  AOI21X1 U355 ( .A(n1435), .B(parityError), .C(n1383), .Y(n248) );
  NAND3X1 U356 ( .A(n1371), .B(n1426), .C(n248), .Y(KEY_ERROR) );
  NOR2X1 U357 ( .A(PROG_ERROR), .B(n223), .Y(n255) );
  NAND2X1 U358 ( .A(n249), .B(n1425), .Y(n1419) );
  NOR2X1 U360 ( .A(n1406), .B(n1419), .Y(n250) );
  NAND3X1 U361 ( .A(n255), .B(n1426), .C(n250), .Y(n1403) );
  NAND2X1 U364 ( .A(n1391), .B(n1411), .Y(n1442) );
  INVX2 U365 ( .A(n1442), .Y(n264) );
  INVX2 U366 ( .A(n1438), .Y(n1420) );
  NAND2X1 U367 ( .A(n264), .B(n1420), .Y(n1444) );
  NOR2X1 U368 ( .A(n1490), .B(n1444), .Y(n1732) );
  NAND2X1 U369 ( .A(keyCount[1]), .B(keyCount[0]), .Y(n257) );
  NAND2X1 U370 ( .A(n1420), .B(n257), .Y(n258) );
  NAND2X1 U371 ( .A(n264), .B(n258), .Y(n1439) );
  INVX2 U372 ( .A(n1439), .Y(n1476) );
  INVX2 U375 ( .A(address[0]), .Y(n263) );
  NAND2X1 U376 ( .A(n53), .B(n263), .Y(n1946) );
  NAND3X1 U377 ( .A(address[6]), .B(address[7]), .C(n1911), .Y(n268) );
  INVX2 U378 ( .A(n268), .Y(n266) );
  NAND2X1 U379 ( .A(n266), .B(n21), .Y(n295) );
  INVX2 U380 ( .A(n295), .Y(n1475) );
  NAND2X1 U381 ( .A(address[0]), .B(address[2]), .Y(n259) );
  OR2X2 U382 ( .A(address[1]), .B(n259), .Y(n1937) );
  INVX2 U383 ( .A(n1937), .Y(n1474) );
  NAND2X1 U384 ( .A(n266), .B(n20), .Y(n1749) );
  INVX2 U385 ( .A(n1749), .Y(n1498) );
  NOR2X1 U386 ( .A(address[2]), .B(address[0]), .Y(n260) );
  NAND2X1 U387 ( .A(n260), .B(n261), .Y(n1912) );
  INVX2 U389 ( .A(n1912), .Y(n1473) );
  INVX2 U390 ( .A(address[3]), .Y(n1478) );
  NAND2X1 U393 ( .A(n266), .B(n23), .Y(n1755) );
  NAND3X1 U394 ( .A(address[2]), .B(n263), .C(n261), .Y(n1933) );
  INVX2 U395 ( .A(RCV_DATA[4]), .Y(n1572) );
  NAND3X1 U396 ( .A(address[1]), .B(n263), .C(n262), .Y(n1922) );
  NAND2X1 U397 ( .A(n2), .B(n129), .Y(n1765) );
  INVX2 U398 ( .A(n1765), .Y(n1472) );
  NAND2X1 U399 ( .A(n2), .B(n125), .Y(n1771) );
  INVX2 U400 ( .A(n1771), .Y(n1471) );
  NAND2X1 U401 ( .A(n81), .B(n25), .Y(n1777) );
  INVX2 U404 ( .A(n1777), .Y(n1470) );
  NAND2X1 U405 ( .A(n81), .B(n17), .Y(n1783) );
  INVX2 U406 ( .A(n1783), .Y(n1469) );
  NAND2X1 U407 ( .A(n81), .B(n19), .Y(n1789) );
  INVX2 U408 ( .A(n1789), .Y(n1468) );
  NAND2X1 U409 ( .A(n81), .B(n21), .Y(n1795) );
  INVX2 U410 ( .A(n1795), .Y(n1467) );
  NAND2X1 U411 ( .A(n4), .B(n1473), .Y(n1801) );
  INVX2 U412 ( .A(n1801), .Y(n1466) );
  NAND2X1 U413 ( .A(n4), .B(n131), .Y(n1807) );
  INVX2 U414 ( .A(n1807), .Y(n1465) );
  NAND2X1 U415 ( .A(n4), .B(n129), .Y(n1814) );
  INVX2 U416 ( .A(n1814), .Y(n1464) );
  NAND2X1 U418 ( .A(n4), .B(n125), .Y(n1820) );
  INVX2 U419 ( .A(n1820), .Y(n1463) );
  NAND2X1 U420 ( .A(n83), .B(n25), .Y(n1826) );
  INVX2 U421 ( .A(n1826), .Y(n1462) );
  NAND2X1 U424 ( .A(n83), .B(n17), .Y(n1832) );
  INVX2 U425 ( .A(n1832), .Y(n1461) );
  NAND2X1 U426 ( .A(n83), .B(n19), .Y(n1838) );
  INVX2 U427 ( .A(n1838), .Y(n1460) );
  NAND2X1 U428 ( .A(n83), .B(n21), .Y(n1844) );
  INVX2 U429 ( .A(n1844), .Y(n1459) );
  NAND2X1 U430 ( .A(n1), .B(n1473), .Y(n1850) );
  INVX2 U431 ( .A(n1850), .Y(n1458) );
  NAND2X1 U432 ( .A(n1), .B(n131), .Y(n1856) );
  INVX2 U435 ( .A(n1856), .Y(n1457) );
  NAND2X1 U436 ( .A(n1), .B(n129), .Y(n1863) );
  INVX2 U437 ( .A(n1863), .Y(n1456) );
  NAND2X1 U438 ( .A(n1), .B(n125), .Y(n1869) );
  INVX2 U439 ( .A(n1869), .Y(n1455) );
  NAND2X1 U440 ( .A(n79), .B(n25), .Y(n1875) );
  INVX2 U441 ( .A(n1875), .Y(n1454) );
  NAND2X1 U442 ( .A(n79), .B(n17), .Y(n1881) );
  INVX2 U443 ( .A(n1881), .Y(n1453) );
  NAND2X1 U444 ( .A(n19), .B(n79), .Y(n1888) );
  INVX2 U445 ( .A(n1888), .Y(n1452) );
  NAND2X1 U446 ( .A(n21), .B(n79), .Y(n1896) );
  INVX2 U447 ( .A(n1896), .Y(n1451) );
  NAND2X1 U448 ( .A(n5), .B(n1473), .Y(n1903) );
  INVX2 U450 ( .A(n1903), .Y(n1450) );
  NAND2X1 U451 ( .A(n5), .B(n131), .Y(n1910) );
  INVX2 U454 ( .A(n1910), .Y(n1449) );
  NAND2X1 U455 ( .A(n5), .B(n129), .Y(n1921) );
  INVX2 U456 ( .A(n1921), .Y(n1448) );
  NAND2X1 U457 ( .A(n5), .B(n125), .Y(n1931) );
  INVX2 U458 ( .A(n1931), .Y(n1447) );
  NAND2X1 U459 ( .A(n25), .B(n6), .Y(n1969) );
  INVX2 U460 ( .A(n1969), .Y(n1446) );
  NAND2X1 U461 ( .A(n6), .B(n17), .Y(n1966) );
  INVX2 U462 ( .A(n1966), .Y(n1445) );
  INVX2 U465 ( .A(RCV_DATA[2]), .Y(n1574) );
  INVX2 U466 ( .A(RCV_DATA[3]), .Y(n1573) );
  INVX2 U467 ( .A(RCV_DATA[5]), .Y(n1571) );
  INVX2 U468 ( .A(currentPlainKey[3]), .Y(n1566) );
  INVX2 U469 ( .A(currentPlainKey[2]), .Y(n1567) );
  INVX2 U470 ( .A(currentPlainKey[1]), .Y(n1568) );
  NAND2X1 U471 ( .A(n187), .B(currentPlainKey[0]), .Y(n277) );
  NAND2X1 U472 ( .A(n188), .B(n1420), .Y(n1361) );
  NAND2X1 U473 ( .A(n11), .B(RCV_DATA[5]), .Y(n1171) );
  OAI21X1 U474 ( .A(n10), .B(n99), .C(n1171), .Y(n265) );
  OAI21X1 U475 ( .A(n1740), .B(n10), .C(n265), .Y(n267) );
  NAND2X1 U476 ( .A(RCV_DATA[6]), .B(n11), .Y(n320) );
  MUX2X1 U477 ( .B(n267), .A(n320), .S(n57), .Y(n271) );
  NAND2X1 U479 ( .A(RCV_DATA[7]), .B(n153), .Y(n1267) );
  INVX2 U480 ( .A(n1267), .Y(n1367) );
  NOR2X1 U483 ( .A(n269), .B(n268), .Y(n270) );
  MUX2X1 U484 ( .B(n271), .A(n210), .S(n270), .Y(n275) );
  NAND2X1 U485 ( .A(n277), .B(n275), .Y(n1601) );
  NAND2X1 U486 ( .A(n185), .B(currentPlainKey[1]), .Y(n291) );
  NAND2X1 U487 ( .A(n1098), .B(RCV_DATA[3]), .Y(n1158) );
  INVX2 U488 ( .A(n1742), .Y(n278) );
  NAND2X1 U489 ( .A(n2), .B(n1473), .Y(n313) );
  INVX2 U490 ( .A(n313), .Y(n376) );
  MUX2X1 U491 ( .B(n278), .A(n222), .S(n376), .Y(n280) );
  NOR2X1 U494 ( .A(n1574), .B(n1755), .Y(n279) );
  AOI21X1 U495 ( .A(n16), .B(n280), .C(n279), .Y(n281) );
  NOR2X1 U496 ( .A(n281), .B(n1361), .Y(n282) );
  AOI21X1 U497 ( .A(n1475), .B(n165), .C(n282), .Y(n284) );
  NAND2X1 U498 ( .A(n11), .B(RCV_DATA[4]), .Y(n1169) );
  MUX2X1 U499 ( .B(n284), .A(n1169), .S(n1498), .Y(n285) );
  INVX2 U500 ( .A(n1171), .Y(n1364) );
  MUX2X1 U501 ( .B(n285), .A(n203), .S(n9), .Y(n286) );
  MUX2X1 U502 ( .B(n286), .A(n320), .S(n10), .Y(n287) );
  MUX2X1 U503 ( .B(n287), .A(n219), .S(n57), .Y(n289) );
  NAND2X1 U504 ( .A(n291), .B(n289), .Y(n1602) );
  NAND2X1 U505 ( .A(n185), .B(currentPlainKey[2]), .Y(n305) );
  NOR2X1 U506 ( .A(n1169), .B(n295), .Y(n301) );
  NAND2X1 U508 ( .A(n2), .B(n119), .Y(n340) );
  NAND2X1 U509 ( .A(n27), .B(n1098), .Y(n331) );
  INVX2 U512 ( .A(n1744), .Y(n296) );
  OAI22X1 U513 ( .A(n133), .B(n340), .C(n331), .D(n296), .Y(n298) );
  OAI22X1 U514 ( .A(n1755), .B(n156), .C(n71), .D(n313), .Y(n297) );
  AOI21X1 U515 ( .A(n16), .B(n298), .C(n297), .Y(n299) );
  MUX2X1 U516 ( .B(n299), .A(n1171), .S(n1498), .Y(n300) );
  NOR2X1 U517 ( .A(n301), .B(n300), .Y(n302) );
  MUX2X1 U518 ( .B(n302), .A(n320), .S(n9), .Y(n303) );
  MUX2X1 U519 ( .B(n303), .A(n219), .S(n10), .Y(n304) );
  NAND2X1 U520 ( .A(n305), .B(n304), .Y(n1603) );
  NAND2X1 U523 ( .A(n186), .B(currentPlainKey[3]), .Y(n327) );
  NAND2X1 U524 ( .A(n1475), .B(n203), .Y(n319) );
  INVX2 U525 ( .A(n331), .Y(n311) );
  NAND2X1 U526 ( .A(n1746), .B(n311), .Y(n312) );
  NAND2X1 U527 ( .A(n2), .B(n131), .Y(n343) );
  INVX2 U528 ( .A(n343), .Y(n422) );
  MUX2X1 U529 ( .B(n312), .A(n135), .S(n422), .Y(n315) );
  OAI22X1 U530 ( .A(n156), .B(n313), .C(n71), .D(n340), .Y(n314) );
  OAI21X1 U531 ( .A(n315), .B(n314), .C(n16), .Y(n317) );
  INVX2 U532 ( .A(n1169), .Y(n1181) );
  INVX2 U533 ( .A(n1755), .Y(n370) );
  NAND2X1 U534 ( .A(n181), .B(n370), .Y(n316) );
  NAND3X1 U535 ( .A(n319), .B(n317), .C(n316), .Y(n321) );
  INVX2 U537 ( .A(n320), .Y(n1360) );
  MUX2X1 U538 ( .B(n321), .A(n195), .S(n1498), .Y(n322) );
  MUX2X1 U541 ( .B(n322), .A(n1267), .S(n9), .Y(n324) );
  INVX2 U542 ( .A(n324), .Y(n326) );
  NAND2X1 U543 ( .A(n327), .B(n326), .Y(n1604) );
  AOI22X1 U544 ( .A(currentPlainKey[4]), .B(n186), .C(n1475), .D(n192), .Y(
        n339) );
  NAND2X1 U545 ( .A(n376), .B(n178), .Y(n336) );
  OAI22X1 U546 ( .A(n160), .B(n340), .C(n71), .D(n343), .Y(n333) );
  NAND2X1 U547 ( .A(n2), .B(n1477), .Y(n380) );
  NAND2X1 U548 ( .A(n343), .B(n380), .Y(n362) );
  INVX2 U549 ( .A(n362), .Y(n418) );
  NAND2X1 U552 ( .A(n1748), .B(n418), .Y(n330) );
  OAI22X1 U553 ( .A(n133), .B(n380), .C(n331), .D(n330), .Y(n332) );
  OAI21X1 U554 ( .A(n333), .B(n332), .C(n16), .Y(n335) );
  NAND2X1 U555 ( .A(n207), .B(n370), .Y(n334) );
  NAND3X1 U556 ( .A(n336), .B(n335), .C(n334), .Y(n337) );
  MUX2X1 U557 ( .B(n337), .A(n219), .S(n1498), .Y(n338) );
  NAND2X1 U558 ( .A(n339), .B(n338), .Y(n1605) );
  NAND2X1 U559 ( .A(n1475), .B(n219), .Y(n360) );
  INVX2 U560 ( .A(n340), .Y(n400) );
  NAND2X1 U561 ( .A(n400), .B(n178), .Y(n351) );
  NOR2X1 U562 ( .A(n160), .B(n343), .Y(n347) );
  INVX2 U563 ( .A(n1752), .Y(n344) );
  NAND3X1 U564 ( .A(n418), .B(n153), .C(n344), .Y(n345) );
  OAI21X1 U565 ( .A(n172), .B(n380), .C(n345), .Y(n346) );
  OAI21X1 U567 ( .A(n347), .B(n346), .C(n27), .Y(n350) );
  NAND2X1 U568 ( .A(n376), .B(n205), .Y(n348) );
  NAND3X1 U571 ( .A(n351), .B(n350), .C(n348), .Y(n352) );
  NAND2X1 U572 ( .A(n16), .B(n352), .Y(n357) );
  AND2X2 U573 ( .A(currentPlainKey[5]), .B(n187), .Y(n353) );
  AOI21X1 U574 ( .A(n195), .B(n370), .C(n353), .Y(n355) );
  NAND3X1 U575 ( .A(n360), .B(n357), .C(n355), .Y(n1606) );
  AOI22X1 U576 ( .A(currentPlainKey[6]), .B(n186), .C(n376), .D(n192), .Y(n375) );
  NAND2X1 U577 ( .A(n400), .B(n205), .Y(n369) );
  NAND2X1 U578 ( .A(n2), .B(n1474), .Y(n392) );
  INVX2 U579 ( .A(n392), .Y(n465) );
  NAND2X1 U582 ( .A(n465), .B(n1132), .Y(n364) );
  NAND2X1 U583 ( .A(n41), .B(n153), .Y(n394) );
  INVX2 U584 ( .A(n394), .Y(n361) );
  NAND2X1 U585 ( .A(n1754), .B(n361), .Y(n363) );
  AOI21X1 U586 ( .A(n364), .B(n363), .C(n362), .Y(n366) );
  OAI22X1 U587 ( .A(n160), .B(n380), .C(n1765), .D(n168), .Y(n365) );
  OAI21X1 U588 ( .A(n366), .B(n365), .C(n27), .Y(n368) );
  NAND2X1 U589 ( .A(n422), .B(n178), .Y(n367) );
  NAND3X1 U590 ( .A(n369), .B(n368), .C(n367), .Y(n373) );
  MUX2X1 U591 ( .B(n373), .A(n219), .S(n370), .Y(n374) );
  NAND2X1 U592 ( .A(n375), .B(n374), .Y(n1607) );
  AOI22X1 U593 ( .A(currentPlainKey[7]), .B(n186), .C(n376), .D(n208), .Y(n391) );
  NAND2X1 U594 ( .A(n422), .B(n205), .Y(n383) );
  NOR2X1 U596 ( .A(n1765), .B(n161), .Y(n378) );
  OAI22X1 U597 ( .A(n173), .B(n392), .C(n1758), .D(n394), .Y(n377) );
  OAI21X1 U600 ( .A(n378), .B(n377), .C(n418), .Y(n382) );
  INVX2 U601 ( .A(n380), .Y(n437) );
  NAND2X1 U602 ( .A(n437), .B(n178), .Y(n381) );
  NAND3X1 U603 ( .A(n383), .B(n382), .C(n381), .Y(n385) );
  NAND2X1 U604 ( .A(n27), .B(n385), .Y(n390) );
  NAND2X1 U605 ( .A(n400), .B(n197), .Y(n387) );
  NAND3X1 U606 ( .A(n391), .B(n390), .C(n387), .Y(n1608) );
  AOI22X1 U607 ( .A(currentPlainKey[8]), .B(n187), .C(n422), .D(n192), .Y(n406) );
  NAND2X1 U608 ( .A(n184), .B(n1472), .Y(n399) );
  OAI22X1 U611 ( .A(n160), .B(n392), .C(n1771), .D(n168), .Y(n396) );
  NAND2X1 U612 ( .A(n2), .B(n7), .Y(n444) );
  NAND2X1 U613 ( .A(n1771), .B(n444), .Y(n427) );
  INVX2 U614 ( .A(n427), .Y(n481) );
  NAND2X1 U615 ( .A(n1761), .B(n481), .Y(n393) );
  OAI22X1 U616 ( .A(n133), .B(n444), .C(n394), .D(n393), .Y(n395) );
  OAI21X1 U617 ( .A(n396), .B(n395), .C(n418), .Y(n398) );
  NAND2X1 U618 ( .A(n437), .B(n205), .Y(n397) );
  NAND3X1 U619 ( .A(n399), .B(n398), .C(n397), .Y(n404) );
  MUX2X1 U620 ( .B(n404), .A(n219), .S(n400), .Y(n405) );
  NAND2X1 U621 ( .A(n406), .B(n405), .Y(n1609) );
  NAND2X1 U622 ( .A(n437), .B(n197), .Y(n425) );
  NAND2X1 U623 ( .A(n465), .B(n178), .Y(n414) );
  NOR2X1 U625 ( .A(n1771), .B(n161), .Y(n411) );
  INVX2 U626 ( .A(n1764), .Y(n407) );
  NAND3X1 U629 ( .A(n481), .B(n153), .C(n407), .Y(n408) );
  OAI21X1 U630 ( .A(n173), .B(n444), .C(n408), .Y(n409) );
  OAI21X1 U631 ( .A(n411), .B(n409), .C(n41), .Y(n413) );
  NAND2X1 U632 ( .A(n206), .B(n1472), .Y(n412) );
  NAND3X1 U633 ( .A(n414), .B(n413), .C(n412), .Y(n416) );
  NAND2X1 U634 ( .A(n418), .B(n416), .Y(n424) );
  AND2X2 U635 ( .A(currentPlainKey[9]), .B(n187), .Y(n419) );
  AOI21X1 U636 ( .A(n422), .B(n209), .C(n419), .Y(n423) );
  NAND3X1 U637 ( .A(n425), .B(n424), .C(n423), .Y(n1610) );
  AOI22X1 U640 ( .A(currentPlainKey[10]), .B(n185), .C(n192), .D(n1472), .Y(
        n440) );
  NAND2X1 U641 ( .A(n184), .B(n1471), .Y(n436) );
  NAND2X1 U642 ( .A(n81), .B(n917), .Y(n455) );
  INVX2 U643 ( .A(n455), .Y(n526) );
  NAND2X1 U644 ( .A(n526), .B(n1132), .Y(n429) );
  NAND2X1 U645 ( .A(n33), .B(n153), .Y(n457) );
  INVX2 U646 ( .A(n457), .Y(n426) );
  NAND2X1 U647 ( .A(n1767), .B(n426), .Y(n428) );
  AOI21X1 U648 ( .A(n429), .B(n428), .C(n427), .Y(n431) );
  OAI22X1 U649 ( .A(n160), .B(n444), .C(n1777), .D(n168), .Y(n430) );
  OAI21X1 U650 ( .A(n431), .B(n430), .C(n41), .Y(n435) );
  NAND2X1 U651 ( .A(n465), .B(n205), .Y(n432) );
  NAND3X1 U652 ( .A(n436), .B(n435), .C(n432), .Y(n438) );
  MUX2X1 U654 ( .B(n438), .A(n219), .S(n437), .Y(n439) );
  NAND2X1 U655 ( .A(n440), .B(n439), .Y(n1611) );
  AOI22X1 U656 ( .A(currentPlainKey[11]), .B(n186), .C(n208), .D(n1472), .Y(
        n454) );
  NAND2X1 U657 ( .A(n206), .B(n1471), .Y(n448) );
  NOR2X1 U660 ( .A(n1777), .B(n161), .Y(n443) );
  OAI22X1 U661 ( .A(n173), .B(n455), .C(n1770), .D(n457), .Y(n441) );
  OAI21X1 U662 ( .A(n443), .B(n441), .C(n481), .Y(n446) );
  INVX2 U663 ( .A(n444), .Y(n498) );
  NAND2X1 U664 ( .A(n498), .B(n178), .Y(n445) );
  NAND3X1 U665 ( .A(n448), .B(n446), .C(n445), .Y(n450) );
  NAND2X1 U666 ( .A(n41), .B(n450), .Y(n453) );
  NAND2X1 U667 ( .A(n465), .B(n197), .Y(n452) );
  NAND3X1 U668 ( .A(n454), .B(n453), .C(n452), .Y(n1612) );
  AOI22X1 U671 ( .A(currentPlainKey[12]), .B(n186), .C(n192), .D(n1471), .Y(
        n468) );
  NAND2X1 U673 ( .A(n184), .B(n1470), .Y(n462) );
  OAI22X1 U674 ( .A(n158), .B(n455), .C(n1783), .D(n168), .Y(n459) );
  NAND2X1 U675 ( .A(n81), .B(n8), .Y(n507) );
  NAND2X1 U676 ( .A(n1783), .B(n507), .Y(n487) );
  INVX2 U677 ( .A(n487), .Y(n541) );
  NAND2X1 U678 ( .A(n1773), .B(n541), .Y(n456) );
  OAI22X1 U679 ( .A(n133), .B(n507), .C(n457), .D(n456), .Y(n458) );
  OAI21X1 U680 ( .A(n459), .B(n458), .C(n481), .Y(n461) );
  NAND2X1 U681 ( .A(n498), .B(n205), .Y(n460) );
  NAND3X1 U682 ( .A(n462), .B(n461), .C(n460), .Y(n466) );
  MUX2X1 U683 ( .B(n466), .A(n219), .S(n465), .Y(n467) );
  NAND2X1 U684 ( .A(n468), .B(n467), .Y(n1613) );
  NAND2X1 U685 ( .A(n498), .B(n197), .Y(n485) );
  NAND2X1 U687 ( .A(n526), .B(n178), .Y(n479) );
  NOR2X1 U688 ( .A(n1783), .B(n161), .Y(n473) );
  INVX2 U691 ( .A(n1776), .Y(n469) );
  NAND3X1 U692 ( .A(n541), .B(n153), .C(n469), .Y(n471) );
  OAI21X1 U693 ( .A(n173), .B(n507), .C(n471), .Y(n472) );
  OAI21X1 U694 ( .A(n473), .B(n472), .C(n33), .Y(n476) );
  NAND2X1 U695 ( .A(n206), .B(n1470), .Y(n474) );
  NAND3X1 U696 ( .A(n479), .B(n476), .C(n474), .Y(n480) );
  NAND2X1 U697 ( .A(n481), .B(n480), .Y(n484) );
  AND2X2 U698 ( .A(currentPlainKey[13]), .B(n185), .Y(n482) );
  AOI21X1 U699 ( .A(n209), .B(n1471), .C(n482), .Y(n483) );
  NAND3X1 U702 ( .A(n485), .B(n484), .C(n483), .Y(n1614) );
  AOI22X1 U703 ( .A(currentPlainKey[14]), .B(n187), .C(n192), .D(n1470), .Y(
        n501) );
  NAND2X1 U704 ( .A(n184), .B(n1469), .Y(n496) );
  NAND2X1 U705 ( .A(n81), .B(n20), .Y(n515) );
  INVX2 U706 ( .A(n515), .Y(n590) );
  NAND2X1 U707 ( .A(n590), .B(n1132), .Y(n489) );
  NAND2X1 U708 ( .A(n35), .B(n153), .Y(n519) );
  INVX2 U709 ( .A(n519), .Y(n486) );
  NAND2X1 U710 ( .A(n1779), .B(n486), .Y(n488) );
  AOI21X1 U711 ( .A(n489), .B(n488), .C(n487), .Y(n493) );
  OAI22X1 U712 ( .A(n158), .B(n507), .C(n1789), .D(n168), .Y(n492) );
  OAI21X1 U713 ( .A(n493), .B(n492), .C(n33), .Y(n495) );
  NAND2X1 U714 ( .A(n526), .B(n205), .Y(n494) );
  NAND3X1 U716 ( .A(n496), .B(n495), .C(n494), .Y(n499) );
  MUX2X1 U717 ( .B(n499), .A(n219), .S(n498), .Y(n500) );
  NAND2X1 U720 ( .A(n501), .B(n500), .Y(n1615) );
  AOI22X1 U721 ( .A(currentPlainKey[15]), .B(n186), .C(n208), .D(n1470), .Y(
        n514) );
  NAND2X1 U722 ( .A(n206), .B(n1469), .Y(n510) );
  NOR2X1 U723 ( .A(n1789), .B(n160), .Y(n506) );
  OAI22X1 U724 ( .A(n173), .B(n515), .C(n1782), .D(n519), .Y(n503) );
  OAI21X1 U725 ( .A(n506), .B(n503), .C(n541), .Y(n509) );
  INVX2 U726 ( .A(n507), .Y(n561) );
  NAND2X1 U727 ( .A(n561), .B(n178), .Y(n508) );
  NAND3X1 U728 ( .A(n510), .B(n509), .C(n508), .Y(n511) );
  NAND2X1 U731 ( .A(n33), .B(n511), .Y(n513) );
  NAND2X1 U732 ( .A(n526), .B(n197), .Y(n512) );
  NAND3X1 U733 ( .A(n514), .B(n513), .C(n512), .Y(n1616) );
  AOI22X1 U734 ( .A(currentPlainKey[16]), .B(n186), .C(n193), .D(n1469), .Y(
        n530) );
  NAND2X1 U735 ( .A(n184), .B(n1468), .Y(n525) );
  OAI22X1 U736 ( .A(n158), .B(n515), .C(n1795), .D(n172), .Y(n521) );
  NAND2X1 U737 ( .A(n81), .B(n23), .Y(n568) );
  NAND2X1 U738 ( .A(n1795), .B(n568), .Y(n550) );
  INVX2 U739 ( .A(n550), .Y(n604) );
  NAND2X1 U740 ( .A(n1785), .B(n604), .Y(n516) );
  OAI22X1 U741 ( .A(n135), .B(n568), .C(n519), .D(n516), .Y(n520) );
  OAI21X1 U742 ( .A(n521), .B(n520), .C(n541), .Y(n523) );
  NAND2X1 U743 ( .A(n561), .B(n205), .Y(n522) );
  NAND3X1 U745 ( .A(n525), .B(n523), .C(n522), .Y(n527) );
  MUX2X1 U746 ( .B(n527), .A(n219), .S(n526), .Y(n528) );
  NAND2X1 U749 ( .A(n530), .B(n528), .Y(n1617) );
  NAND2X1 U750 ( .A(n561), .B(n197), .Y(n548) );
  NAND2X1 U751 ( .A(n590), .B(n178), .Y(n539) );
  NOR2X1 U752 ( .A(n1795), .B(n160), .Y(n536) );
  INVX2 U753 ( .A(n1788), .Y(n533) );
  NAND3X1 U754 ( .A(n604), .B(n153), .C(n533), .Y(n534) );
  OAI21X1 U755 ( .A(n173), .B(n568), .C(n534), .Y(n535) );
  OAI21X1 U756 ( .A(n536), .B(n535), .C(n35), .Y(n538) );
  NAND2X1 U757 ( .A(n206), .B(n1468), .Y(n537) );
  NAND3X1 U760 ( .A(n539), .B(n538), .C(n537), .Y(n540) );
  NAND2X1 U761 ( .A(n541), .B(n540), .Y(n547) );
  AND2X2 U762 ( .A(currentPlainKey[17]), .B(n186), .Y(n542) );
  AOI21X1 U763 ( .A(n209), .B(n1469), .C(n542), .Y(n543) );
  NAND3X1 U764 ( .A(n548), .B(n547), .C(n543), .Y(n1618) );
  AOI22X1 U765 ( .A(currentPlainKey[18]), .B(n186), .C(n192), .D(n1468), .Y(
        n565) );
  NAND2X1 U766 ( .A(n184), .B(n1467), .Y(n559) );
  NAND2X1 U767 ( .A(n4), .B(n119), .Y(n578) );
  INVX2 U768 ( .A(n578), .Y(n650) );
  NAND2X1 U769 ( .A(n650), .B(n1132), .Y(n552) );
  NAND2X1 U770 ( .A(n43), .B(n153), .Y(n580) );
  INVX2 U771 ( .A(n580), .Y(n549) );
  NAND2X1 U772 ( .A(n1791), .B(n549), .Y(n551) );
  AOI21X1 U774 ( .A(n552), .B(n551), .C(n550), .Y(n555) );
  OAI22X1 U775 ( .A(n158), .B(n568), .C(n1801), .D(n168), .Y(n554) );
  OAI21X1 U778 ( .A(n555), .B(n554), .C(n35), .Y(n557) );
  NAND2X1 U779 ( .A(n590), .B(n205), .Y(n556) );
  NAND3X1 U780 ( .A(n559), .B(n557), .C(n556), .Y(n563) );
  MUX2X1 U781 ( .B(n563), .A(n217), .S(n561), .Y(n564) );
  NAND2X1 U782 ( .A(n565), .B(n564), .Y(n1619) );
  AOI22X1 U783 ( .A(currentPlainKey[19]), .B(n186), .C(n208), .D(n1468), .Y(
        n577) );
  NAND2X1 U784 ( .A(n206), .B(n1467), .Y(n571) );
  NOR2X1 U785 ( .A(n1801), .B(n160), .Y(n567) );
  OAI22X1 U786 ( .A(n71), .B(n578), .C(n1794), .D(n580), .Y(n566) );
  OAI21X1 U789 ( .A(n567), .B(n566), .C(n604), .Y(n570) );
  INVX2 U790 ( .A(n568), .Y(n622) );
  NAND2X1 U791 ( .A(n622), .B(n180), .Y(n569) );
  NAND3X1 U792 ( .A(n571), .B(n570), .C(n569), .Y(n572) );
  NAND2X1 U793 ( .A(n35), .B(n572), .Y(n576) );
  NAND2X1 U794 ( .A(n590), .B(n197), .Y(n573) );
  NAND3X1 U795 ( .A(n577), .B(n576), .C(n573), .Y(n1620) );
  AOI22X1 U796 ( .A(currentPlainKey[20]), .B(n186), .C(n193), .D(n1467), .Y(
        n593) );
  NAND2X1 U797 ( .A(n184), .B(n1466), .Y(n587) );
  OAI22X1 U798 ( .A(n158), .B(n578), .C(n1807), .D(n172), .Y(n583) );
  NAND2X1 U799 ( .A(n4), .B(n1477), .Y(n630) );
  NAND2X1 U800 ( .A(n1807), .B(n630), .Y(n611) );
  INVX2 U801 ( .A(n611), .Y(n665) );
  NAND2X1 U802 ( .A(n1797), .B(n665), .Y(n579) );
  OAI22X1 U804 ( .A(n135), .B(n630), .C(n580), .D(n579), .Y(n582) );
  OAI21X1 U805 ( .A(n583), .B(n582), .C(n604), .Y(n585) );
  NAND2X1 U808 ( .A(n622), .B(n205), .Y(n584) );
  NAND3X1 U809 ( .A(n587), .B(n585), .C(n584), .Y(n591) );
  MUX2X1 U810 ( .B(n591), .A(n217), .S(n590), .Y(n592) );
  NAND2X1 U811 ( .A(n593), .B(n592), .Y(n1621) );
  NAND2X1 U812 ( .A(n622), .B(n197), .Y(n609) );
  NAND2X1 U813 ( .A(n650), .B(n180), .Y(n600) );
  NOR2X1 U814 ( .A(n1807), .B(n160), .Y(n597) );
  INVX2 U815 ( .A(n1800), .Y(n594) );
  NAND3X1 U816 ( .A(n665), .B(n153), .C(n594), .Y(n595) );
  OAI21X1 U819 ( .A(n173), .B(n630), .C(n595), .Y(n596) );
  OAI21X1 U820 ( .A(n597), .B(n596), .C(n43), .Y(n599) );
  NAND2X1 U821 ( .A(n205), .B(n1466), .Y(n598) );
  NAND3X1 U822 ( .A(n600), .B(n599), .C(n598), .Y(n603) );
  NAND2X1 U823 ( .A(n604), .B(n603), .Y(n607) );
  AND2X2 U824 ( .A(currentPlainKey[21]), .B(n187), .Y(n605) );
  AOI21X1 U825 ( .A(n209), .B(n1467), .C(n605), .Y(n606) );
  NAND3X1 U826 ( .A(n609), .B(n607), .C(n606), .Y(n1622) );
  AOI22X1 U827 ( .A(currentPlainKey[22]), .B(n186), .C(n193), .D(n1466), .Y(
        n625) );
  NAND2X1 U828 ( .A(n183), .B(n1465), .Y(n621) );
  NAND2X1 U829 ( .A(n4), .B(n1474), .Y(n639) );
  INVX2 U830 ( .A(n639), .Y(n710) );
  NAND2X1 U831 ( .A(n710), .B(n1132), .Y(n614) );
  NAND2X1 U833 ( .A(n45), .B(n153), .Y(n644) );
  INVX2 U834 ( .A(n644), .Y(n610) );
  NAND2X1 U837 ( .A(n1803), .B(n610), .Y(n612) );
  AOI21X1 U838 ( .A(n614), .B(n612), .C(n611), .Y(n618) );
  OAI22X1 U839 ( .A(n158), .B(n630), .C(n1814), .D(n172), .Y(n617) );
  OAI21X1 U840 ( .A(n618), .B(n617), .C(n43), .Y(n620) );
  NAND2X1 U841 ( .A(n650), .B(n205), .Y(n619) );
  NAND3X1 U842 ( .A(n621), .B(n620), .C(n619), .Y(n623) );
  MUX2X1 U843 ( .B(n623), .A(n217), .S(n622), .Y(n624) );
  NAND2X1 U844 ( .A(n625), .B(n624), .Y(n1623) );
  AOI22X1 U845 ( .A(currentPlainKey[23]), .B(n186), .C(n208), .D(n1466), .Y(
        n638) );
  NAND2X1 U848 ( .A(n205), .B(n1465), .Y(n633) );
  NOR2X1 U849 ( .A(n1814), .B(n160), .Y(n627) );
  OAI22X1 U850 ( .A(n71), .B(n639), .C(n1806), .D(n644), .Y(n626) );
  OAI21X1 U851 ( .A(n627), .B(n626), .C(n665), .Y(n632) );
  INVX2 U852 ( .A(n630), .Y(n682) );
  NAND2X1 U853 ( .A(n682), .B(n180), .Y(n631) );
  NAND3X1 U854 ( .A(n633), .B(n632), .C(n631), .Y(n634) );
  NAND2X1 U855 ( .A(n43), .B(n634), .Y(n637) );
  NAND2X1 U856 ( .A(n650), .B(n197), .Y(n636) );
  NAND3X1 U857 ( .A(n638), .B(n637), .C(n636), .Y(n1624) );
  AOI22X1 U858 ( .A(currentPlainKey[24]), .B(n186), .C(n193), .D(n1465), .Y(
        n653) );
  NAND2X1 U859 ( .A(n183), .B(n1464), .Y(n649) );
  OAI22X1 U860 ( .A(n158), .B(n639), .C(n1820), .D(n172), .Y(n646) );
  NAND2X1 U862 ( .A(n4), .B(n7), .Y(n690) );
  NAND2X1 U863 ( .A(n1820), .B(n690), .Y(n674) );
  INVX2 U866 ( .A(n674), .Y(n728) );
  NAND2X1 U867 ( .A(n1810), .B(n728), .Y(n641) );
  OAI22X1 U868 ( .A(n135), .B(n690), .C(n644), .D(n641), .Y(n645) );
  OAI21X1 U869 ( .A(n646), .B(n645), .C(n665), .Y(n648) );
  NAND2X1 U870 ( .A(n682), .B(n205), .Y(n647) );
  NAND3X1 U871 ( .A(n649), .B(n648), .C(n647), .Y(n651) );
  MUX2X1 U872 ( .B(n651), .A(n217), .S(n650), .Y(n652) );
  NAND2X1 U873 ( .A(n653), .B(n652), .Y(n1625) );
  NAND2X1 U874 ( .A(n682), .B(n195), .Y(n670) );
  NAND2X1 U877 ( .A(n710), .B(n180), .Y(n662) );
  NOR2X1 U878 ( .A(n1820), .B(n160), .Y(n659) );
  INVX2 U879 ( .A(n1813), .Y(n654) );
  NAND3X1 U880 ( .A(n728), .B(n153), .C(n654), .Y(n657) );
  OAI21X1 U881 ( .A(n173), .B(n690), .C(n657), .Y(n658) );
  OAI21X1 U882 ( .A(n659), .B(n658), .C(n45), .Y(n661) );
  NAND2X1 U883 ( .A(n206), .B(n1464), .Y(n660) );
  NAND3X1 U884 ( .A(n662), .B(n661), .C(n660), .Y(n663) );
  NAND2X1 U885 ( .A(n665), .B(n663), .Y(n668) );
  AND2X2 U886 ( .A(currentPlainKey[25]), .B(n187), .Y(n666) );
  AOI21X1 U887 ( .A(n209), .B(n1465), .C(n666), .Y(n667) );
  NAND3X1 U888 ( .A(n670), .B(n668), .C(n667), .Y(n1626) );
  AOI22X1 U889 ( .A(currentPlainKey[26]), .B(n186), .C(n193), .D(n1464), .Y(
        n687) );
  NAND2X1 U891 ( .A(n183), .B(n1463), .Y(n681) );
  NAND2X1 U892 ( .A(n83), .B(n917), .Y(n702) );
  INVX2 U893 ( .A(n702), .Y(n773) );
  NAND2X1 U894 ( .A(n773), .B(n1132), .Y(n676) );
  NAND2X1 U897 ( .A(n37), .B(n153), .Y(n704) );
  INVX2 U898 ( .A(n704), .Y(n672) );
  NAND2X1 U899 ( .A(n1816), .B(n672), .Y(n675) );
  AOI21X1 U900 ( .A(n676), .B(n675), .C(n674), .Y(n678) );
  OAI22X1 U901 ( .A(n158), .B(n690), .C(n1826), .D(n172), .Y(n677) );
  OAI21X1 U902 ( .A(n678), .B(n677), .C(n45), .Y(n680) );
  NAND2X1 U903 ( .A(n710), .B(n205), .Y(n679) );
  NAND3X1 U904 ( .A(n681), .B(n680), .C(n679), .Y(n683) );
  MUX2X1 U905 ( .B(n683), .A(n217), .S(n682), .Y(n684) );
  NAND2X1 U908 ( .A(n687), .B(n684), .Y(n1627) );
  AOI22X1 U910 ( .A(currentPlainKey[27]), .B(n186), .C(n208), .D(n1464), .Y(
        n701) );
  NAND2X1 U911 ( .A(n206), .B(n1463), .Y(n694) );
  NOR2X1 U912 ( .A(n1826), .B(n161), .Y(n689) );
  OAI22X1 U913 ( .A(n71), .B(n702), .C(n1819), .D(n704), .Y(n688) );
  OAI21X1 U914 ( .A(n689), .B(n688), .C(n728), .Y(n693) );
  INVX2 U915 ( .A(n690), .Y(n744) );
  NAND2X1 U916 ( .A(n744), .B(n178), .Y(n691) );
  NAND3X1 U917 ( .A(n694), .B(n693), .C(n691), .Y(n695) );
  NAND2X1 U918 ( .A(n45), .B(n695), .Y(n698) );
  NAND2X1 U919 ( .A(n710), .B(n195), .Y(n696) );
  NAND3X1 U920 ( .A(n701), .B(n698), .C(n696), .Y(n1628) );
  AOI22X1 U921 ( .A(currentPlainKey[28]), .B(n185), .C(n193), .D(n1463), .Y(
        n715) );
  NAND2X1 U922 ( .A(n183), .B(n1462), .Y(n709) );
  OAI22X1 U924 ( .A(n158), .B(n702), .C(n1832), .D(n172), .Y(n706) );
  NAND2X1 U925 ( .A(n83), .B(n8), .Y(n752) );
  NAND2X1 U928 ( .A(n1832), .B(n752), .Y(n734) );
  INVX2 U929 ( .A(n734), .Y(n789) );
  NAND2X1 U930 ( .A(n1822), .B(n789), .Y(n703) );
  OAI22X1 U931 ( .A(n135), .B(n752), .C(n704), .D(n703), .Y(n705) );
  OAI21X1 U932 ( .A(n706), .B(n705), .C(n728), .Y(n708) );
  NAND2X1 U933 ( .A(n744), .B(n205), .Y(n707) );
  NAND3X1 U934 ( .A(n709), .B(n708), .C(n707), .Y(n711) );
  MUX2X1 U935 ( .B(n711), .A(n217), .S(n710), .Y(n714) );
  NAND2X1 U936 ( .A(n715), .B(n714), .Y(n1629) );
  NAND2X1 U939 ( .A(n744), .B(n195), .Y(n732) );
  NAND2X1 U940 ( .A(n773), .B(n180), .Y(n723) );
  NOR2X1 U941 ( .A(n1832), .B(n160), .Y(n720) );
  INVX2 U942 ( .A(n1825), .Y(n716) );
  NAND3X1 U943 ( .A(n789), .B(n153), .C(n716), .Y(n717) );
  OAI21X1 U944 ( .A(n173), .B(n752), .C(n717), .Y(n718) );
  OAI21X1 U945 ( .A(n720), .B(n718), .C(n37), .Y(n722) );
  NAND2X1 U946 ( .A(n205), .B(n1462), .Y(n721) );
  NAND3X1 U947 ( .A(n723), .B(n722), .C(n721), .Y(n725) );
  NAND2X1 U948 ( .A(n728), .B(n725), .Y(n731) );
  AND2X2 U949 ( .A(currentPlainKey[29]), .B(n187), .Y(n729) );
  AOI21X1 U950 ( .A(n209), .B(n1463), .C(n729), .Y(n730) );
  NAND3X1 U951 ( .A(n732), .B(n731), .C(n730), .Y(n1630) );
  AOI22X1 U953 ( .A(currentPlainKey[30]), .B(n185), .C(n195), .D(n1462), .Y(
        n748) );
  NAND2X1 U954 ( .A(n183), .B(n1461), .Y(n743) );
  NAND2X1 U957 ( .A(n83), .B(n20), .Y(n762) );
  INVX2 U958 ( .A(n762), .Y(n834) );
  NAND2X1 U959 ( .A(n834), .B(n1132), .Y(n736) );
  NAND2X1 U960 ( .A(n39), .B(n153), .Y(n764) );
  INVX2 U961 ( .A(n764), .Y(n733) );
  NAND2X1 U962 ( .A(n1828), .B(n733), .Y(n735) );
  AOI21X1 U963 ( .A(n736), .B(n735), .C(n734), .Y(n738) );
  OAI22X1 U964 ( .A(n158), .B(n752), .C(n1838), .D(n71), .Y(n737) );
  OAI21X1 U965 ( .A(n738), .B(n737), .C(n37), .Y(n742) );
  NAND2X1 U968 ( .A(n773), .B(n203), .Y(n741) );
  NAND3X1 U969 ( .A(n743), .B(n742), .C(n741), .Y(n745) );
  MUX2X1 U970 ( .B(n745), .A(n217), .S(n744), .Y(n747) );
  NAND2X1 U971 ( .A(n748), .B(n747), .Y(n1631) );
  AOI22X1 U972 ( .A(currentPlainKey[31]), .B(n185), .C(n208), .D(n1462), .Y(
        n761) );
  NAND2X1 U973 ( .A(n206), .B(n1461), .Y(n757) );
  NOR2X1 U974 ( .A(n1838), .B(n160), .Y(n750) );
  OAI22X1 U975 ( .A(n71), .B(n762), .C(n1831), .D(n764), .Y(n749) );
  OAI21X1 U976 ( .A(n750), .B(n749), .C(n789), .Y(n756) );
  INVX2 U977 ( .A(n752), .Y(n806) );
  NAND2X1 U978 ( .A(n806), .B(n181), .Y(n755) );
  NAND3X1 U979 ( .A(n757), .B(n756), .C(n755), .Y(n758) );
  NAND2X1 U980 ( .A(n37), .B(n758), .Y(n760) );
  NAND2X1 U982 ( .A(n773), .B(n195), .Y(n759) );
  NAND3X1 U983 ( .A(n761), .B(n760), .C(n759), .Y(n1632) );
  AOI22X1 U986 ( .A(currentPlainKey[32]), .B(n185), .C(n195), .D(n1461), .Y(
        n777) );
  NAND2X1 U987 ( .A(n183), .B(n1460), .Y(n772) );
  OAI22X1 U988 ( .A(n158), .B(n762), .C(n1844), .D(n172), .Y(n769) );
  NAND2X1 U989 ( .A(n83), .B(n23), .Y(n815) );
  NAND2X1 U990 ( .A(n1844), .B(n815), .Y(n795) );
  INVX2 U991 ( .A(n795), .Y(n849) );
  NAND2X1 U992 ( .A(n1834), .B(n849), .Y(n763) );
  OAI22X1 U993 ( .A(n135), .B(n815), .C(n764), .D(n763), .Y(n765) );
  OAI21X1 U994 ( .A(n769), .B(n765), .C(n789), .Y(n771) );
  NAND2X1 U997 ( .A(n806), .B(n203), .Y(n770) );
  NAND3X1 U998 ( .A(n772), .B(n771), .C(n770), .Y(n774) );
  MUX2X1 U999 ( .B(n774), .A(n217), .S(n773), .Y(n776) );
  NAND2X1 U1000 ( .A(n777), .B(n776), .Y(n1633) );
  NAND2X1 U1001 ( .A(n806), .B(n195), .Y(n793) );
  NAND2X1 U1002 ( .A(n834), .B(n181), .Y(n787) );
  NOR2X1 U1003 ( .A(n1844), .B(n160), .Y(n783) );
  INVX2 U1004 ( .A(n1837), .Y(n778) );
  NAND3X1 U1005 ( .A(n849), .B(n153), .C(n778), .Y(n779) );
  OAI21X1 U1006 ( .A(n173), .B(n815), .C(n779), .Y(n781) );
  OAI21X1 U1007 ( .A(n783), .B(n781), .C(n39), .Y(n786) );
  NAND2X1 U1008 ( .A(n206), .B(n1460), .Y(n785) );
  NAND3X1 U1009 ( .A(n787), .B(n786), .C(n785), .Y(n788) );
  NAND2X1 U1011 ( .A(n789), .B(n788), .Y(n792) );
  AND2X2 U1012 ( .A(currentPlainKey[33]), .B(n187), .Y(n790) );
  AOI21X1 U1013 ( .A(n209), .B(n1461), .C(n790), .Y(n791) );
  NAND3X1 U1016 ( .A(n793), .B(n792), .C(n791), .Y(n1634) );
  AOI22X1 U1017 ( .A(currentPlainKey[34]), .B(n185), .C(n193), .D(n1460), .Y(
        n812) );
  NAND2X1 U1018 ( .A(n183), .B(n1459), .Y(n805) );
  NAND2X1 U1019 ( .A(n1), .B(n119), .Y(n825) );
  INVX2 U1020 ( .A(n825), .Y(n897) );
  NAND2X1 U1021 ( .A(n897), .B(n1132), .Y(n799) );
  NAND2X1 U1022 ( .A(n47), .B(n153), .Y(n827) );
  INVX2 U1023 ( .A(n827), .Y(n794) );
  NAND2X1 U1024 ( .A(n1840), .B(n794), .Y(n798) );
  AOI21X1 U1027 ( .A(n799), .B(n798), .C(n795), .Y(n801) );
  OAI22X1 U1028 ( .A(n158), .B(n815), .C(n1850), .D(n172), .Y(n800) );
  OAI21X1 U1029 ( .A(n801), .B(n800), .C(n39), .Y(n804) );
  NAND2X1 U1030 ( .A(n834), .B(n203), .Y(n802) );
  NAND3X1 U1031 ( .A(n805), .B(n804), .C(n802), .Y(n807) );
  MUX2X1 U1032 ( .B(n807), .A(n217), .S(n806), .Y(n809) );
  NAND2X1 U1033 ( .A(n812), .B(n809), .Y(n1635) );
  AOI22X1 U1034 ( .A(currentPlainKey[35]), .B(n185), .C(n209), .D(n1460), .Y(
        n822) );
  NAND2X1 U1035 ( .A(n206), .B(n1459), .Y(n818) );
  NOR2X1 U1036 ( .A(n1850), .B(n160), .Y(n814) );
  OAI22X1 U1037 ( .A(n71), .B(n825), .C(n1843), .D(n827), .Y(n813) );
  OAI21X1 U1038 ( .A(n814), .B(n813), .C(n849), .Y(n817) );
  INVX2 U1039 ( .A(n815), .Y(n869) );
  NAND2X1 U1040 ( .A(n869), .B(n180), .Y(n816) );
  NAND3X1 U1042 ( .A(n818), .B(n817), .C(n816), .Y(n819) );
  NAND2X1 U1043 ( .A(n39), .B(n819), .Y(n821) );
  NAND2X1 U1047 ( .A(n834), .B(n195), .Y(n820) );
  NAND3X1 U1048 ( .A(n822), .B(n821), .C(n820), .Y(n1636) );
  AOI22X1 U1049 ( .A(currentPlainKey[36]), .B(n185), .C(n195), .D(n1459), .Y(
        n840) );
  NAND2X1 U1050 ( .A(n183), .B(n1458), .Y(n833) );
  OAI22X1 U1051 ( .A(n156), .B(n825), .C(n1856), .D(n172), .Y(n829) );
  NAND2X1 U1052 ( .A(n1), .B(n1477), .Y(n875) );
  NAND2X1 U1053 ( .A(n1856), .B(n875), .Y(n858) );
  INVX2 U1054 ( .A(n858), .Y(n911) );
  NAND2X1 U1055 ( .A(n1846), .B(n911), .Y(n826) );
  OAI22X1 U1056 ( .A(n135), .B(n875), .C(n827), .D(n826), .Y(n828) );
  OAI21X1 U1060 ( .A(n829), .B(n828), .C(n849), .Y(n832) );
  NAND2X1 U1061 ( .A(n869), .B(n203), .Y(n831) );
  NAND3X1 U1062 ( .A(n833), .B(n832), .C(n831), .Y(n836) );
  MUX2X1 U1063 ( .B(n836), .A(n217), .S(n834), .Y(n839) );
  NAND2X1 U1064 ( .A(n840), .B(n839), .Y(n1637) );
  NAND2X1 U1065 ( .A(n869), .B(n195), .Y(n855) );
  NAND2X1 U1066 ( .A(n897), .B(n181), .Y(n847) );
  NOR2X1 U1067 ( .A(n1856), .B(n161), .Y(n844) );
  INVX2 U1068 ( .A(n1849), .Y(n841) );
  NAND3X1 U1069 ( .A(n911), .B(n153), .C(n841), .Y(n842) );
  OAI21X1 U1070 ( .A(n168), .B(n875), .C(n842), .Y(n843) );
  OAI21X1 U1071 ( .A(n844), .B(n843), .C(n47), .Y(n846) );
  NAND2X1 U1072 ( .A(n206), .B(n1458), .Y(n845) );
  NAND3X1 U1073 ( .A(n847), .B(n846), .C(n845), .Y(n848) );
  NAND2X1 U1075 ( .A(n849), .B(n848), .Y(n854) );
  AND2X2 U1076 ( .A(currentPlainKey[37]), .B(n186), .Y(n852) );
  AOI21X1 U1080 ( .A(n210), .B(n1459), .C(n852), .Y(n853) );
  NAND3X1 U1081 ( .A(n855), .B(n854), .C(n853), .Y(n1638) );
  AOI22X1 U1082 ( .A(currentPlainKey[38]), .B(n185), .C(n193), .D(n1458), .Y(
        n872) );
  NAND2X1 U1083 ( .A(n183), .B(n1457), .Y(n868) );
  NAND2X1 U1084 ( .A(n1), .B(n1474), .Y(n885) );
  INVX2 U1085 ( .A(n885), .Y(n958) );
  NAND2X1 U1086 ( .A(n958), .B(n1132), .Y(n860) );
  NAND2X1 U1087 ( .A(n49), .B(n153), .Y(n888) );
  INVX2 U1088 ( .A(n888), .Y(n856) );
  NAND2X1 U1089 ( .A(n1852), .B(n856), .Y(n859) );
  AOI21X1 U1093 ( .A(n860), .B(n859), .C(n858), .Y(n863) );
  OAI22X1 U1094 ( .A(n156), .B(n875), .C(n1863), .D(n172), .Y(n861) );
  OAI21X1 U1095 ( .A(n863), .B(n861), .C(n47), .Y(n867) );
  NAND2X1 U1096 ( .A(n897), .B(n203), .Y(n866) );
  NAND3X1 U1097 ( .A(n868), .B(n867), .C(n866), .Y(n870) );
  MUX2X1 U1098 ( .B(n870), .A(n217), .S(n869), .Y(n871) );
  NAND2X1 U1099 ( .A(n872), .B(n871), .Y(n1639) );
  AOI22X1 U1100 ( .A(currentPlainKey[39]), .B(n185), .C(n208), .D(n1458), .Y(
        n884) );
  NAND2X1 U1101 ( .A(n206), .B(n1457), .Y(n880) );
  NOR2X1 U1102 ( .A(n1863), .B(n161), .Y(n874) );
  OAI22X1 U1103 ( .A(n173), .B(n885), .C(n1855), .D(n888), .Y(n873) );
  OAI21X1 U1104 ( .A(n874), .B(n873), .C(n911), .Y(n879) );
  INVX2 U1105 ( .A(n875), .Y(n930) );
  NAND2X1 U1106 ( .A(n930), .B(n181), .Y(n876) );
  NAND3X1 U1107 ( .A(n880), .B(n879), .C(n876), .Y(n881) );
  NAND2X1 U1108 ( .A(n47), .B(n881), .Y(n883) );
  NAND2X1 U1109 ( .A(n897), .B(n195), .Y(n882) );
  NAND3X1 U1110 ( .A(n884), .B(n883), .C(n882), .Y(n1640) );
  AOI22X1 U1114 ( .A(currentPlainKey[40]), .B(n185), .C(n193), .D(n1457), .Y(
        n900) );
  NAND2X1 U1115 ( .A(n183), .B(n1456), .Y(n896) );
  OAI22X1 U1116 ( .A(n156), .B(n885), .C(n1869), .D(n172), .Y(n890) );
  NAND2X1 U1117 ( .A(n1), .B(n7), .Y(n938) );
  NAND2X1 U1118 ( .A(n1869), .B(n938), .Y(n920) );
  INVX2 U1119 ( .A(n920), .Y(n974) );
  NAND2X1 U1120 ( .A(n1859), .B(n974), .Y(n887) );
  OAI22X1 U1121 ( .A(n135), .B(n938), .C(n888), .D(n887), .Y(n889) );
  OAI21X1 U1122 ( .A(n890), .B(n889), .C(n911), .Y(n894) );
  NAND2X1 U1123 ( .A(n930), .B(n203), .Y(n892) );
  NAND3X1 U1124 ( .A(n896), .B(n894), .C(n892), .Y(n898) );
  MUX2X1 U1125 ( .B(n898), .A(n217), .S(n897), .Y(n899) );
  NAND2X1 U1129 ( .A(n900), .B(n899), .Y(n1641) );
  NAND2X1 U1130 ( .A(n930), .B(n195), .Y(n916) );
  NAND2X1 U1131 ( .A(n958), .B(n180), .Y(n909) );
  NOR2X1 U1132 ( .A(n1869), .B(n161), .Y(n904) );
  INVX2 U1133 ( .A(n1862), .Y(n901) );
  NAND3X1 U1134 ( .A(n974), .B(n153), .C(n901), .Y(n902) );
  OAI21X1 U1135 ( .A(n173), .B(n938), .C(n902), .Y(n903) );
  OAI21X1 U1136 ( .A(n904), .B(n903), .C(n49), .Y(n906) );
  NAND2X1 U1137 ( .A(n206), .B(n1456), .Y(n905) );
  NAND3X1 U1138 ( .A(n909), .B(n906), .C(n905), .Y(n910) );
  NAND2X1 U1139 ( .A(n911), .B(n910), .Y(n915) );
  AND2X2 U1140 ( .A(currentPlainKey[41]), .B(n185), .Y(n912) );
  AOI21X1 U1141 ( .A(n210), .B(n1457), .C(n912), .Y(n913) );
  NAND3X1 U1142 ( .A(n916), .B(n915), .C(n913), .Y(n1642) );
  AOI22X1 U1143 ( .A(currentPlainKey[42]), .B(n185), .C(n193), .D(n1456), .Y(
        n933) );
  NAND2X1 U1144 ( .A(n183), .B(n1455), .Y(n929) );
  NAND2X1 U1145 ( .A(n79), .B(n917), .Y(n950) );
  INVX2 U1146 ( .A(n950), .Y(n1021) );
  NAND2X1 U1147 ( .A(n1021), .B(n1132), .Y(n924) );
  NAND2X1 U1148 ( .A(n31), .B(n153), .Y(n952) );
  INVX2 U1149 ( .A(n952), .Y(n918) );
  NAND2X1 U1150 ( .A(n1865), .B(n918), .Y(n923) );
  AOI21X1 U1151 ( .A(n924), .B(n923), .C(n920), .Y(n926) );
  OAI22X1 U1152 ( .A(n156), .B(n938), .C(n1875), .D(n172), .Y(n925) );
  OAI21X1 U1153 ( .A(n926), .B(n925), .C(n49), .Y(n928) );
  NAND2X1 U1158 ( .A(n958), .B(n203), .Y(n927) );
  NAND3X1 U1159 ( .A(n929), .B(n928), .C(n927), .Y(n931) );
  MUX2X1 U1160 ( .B(n931), .A(n210), .S(n930), .Y(n932) );
  NAND2X1 U1161 ( .A(n933), .B(n932), .Y(n1643) );
  AOI22X1 U1162 ( .A(currentPlainKey[43]), .B(n185), .C(n209), .D(n1456), .Y(
        n947) );
  NAND2X1 U1163 ( .A(n206), .B(n1455), .Y(n942) );
  NOR2X1 U1164 ( .A(n1875), .B(n161), .Y(n937) );
  OAI22X1 U1165 ( .A(n173), .B(n950), .C(n1868), .D(n952), .Y(n936) );
  OAI21X1 U1166 ( .A(n937), .B(n936), .C(n974), .Y(n940) );
  INVX2 U1167 ( .A(n938), .Y(n993) );
  NAND2X1 U1168 ( .A(n993), .B(n181), .Y(n939) );
  NAND3X1 U1169 ( .A(n942), .B(n940), .C(n939), .Y(n943) );
  NAND2X1 U1170 ( .A(n49), .B(n943), .Y(n945) );
  NAND2X1 U1171 ( .A(n958), .B(n195), .Y(n944) );
  NAND3X1 U1172 ( .A(n947), .B(n945), .C(n944), .Y(n1644) );
  AOI22X1 U1173 ( .A(currentPlainKey[44]), .B(n185), .C(n193), .D(n1455), .Y(
        n963) );
  NAND2X1 U1174 ( .A(n181), .B(n1454), .Y(n957) );
  OAI22X1 U1175 ( .A(n156), .B(n950), .C(n1881), .D(n168), .Y(n954) );
  NAND2X1 U1176 ( .A(n79), .B(n8), .Y(n999) );
  NAND2X1 U1177 ( .A(n1881), .B(n999), .Y(n982) );
  INVX2 U1178 ( .A(n982), .Y(n1036) );
  NAND2X1 U1179 ( .A(n1871), .B(n1036), .Y(n951) );
  OAI22X1 U1180 ( .A(n135), .B(n999), .C(n952), .D(n951), .Y(n953) );
  OAI21X1 U1181 ( .A(n954), .B(n953), .C(n974), .Y(n956) );
  NAND2X1 U1188 ( .A(n993), .B(n203), .Y(n955) );
  NAND3X1 U1191 ( .A(n957), .B(n956), .C(n955), .Y(n959) );
  MUX2X1 U1192 ( .B(n959), .A(n210), .S(n958), .Y(n960) );
  NAND2X1 U1193 ( .A(n963), .B(n960), .Y(n1645) );
  NAND2X1 U1194 ( .A(n993), .B(n197), .Y(n980) );
  NAND2X1 U1195 ( .A(n1021), .B(n180), .Y(n971) );
  NOR2X1 U1196 ( .A(n1881), .B(n161), .Y(n967) );
  INVX2 U1197 ( .A(n1874), .Y(n964) );
  NAND3X1 U1198 ( .A(n1036), .B(n153), .C(n964), .Y(n965) );
  OAI21X1 U1200 ( .A(n172), .B(n999), .C(n965), .Y(n966) );
  OAI21X1 U1201 ( .A(n967), .B(n966), .C(n31), .Y(n970) );
  NAND2X1 U1202 ( .A(n206), .B(n1454), .Y(n969) );
  NAND3X1 U1203 ( .A(n971), .B(n970), .C(n969), .Y(n972) );
  NAND2X1 U1204 ( .A(n974), .B(n972), .Y(n979) );
  AND2X2 U1205 ( .A(currentPlainKey[45]), .B(n187), .Y(n977) );
  AOI21X1 U1206 ( .A(n209), .B(n1455), .C(n977), .Y(n978) );
  NAND3X1 U1207 ( .A(n980), .B(n979), .C(n978), .Y(n1646) );
  AOI22X1 U1208 ( .A(currentPlainKey[46]), .B(n187), .C(n193), .D(n1454), .Y(
        n996) );
  NAND2X1 U1209 ( .A(n181), .B(n1453), .Y(n992) );
  NAND2X1 U1210 ( .A(n20), .B(n79), .Y(n1010) );
  INVX2 U1211 ( .A(n1010), .Y(n1079) );
  NAND2X1 U1212 ( .A(n1079), .B(n1132), .Y(n984) );
  NAND2X1 U1213 ( .A(n29), .B(n153), .Y(n1013) );
  INVX2 U1214 ( .A(n1013), .Y(n981) );
  NAND2X1 U1215 ( .A(n1877), .B(n981), .Y(n983) );
  AOI21X1 U1216 ( .A(n984), .B(n983), .C(n982), .Y(n986) );
  OAI22X1 U1217 ( .A(n156), .B(n999), .C(n1888), .D(n168), .Y(n985) );
  OAI21X1 U1218 ( .A(n986), .B(n985), .C(n31), .Y(n991) );
  NAND2X1 U1219 ( .A(n1021), .B(n205), .Y(n987) );
  NAND3X1 U1221 ( .A(n992), .B(n991), .C(n987), .Y(n994) );
  MUX2X1 U1222 ( .B(n994), .A(n210), .S(n993), .Y(n995) );
  NAND2X1 U1223 ( .A(n996), .B(n995), .Y(n1647) );
  AOI22X1 U1224 ( .A(currentPlainKey[47]), .B(n187), .C(n208), .D(n1454), .Y(
        n1009) );
  NAND2X1 U1225 ( .A(n206), .B(n1453), .Y(n1003) );
  NOR2X1 U1226 ( .A(n1888), .B(n161), .Y(n998) );
  OAI22X1 U1227 ( .A(n71), .B(n1010), .C(n1880), .D(n1013), .Y(n997) );
  OAI21X1 U1228 ( .A(n998), .B(n997), .C(n1036), .Y(n1001) );
  INVX2 U1229 ( .A(n999), .Y(n1053) );
  NAND2X1 U1230 ( .A(n1053), .B(n180), .Y(n1000) );
  NAND3X1 U1231 ( .A(n1003), .B(n1001), .C(n1000), .Y(n1005) );
  NAND2X1 U1232 ( .A(n31), .B(n1005), .Y(n1008) );
  NAND2X1 U1233 ( .A(n1021), .B(n197), .Y(n1007) );
  NAND3X1 U1234 ( .A(n1009), .B(n1008), .C(n1007), .Y(n1648) );
  AOI22X1 U1235 ( .A(currentPlainKey[48]), .B(n185), .C(n193), .D(n1453), .Y(
        n1024) );
  NAND2X1 U1236 ( .A(n181), .B(n1452), .Y(n1020) );
  OAI22X1 U1237 ( .A(n156), .B(n1010), .C(n1896), .D(n168), .Y(n1015) );
  NAND2X1 U1238 ( .A(n79), .B(n23), .Y(n1059) );
  NAND2X1 U1239 ( .A(n1896), .B(n1059), .Y(n1043) );
  INVX2 U1240 ( .A(n1043), .Y(n1093) );
  NAND2X1 U1241 ( .A(n1883), .B(n1093), .Y(n1012) );
  OAI22X1 U1242 ( .A(n135), .B(n1059), .C(n1013), .D(n1012), .Y(n1014) );
  OAI21X1 U1243 ( .A(n1015), .B(n1014), .C(n1036), .Y(n1017) );
  NAND2X1 U1244 ( .A(n1053), .B(n203), .Y(n1016) );
  NAND3X1 U1245 ( .A(n1020), .B(n1017), .C(n1016), .Y(n1022) );
  MUX2X1 U1246 ( .B(n1022), .A(n210), .S(n1021), .Y(n1023) );
  NAND2X1 U1247 ( .A(n1024), .B(n1023), .Y(n1649) );
  NAND2X1 U1248 ( .A(n1053), .B(n197), .Y(n1041) );
  NAND2X1 U1249 ( .A(n1079), .B(n180), .Y(n1032) );
  NOR2X1 U1250 ( .A(n1896), .B(n161), .Y(n1028) );
  INVX2 U1251 ( .A(n1887), .Y(n1025) );
  NAND3X1 U1252 ( .A(n1093), .B(n153), .C(n1025), .Y(n1026) );
  OAI21X1 U1253 ( .A(n168), .B(n1059), .C(n1026), .Y(n1027) );
  OAI21X1 U1254 ( .A(n1028), .B(n1027), .C(n29), .Y(n1030) );
  NAND2X1 U1255 ( .A(n206), .B(n1452), .Y(n1029) );
  NAND3X1 U1256 ( .A(n1032), .B(n1030), .C(n1029), .Y(n1035) );
  NAND2X1 U1257 ( .A(n1036), .B(n1035), .Y(n1040) );
  AND2X2 U1258 ( .A(currentPlainKey[49]), .B(n187), .Y(n1037) );
  AOI21X1 U1259 ( .A(n209), .B(n1453), .C(n1037), .Y(n1039) );
  NAND3X1 U1260 ( .A(n1041), .B(n1040), .C(n1039), .Y(n1650) );
  AOI22X1 U1261 ( .A(currentPlainKey[50]), .B(n186), .C(n192), .D(n1452), .Y(
        n1056) );
  NAND2X1 U1262 ( .A(n183), .B(n1451), .Y(n1052) );
  NAND2X1 U1263 ( .A(n5), .B(n119), .Y(n1069) );
  INVX2 U1264 ( .A(n1069), .Y(n1140) );
  NAND2X1 U1265 ( .A(n1140), .B(n1132), .Y(n1045) );
  NAND2X1 U1266 ( .A(n51), .B(n153), .Y(n1071) );
  INVX2 U1267 ( .A(n1071), .Y(n1042) );
  NAND2X1 U1268 ( .A(n1891), .B(n1042), .Y(n1044) );
  AOI21X1 U1269 ( .A(n1045), .B(n1044), .C(n1043), .Y(n1049) );
  OAI22X1 U1270 ( .A(n158), .B(n1059), .C(n1903), .D(n168), .Y(n1048) );
  OAI21X1 U1271 ( .A(n1049), .B(n1048), .C(n29), .Y(n1051) );
  NAND2X1 U1272 ( .A(n1079), .B(n203), .Y(n1050) );
  NAND3X1 U1275 ( .A(n1052), .B(n1051), .C(n1050), .Y(n1054) );
  MUX2X1 U1276 ( .B(n1054), .A(n210), .S(n1053), .Y(n1055) );
  NAND2X1 U1277 ( .A(n1056), .B(n1055), .Y(n1651) );
  AOI22X1 U1278 ( .A(currentPlainKey[51]), .B(n187), .C(n208), .D(n1452), .Y(
        n1068) );
  NAND2X1 U1279 ( .A(n207), .B(n1451), .Y(n1064) );
  NOR2X1 U1280 ( .A(n1903), .B(n161), .Y(n1058) );
  OAI22X1 U1281 ( .A(n173), .B(n1069), .C(n1895), .D(n1071), .Y(n1057) );
  OAI21X1 U1282 ( .A(n1058), .B(n1057), .C(n1093), .Y(n1061) );
  INVX2 U1283 ( .A(n1059), .Y(n1114) );
  NAND2X1 U1284 ( .A(n1114), .B(n180), .Y(n1060) );
  NAND3X1 U1285 ( .A(n1064), .B(n1061), .C(n1060), .Y(n1065) );
  NAND2X1 U1286 ( .A(n29), .B(n1065), .Y(n1067) );
  NAND2X1 U1287 ( .A(n1079), .B(n197), .Y(n1066) );
  NAND3X1 U1288 ( .A(n1068), .B(n1067), .C(n1066), .Y(n1652) );
  AOI22X1 U1289 ( .A(currentPlainKey[52]), .B(n187), .C(n192), .D(n1451), .Y(
        n1082) );
  NAND2X1 U1290 ( .A(n181), .B(n1450), .Y(n1076) );
  OAI22X1 U1291 ( .A(n156), .B(n1069), .C(n1910), .D(n168), .Y(n1073) );
  NAND2X1 U1292 ( .A(n5), .B(n1477), .Y(n1118) );
  NAND2X1 U1293 ( .A(n1910), .B(n1118), .Y(n1099) );
  INVX2 U1294 ( .A(n1099), .Y(n1153) );
  NAND2X1 U1295 ( .A(n1898), .B(n1153), .Y(n1070) );
  OAI22X1 U1296 ( .A(n1118), .B(n133), .C(n1071), .D(n1070), .Y(n1072) );
  OAI21X1 U1297 ( .A(n1073), .B(n1072), .C(n1093), .Y(n1075) );
  NAND2X1 U1298 ( .A(n1114), .B(n203), .Y(n1074) );
  NAND3X1 U1299 ( .A(n1076), .B(n1075), .C(n1074), .Y(n1080) );
  MUX2X1 U1300 ( .B(n1080), .A(n210), .S(n1079), .Y(n1081) );
  NAND2X1 U1301 ( .A(n1082), .B(n1081), .Y(n1653) );
  NAND2X1 U1302 ( .A(n1114), .B(n197), .Y(n1097) );
  NAND2X1 U1303 ( .A(n1140), .B(n180), .Y(n1091) );
  NOR2X1 U1304 ( .A(n1910), .B(n161), .Y(n1086) );
  INVX2 U1306 ( .A(n1902), .Y(n1083) );
  NAND3X1 U1307 ( .A(n1153), .B(n153), .C(n1083), .Y(n1084) );
  OAI21X1 U1308 ( .A(n173), .B(n1118), .C(n1084), .Y(n1085) );
  OAI21X1 U1309 ( .A(n1086), .B(n1085), .C(n51), .Y(n1088) );
  NAND2X1 U1310 ( .A(n206), .B(n1450), .Y(n1087) );
  NAND3X1 U1311 ( .A(n1091), .B(n1088), .C(n1087), .Y(n1092) );
  NAND2X1 U1312 ( .A(n1093), .B(n1092), .Y(n1096) );
  AND2X2 U1313 ( .A(currentPlainKey[53]), .B(n187), .Y(n1094) );
  AOI21X1 U1316 ( .A(n209), .B(n1451), .C(n1094), .Y(n1095) );
  NAND3X1 U1317 ( .A(n1097), .B(n1096), .C(n1095), .Y(n1654) );
  AOI22X1 U1318 ( .A(currentPlainKey[54]), .B(n185), .C(n192), .D(n1450), .Y(
        n1117) );
  NAND2X1 U1319 ( .A(n181), .B(n1449), .Y(n1113) );
  NAND2X1 U1320 ( .A(n5), .B(n1474), .Y(n1121) );
  NAND2X1 U1321 ( .A(n1921), .B(n1121), .Y(n1134) );
  INVX2 U1322 ( .A(n1134), .Y(n1174) );
  NAND3X1 U1323 ( .A(n1905), .B(n153), .C(n1174), .Y(n1102) );
  INVX2 U1324 ( .A(n1121), .Y(n1190) );
  NAND2X1 U1325 ( .A(n1132), .B(n1190), .Y(n1100) );
  AOI21X1 U1326 ( .A(n1102), .B(n1100), .C(n1099), .Y(n1110) );
  OAI22X1 U1327 ( .A(n1921), .B(n71), .C(n156), .D(n1118), .Y(n1109) );
  OAI21X1 U1328 ( .A(n1110), .B(n1109), .C(n51), .Y(n1112) );
  NAND2X1 U1329 ( .A(n1140), .B(n203), .Y(n1111) );
  NAND3X1 U1330 ( .A(n1113), .B(n1112), .C(n1111), .Y(n1115) );
  MUX2X1 U1331 ( .B(n1115), .A(n210), .S(n1114), .Y(n1116) );
  NAND2X1 U1332 ( .A(n1117), .B(n1116), .Y(n1655) );
  NAND2X1 U1333 ( .A(n1140), .B(n197), .Y(n1131) );
  INVX2 U1334 ( .A(n1118), .Y(n1165) );
  NAND2X1 U1335 ( .A(n1165), .B(n178), .Y(n1126) );
  NOR2X1 U1336 ( .A(n1921), .B(n161), .Y(n1123) );
  INVX2 U1337 ( .A(n1909), .Y(n1119) );
  NAND3X1 U1338 ( .A(n1174), .B(n11), .C(n1119), .Y(n1120) );
  OAI21X1 U1339 ( .A(n1121), .B(n71), .C(n1120), .Y(n1122) );
  OAI21X1 U1340 ( .A(n1123), .B(n1122), .C(n1153), .Y(n1125) );
  NAND2X1 U1341 ( .A(n207), .B(n1449), .Y(n1124) );
  NAND3X1 U1342 ( .A(n1126), .B(n1125), .C(n1124), .Y(n1127) );
  NAND2X1 U1343 ( .A(n51), .B(n1127), .Y(n1130) );
  AND2X2 U1344 ( .A(currentPlainKey[55]), .B(n187), .Y(n1128) );
  AOI21X1 U1345 ( .A(n209), .B(n1450), .C(n1128), .Y(n1129) );
  NAND3X1 U1346 ( .A(n1131), .B(n1130), .C(n1129), .Y(n1656) );
  AOI22X1 U1347 ( .A(currentPlainKey[56]), .B(n186), .C(n192), .D(n1449), .Y(
        n1145) );
  NAND2X1 U1348 ( .A(n181), .B(n1448), .Y(n1139) );
  NAND2X1 U1349 ( .A(n5), .B(n7), .Y(n1170) );
  NAND3X1 U1350 ( .A(n1098), .B(n1170), .C(n1931), .Y(n1146) );
  INVX2 U1351 ( .A(n1146), .Y(n1196) );
  INVX2 U1352 ( .A(n1170), .Y(n1266) );
  AOI22X1 U1353 ( .A(n1915), .B(n1196), .C(n1132), .D(n1266), .Y(n1135) );
  AOI22X1 U1354 ( .A(n166), .B(n1190), .C(n175), .D(n1447), .Y(n1133) );
  OAI21X1 U1355 ( .A(n1135), .B(n1134), .C(n1133), .Y(n1136) );
  NAND2X1 U1356 ( .A(n1153), .B(n1136), .Y(n1138) );
  NAND2X1 U1357 ( .A(n1165), .B(n203), .Y(n1137) );
  NAND3X1 U1358 ( .A(n1139), .B(n1138), .C(n1137), .Y(n1141) );
  MUX2X1 U1359 ( .B(n1141), .A(n210), .S(n1140), .Y(n1142) );
  NAND2X1 U1360 ( .A(n1145), .B(n1142), .Y(n1657) );
  AOI22X1 U1361 ( .A(currentPlainKey[57]), .B(n187), .C(n208), .D(n1449), .Y(
        n1156) );
  NAND2X1 U1362 ( .A(n207), .B(n1448), .Y(n1151) );
  NOR2X1 U1363 ( .A(n1920), .B(n1146), .Y(n1148) );
  OAI22X1 U1364 ( .A(n1931), .B(n156), .C(n1170), .D(n168), .Y(n1147) );
  OAI21X1 U1365 ( .A(n1148), .B(n1147), .C(n1174), .Y(n1150) );
  NAND2X1 U1366 ( .A(n1190), .B(n178), .Y(n1149) );
  NAND3X1 U1367 ( .A(n1151), .B(n1150), .C(n1149), .Y(n1152) );
  NAND2X1 U1368 ( .A(n1153), .B(n1152), .Y(n1155) );
  NAND2X1 U1369 ( .A(n1165), .B(n197), .Y(n1154) );
  NAND3X1 U1370 ( .A(n1156), .B(n1155), .C(n1154), .Y(n1658) );
  AOI22X1 U1371 ( .A(currentPlainKey[58]), .B(n187), .C(n192), .D(n1448), .Y(
        n1168) );
  NAND2X1 U1372 ( .A(n181), .B(n1447), .Y(n1164) );
  NAND2X1 U1373 ( .A(n1196), .B(n1969), .Y(n1183) );
  INVX2 U1374 ( .A(n1925), .Y(n1157) );
  NOR2X1 U1375 ( .A(n1183), .B(n1157), .Y(n1161) );
  OAI22X1 U1376 ( .A(n1969), .B(n71), .C(n1170), .D(n156), .Y(n1159) );
  OAI21X1 U1377 ( .A(n1161), .B(n1159), .C(n1174), .Y(n1163) );
  NAND2X1 U1378 ( .A(n1190), .B(n203), .Y(n1162) );
  NAND3X1 U1379 ( .A(n1164), .B(n1163), .C(n1162), .Y(n1166) );
  MUX2X1 U1380 ( .B(n1166), .A(n210), .S(n1165), .Y(n1167) );
  NAND2X1 U1381 ( .A(n1168), .B(n1167), .Y(n1659) );
  AOI22X1 U1382 ( .A(currentPlainKey[59]), .B(n187), .C(n208), .D(n1448), .Y(
        n1180) );
  OAI22X1 U1383 ( .A(n1931), .B(n1171), .C(n1170), .D(n1169), .Y(n1176) );
  INVX2 U1384 ( .A(n1930), .Y(n1173) );
  NAND3X1 U1385 ( .A(RCV_DATA[3]), .B(n1446), .C(n1196), .Y(n1172) );
  OAI21X1 U1386 ( .A(n1183), .B(n1173), .C(n1172), .Y(n1175) );
  OAI21X1 U1387 ( .A(n1176), .B(n1175), .C(n1174), .Y(n1179) );
  NAND2X1 U1388 ( .A(n1190), .B(n197), .Y(n1177) );
  NAND3X1 U1389 ( .A(n1180), .B(n1179), .C(n1177), .Y(n1660) );
  AOI22X1 U1390 ( .A(currentPlainKey[60]), .B(n185), .C(n192), .D(n1447), .Y(
        n1193) );
  NAND2X1 U1391 ( .A(n183), .B(n1446), .Y(n1189) );
  AOI22X1 U1392 ( .A(n1493), .B(RCV_DATA[3]), .C(n1445), .D(RCV_DATA[2]), .Y(
        n1182) );
  OAI21X1 U1393 ( .A(n222), .B(n1963), .C(n1182), .Y(n1185) );
  INVX2 U1394 ( .A(n1183), .Y(n1184) );
  OAI21X1 U1395 ( .A(n55), .B(n1185), .C(n1184), .Y(n1188) );
  NAND2X1 U1396 ( .A(n207), .B(n1266), .Y(n1187) );
  NAND3X1 U1397 ( .A(n1189), .B(n1188), .C(n1187), .Y(n1191) );
  MUX2X1 U1398 ( .B(n1191), .A(n210), .S(n1190), .Y(n1192) );
  NAND2X1 U1399 ( .A(n1193), .B(n1192), .Y(n1661) );
  AOI22X1 U1400 ( .A(currentPlainKey[61]), .B(n187), .C(n208), .D(n1447), .Y(
        n1263) );
  NAND2X1 U1401 ( .A(n1446), .B(RCV_DATA[5]), .Y(n1194) );
  NAND2X1 U1402 ( .A(n1944), .B(n1194), .Y(n1195) );
  NAND2X1 U1403 ( .A(n1196), .B(n1195), .Y(n1262) );
  NAND2X1 U1404 ( .A(n1266), .B(n197), .Y(n1261) );
  NAND3X1 U1405 ( .A(n1263), .B(n1262), .C(n1261), .Y(n1662) );
  AND2X2 U1406 ( .A(n187), .B(currentPlainKey[62]), .Y(n1264) );
  AOI21X1 U1407 ( .A(n195), .B(n1446), .C(n1264), .Y(n1359) );
  NOR2X1 U1408 ( .A(n1446), .B(n99), .Y(n1265) );
  OAI21X1 U1409 ( .A(n1954), .B(n1953), .C(n1265), .Y(n1268) );
  MUX2X1 U1410 ( .B(n1268), .A(n1267), .S(n1266), .Y(n1357) );
  INVX2 U1411 ( .A(n1357), .Y(n1358) );
  NAND2X1 U1412 ( .A(n1359), .B(n1358), .Y(n1663) );
  NAND2X1 U1413 ( .A(n186), .B(currentPlainKey[63]), .Y(n1370) );
  NAND2X1 U1414 ( .A(n197), .B(n1493), .Y(n1366) );
  NOR2X1 U1415 ( .A(n1445), .B(n99), .Y(n1363) );
  INVX2 U1416 ( .A(n1968), .Y(n1362) );
  OAI21X1 U1417 ( .A(n203), .B(n1363), .C(n1362), .Y(n1365) );
  NAND2X1 U1418 ( .A(n1366), .B(n1365), .Y(n1368) );
  MUX2X1 U1419 ( .B(n1368), .A(n217), .S(n1446), .Y(n1369) );
  NAND2X1 U1420 ( .A(n1370), .B(n1369), .Y(n1664) );
  NAND2X1 U1421 ( .A(n1371), .B(n1414), .Y(n1382) );
  INVX2 U1422 ( .A(n1382), .Y(n1372) );
  NAND3X1 U1423 ( .A(n1372), .B(n233), .C(n1426), .Y(n1380) );
  INVX2 U1424 ( .A(n1380), .Y(n1378) );
  NAND2X1 U1425 ( .A(n1378), .B(keyCount[3]), .Y(n1381) );
  NAND2X1 U1426 ( .A(address[0]), .B(n1380), .Y(n1373) );
  NAND2X1 U1427 ( .A(n1381), .B(n1373), .Y(n1600) );
  NAND2X1 U1428 ( .A(address[1]), .B(n1380), .Y(n1374) );
  NAND2X1 U1429 ( .A(n1381), .B(n1374), .Y(n1599) );
  NAND2X1 U1430 ( .A(address[2]), .B(n1380), .Y(n1375) );
  NAND2X1 U1431 ( .A(n1381), .B(n1375), .Y(n1598) );
  MUX2X1 U1432 ( .B(address[3]), .A(keyCount[0]), .S(n1378), .Y(n1376) );
  NAND2X1 U1433 ( .A(n1381), .B(n1376), .Y(n1597) );
  MUX2X1 U1434 ( .B(address[4]), .A(keyCount[1]), .S(n1378), .Y(n1377) );
  NAND2X1 U1435 ( .A(n1381), .B(n1377), .Y(n1596) );
  MUX2X1 U1436 ( .B(address[5]), .A(keyCount[2]), .S(n1378), .Y(n1379) );
  NAND2X1 U1437 ( .A(n1381), .B(n1379), .Y(n1595) );
  OAI21X1 U1438 ( .A(n1499), .B(n1378), .C(n1381), .Y(n1594) );
  OAI21X1 U1439 ( .A(n1491), .B(n1378), .C(n1381), .Y(n1593) );
  OAI21X1 U1440 ( .A(n1383), .B(n1382), .C(parityError), .Y(n1386) );
  OAI21X1 U1441 ( .A(n2037), .B(n2036), .C(n1384), .Y(n1385) );
  NAND2X1 U1442 ( .A(n1386), .B(n1385), .Y(nextParityError) );
  NOR2X1 U1443 ( .A(keyCount[0]), .B(n1438), .Y(n1387) );
  NOR2X1 U1444 ( .A(n1387), .B(n1442), .Y(n1390) );
  INVX2 U1445 ( .A(n1444), .Y(n1388) );
  NAND2X1 U1446 ( .A(keyCount[0]), .B(n1388), .Y(n1389) );
  MUX2X1 U1447 ( .B(n1390), .A(n1389), .S(n1490), .Y(n1583) );
  NAND2X1 U1448 ( .A(n1391), .B(CLR_RBUFF), .Y(n1405) );
  INVX2 U1449 ( .A(n1405), .Y(n1400) );
  NAND2X1 U1450 ( .A(N1799), .B(n1400), .Y(n1392) );
  OAI21X1 U1451 ( .A(n1489), .B(n1393), .C(n1392), .Y(n1592) );
  NAND2X1 U1452 ( .A(N1798), .B(n1400), .Y(n1394) );
  OAI21X1 U1453 ( .A(n1488), .B(n1395), .C(n1394), .Y(n1591) );
  NAND2X1 U1454 ( .A(N1797), .B(n1400), .Y(n1396) );
  OAI21X1 U1455 ( .A(n1487), .B(n1395), .C(n1396), .Y(n1590) );
  NAND2X1 U1456 ( .A(N1796), .B(n1400), .Y(n1397) );
  OAI21X1 U1457 ( .A(n1486), .B(n1393), .C(n1397), .Y(n1589) );
  NAND2X1 U1458 ( .A(N1795), .B(n1400), .Y(n1398) );
  OAI21X1 U1459 ( .A(n1485), .B(n1399), .C(n1398), .Y(n1588) );
  NAND2X1 U1460 ( .A(N1794), .B(n1400), .Y(n1401) );
  OAI21X1 U1461 ( .A(n1484), .B(n1399), .C(n1401), .Y(n1587) );
  INVX2 U1462 ( .A(N1793), .Y(n1402) );
  OAI22X1 U1463 ( .A(n1483), .B(n1393), .C(n1405), .D(n1402), .Y(n1586) );
  INVX2 U1464 ( .A(N1792), .Y(n1404) );
  OAI22X1 U1465 ( .A(n1482), .B(n1395), .C(n1405), .D(n1404), .Y(n1585) );
  AOI21X1 U1466 ( .A(N694), .B(RBUF_FULL), .C(n1730), .Y(n1407) );
  NAND2X1 U1467 ( .A(n1407), .B(n1406), .Y(n1410) );
  NAND2X1 U1468 ( .A(n1408), .B(n115), .Y(n1409) );
  NAND2X1 U1469 ( .A(n1409), .B(n1424), .Y(n1431) );
  NAND2X1 U1470 ( .A(n1410), .B(n1431), .Y(n1421) );
  INVX2 U1471 ( .A(n1421), .Y(n1412) );
  OAI21X1 U1472 ( .A(n1412), .B(n115), .C(n1411), .Y(n1579) );
  AND2X2 U1473 ( .A(n1425), .B(n1426), .Y(n1418) );
  OAI21X1 U1474 ( .A(OE), .B(SBE), .C(n1406), .Y(n1417) );
  OAI22X1 U1475 ( .A(RBUF_FULL), .B(n1414), .C(n1413), .D(n1431), .Y(n1415) );
  AOI21X1 U1476 ( .A(n1420), .B(n1433), .C(n1415), .Y(n1416) );
  NAND3X1 U1477 ( .A(n1418), .B(n1417), .C(n1416), .Y(n1581) );
  AOI21X1 U1478 ( .A(state[1]), .B(n1421), .C(n1420), .Y(n1422) );
  NAND2X1 U1479 ( .A(n113), .B(n1422), .Y(n1582) );
  INVX2 U1480 ( .A(RBUF_FULL), .Y(n1423) );
  AOI21X1 U1481 ( .A(n1425), .B(n1424), .C(n1423), .Y(n1430) );
  NAND2X1 U1482 ( .A(n1570), .B(n1576), .Y(n1428) );
  OAI21X1 U1483 ( .A(n1428), .B(n1427), .C(n1426), .Y(n1429) );
  NOR2X1 U1484 ( .A(n1430), .B(n1429), .Y(n1437) );
  INVX2 U1485 ( .A(n1731), .Y(n1433) );
  OAI22X1 U1486 ( .A(n1438), .B(n1433), .C(n1432), .D(n1431), .Y(n1434) );
  NOR2X1 U1487 ( .A(n1435), .B(n1434), .Y(n1436) );
  NAND2X1 U1488 ( .A(n1437), .B(n1436), .Y(n1580) );
  NOR2X1 U1489 ( .A(keyCount[2]), .B(n1438), .Y(n1440) );
  OAI21X1 U1490 ( .A(n1440), .B(n1439), .C(keyCount[3]), .Y(n1441) );
  OAI21X1 U1491 ( .A(n1731), .B(n1444), .C(n1441), .Y(n1578) );
  NAND2X1 U1492 ( .A(n1442), .B(keyCount[0]), .Y(n1443) );
  OAI21X1 U1493 ( .A(keyCount[0]), .B(n1444), .C(n1443), .Y(n1577) );
  INVX2 U1494 ( .A(keyCount[3]), .Y(N694) );
  INVX2 U1495 ( .A(keyCount[0]), .Y(n1479) );
  INVX2 U1496 ( .A(keyCount[2]), .Y(n1480) );
  INVX2 U1497 ( .A(parityAccumulator[0]), .Y(n1482) );
  INVX2 U1498 ( .A(parityAccumulator[1]), .Y(n1483) );
  INVX2 U1499 ( .A(parityAccumulator[2]), .Y(n1484) );
  INVX2 U1500 ( .A(parityAccumulator[3]), .Y(n1485) );
  INVX2 U1501 ( .A(parityAccumulator[4]), .Y(n1486) );
  INVX2 U1502 ( .A(parityAccumulator[5]), .Y(n1487) );
  INVX2 U1503 ( .A(parityAccumulator[6]), .Y(n1488) );
  INVX2 U1504 ( .A(parityAccumulator[7]), .Y(n1489) );
  INVX2 U1505 ( .A(keyCount[1]), .Y(n1490) );
  INVX2 U1506 ( .A(address[7]), .Y(n1491) );
  INVX2 U1507 ( .A(n1945), .Y(n1492) );
  INVX2 U1508 ( .A(n1967), .Y(n1493) );
  INVX2 U1509 ( .A(n1963), .Y(n1494) );
  INVX2 U1510 ( .A(n1962), .Y(n1495) );
  INVX2 U1511 ( .A(n1959), .Y(n1496) );
  INVX2 U1512 ( .A(n1957), .Y(n1497) );
  INVX2 U1513 ( .A(address[6]), .Y(n1499) );
  INVX2 U1514 ( .A(n1923), .Y(n1500) );
  INVX2 U1515 ( .A(n1927), .Y(n1501) );
  INVX2 U1516 ( .A(n1938), .Y(n1502) );
  INVX2 U1517 ( .A(n1956), .Y(n1503) );
  INVX2 U1518 ( .A(address[5]), .Y(n1504) );
  INVX2 U1519 ( .A(address[4]), .Y(n1505) );
  INVX2 U1520 ( .A(currentPlainKey[63]), .Y(n1506) );
  INVX2 U1521 ( .A(currentPlainKey[62]), .Y(n1507) );
  INVX2 U1522 ( .A(currentPlainKey[61]), .Y(n1508) );
  INVX2 U1523 ( .A(currentPlainKey[60]), .Y(n1509) );
  INVX2 U1524 ( .A(currentPlainKey[59]), .Y(n1510) );
  INVX2 U1525 ( .A(currentPlainKey[58]), .Y(n1511) );
  INVX2 U1526 ( .A(currentPlainKey[57]), .Y(n1512) );
  INVX2 U1527 ( .A(currentPlainKey[56]), .Y(n1513) );
  INVX2 U1528 ( .A(currentPlainKey[55]), .Y(n1514) );
  INVX2 U1529 ( .A(currentPlainKey[54]), .Y(n1515) );
  INVX2 U1530 ( .A(currentPlainKey[53]), .Y(n1516) );
  INVX2 U1531 ( .A(currentPlainKey[52]), .Y(n1517) );
  INVX2 U1532 ( .A(currentPlainKey[51]), .Y(n1518) );
  INVX2 U1533 ( .A(currentPlainKey[50]), .Y(n1519) );
  INVX2 U1534 ( .A(currentPlainKey[49]), .Y(n1520) );
  INVX2 U1535 ( .A(currentPlainKey[48]), .Y(n1521) );
  INVX2 U1536 ( .A(currentPlainKey[47]), .Y(n1522) );
  INVX2 U1537 ( .A(currentPlainKey[46]), .Y(n1523) );
  INVX2 U1538 ( .A(currentPlainKey[45]), .Y(n1524) );
  INVX2 U1539 ( .A(currentPlainKey[44]), .Y(n1525) );
  INVX2 U1540 ( .A(currentPlainKey[43]), .Y(n1526) );
  INVX2 U1541 ( .A(currentPlainKey[42]), .Y(n1527) );
  INVX2 U1542 ( .A(currentPlainKey[41]), .Y(n1528) );
  INVX2 U1543 ( .A(currentPlainKey[40]), .Y(n1529) );
  INVX2 U1544 ( .A(currentPlainKey[39]), .Y(n1530) );
  INVX2 U1545 ( .A(currentPlainKey[38]), .Y(n1531) );
  INVX2 U1546 ( .A(currentPlainKey[37]), .Y(n1532) );
  INVX2 U1547 ( .A(currentPlainKey[36]), .Y(n1533) );
  INVX2 U1548 ( .A(currentPlainKey[35]), .Y(n1534) );
  INVX2 U1549 ( .A(currentPlainKey[34]), .Y(n1535) );
  INVX2 U1550 ( .A(currentPlainKey[33]), .Y(n1536) );
  INVX2 U1551 ( .A(currentPlainKey[32]), .Y(n1537) );
  INVX2 U1552 ( .A(currentPlainKey[31]), .Y(n1538) );
  INVX2 U1553 ( .A(currentPlainKey[30]), .Y(n1539) );
  INVX2 U1554 ( .A(currentPlainKey[29]), .Y(n1540) );
  INVX2 U1555 ( .A(currentPlainKey[28]), .Y(n1541) );
  INVX2 U1556 ( .A(currentPlainKey[27]), .Y(n1542) );
  INVX2 U1557 ( .A(currentPlainKey[26]), .Y(n1543) );
  INVX2 U1558 ( .A(currentPlainKey[25]), .Y(n1544) );
  INVX2 U1559 ( .A(currentPlainKey[24]), .Y(n1545) );
  INVX2 U1560 ( .A(currentPlainKey[23]), .Y(n1546) );
  INVX2 U1561 ( .A(currentPlainKey[22]), .Y(n1547) );
  INVX2 U1562 ( .A(currentPlainKey[21]), .Y(n1548) );
  INVX2 U1563 ( .A(currentPlainKey[20]), .Y(n1549) );
  INVX2 U1564 ( .A(currentPlainKey[19]), .Y(n1550) );
  INVX2 U1565 ( .A(currentPlainKey[18]), .Y(n1551) );
  INVX2 U1566 ( .A(currentPlainKey[17]), .Y(n1552) );
  INVX2 U1567 ( .A(currentPlainKey[16]), .Y(n1553) );
  INVX2 U1568 ( .A(currentPlainKey[15]), .Y(n1554) );
  INVX2 U1569 ( .A(currentPlainKey[14]), .Y(n1555) );
  INVX2 U1570 ( .A(currentPlainKey[13]), .Y(n1556) );
  INVX2 U1571 ( .A(currentPlainKey[12]), .Y(n1557) );
  INVX2 U1572 ( .A(currentPlainKey[11]), .Y(n1558) );
  INVX2 U1573 ( .A(currentPlainKey[10]), .Y(n1559) );
  INVX2 U1574 ( .A(currentPlainKey[9]), .Y(n1560) );
  INVX2 U1575 ( .A(currentPlainKey[8]), .Y(n1561) );
  INVX2 U1576 ( .A(currentPlainKey[7]), .Y(n1562) );
  INVX2 U1577 ( .A(currentPlainKey[6]), .Y(n1563) );
  INVX2 U1578 ( .A(currentPlainKey[5]), .Y(n1564) );
  INVX2 U1579 ( .A(currentPlainKey[4]), .Y(n1565) );
  INVX2 U1580 ( .A(currentPlainKey[0]), .Y(n1569) );
  INVX2 U1581 ( .A(SBE), .Y(n1570) );
  INVX2 U1582 ( .A(OE), .Y(n1576) );
endmodule


module uart_timer_0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module uart_timer_0 ( CLK, RST, TIMER_TRIG, STOP_RCVING, SHIFT_STROBE );
  input CLK, RST, TIMER_TRIG;
  output STOP_RCVING, SHIFT_STROBE;
  wire   N26, N27, N28, N29, N30, N31, N32, N33, N60, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110;
  wire   [7:0] state;
  wire   [7:0] nextState;
  assign SHIFT_STROBE = N60;

  OR2X2 U21 ( .A(state[7]), .B(n95), .Y(n96) );
  OAI21X1 U38 ( .A(n20), .B(n27), .C(n110), .Y(n81) );
  NAND2X1 U39 ( .A(N33), .B(n109), .Y(n110) );
  OAI21X1 U40 ( .A(n26), .B(n20), .C(n108), .Y(n80) );
  NAND2X1 U41 ( .A(N32), .B(n109), .Y(n108) );
  OAI21X1 U42 ( .A(n25), .B(n20), .C(n107), .Y(n79) );
  NAND2X1 U43 ( .A(N31), .B(n109), .Y(n107) );
  OAI21X1 U44 ( .A(n20), .B(n24), .C(n106), .Y(n78) );
  NAND2X1 U45 ( .A(N30), .B(n109), .Y(n106) );
  OAI21X1 U46 ( .A(n23), .B(n20), .C(n105), .Y(n77) );
  NAND2X1 U47 ( .A(N29), .B(n109), .Y(n105) );
  OAI21X1 U48 ( .A(n22), .B(n20), .C(n104), .Y(n76) );
  NAND2X1 U49 ( .A(N28), .B(n109), .Y(n104) );
  OAI21X1 U50 ( .A(n20), .B(n21), .C(n103), .Y(n75) );
  NAND2X1 U51 ( .A(N27), .B(n109), .Y(n103) );
  OAI21X1 U52 ( .A(n19), .B(n20), .C(n102), .Y(n74) );
  NAND2X1 U53 ( .A(N26), .B(n109), .Y(n102) );
  NOR2X1 U54 ( .A(n101), .B(n73), .Y(n109) );
  NOR2X1 U55 ( .A(n73), .B(TIMER_TRIG), .Y(n101) );
  NOR2X1 U56 ( .A(n100), .B(n99), .Y(n73) );
  NAND3X1 U57 ( .A(nextState[6]), .B(nextState[5]), .C(n98), .Y(n99) );
  NOR2X1 U58 ( .A(n22), .B(n23), .Y(n98) );
  NAND3X1 U59 ( .A(nextState[0]), .B(n21), .C(n97), .Y(n100) );
  NOR2X1 U60 ( .A(nextState[7]), .B(nextState[4]), .Y(n97) );
  NOR2X1 U61 ( .A(state[0]), .B(n96), .Y(N60) );
  AOI21X1 U62 ( .A(n94), .B(n32), .C(n93), .Y(n95) );
  OAI21X1 U63 ( .A(n33), .B(n92), .C(n91), .Y(n93) );
  NAND3X1 U64 ( .A(state[6]), .B(state[1]), .C(n90), .Y(n91) );
  AOI21X1 U65 ( .A(n89), .B(n88), .C(state[3]), .Y(n90) );
  NAND3X1 U66 ( .A(n33), .B(n31), .C(state[4]), .Y(n88) );
  NAND3X1 U67 ( .A(state[2]), .B(n32), .C(state[5]), .Y(n89) );
  NAND2X1 U68 ( .A(state[4]), .B(n87), .Y(n92) );
  OAI21X1 U69 ( .A(state[2]), .B(n28), .C(n86), .Y(n94) );
  NAND3X1 U70 ( .A(state[2]), .B(n29), .C(n30), .Y(n86) );
  OAI22X1 U71 ( .A(state[6]), .B(n84), .C(n29), .D(n85), .Y(n87) );
  NAND3X1 U72 ( .A(n34), .B(n31), .C(state[3]), .Y(n85) );
  AOI22X1 U73 ( .A(n83), .B(state[1]), .C(n82), .D(state[5]), .Y(n84) );
  XOR2X1 U74 ( .A(n34), .B(state[3]), .Y(n82) );
  NOR2X1 U75 ( .A(state[5]), .B(state[3]), .Y(n83) );
  uart_timer_0_DW01_inc_0 add_39 ( .A(nextState), .SUM({N33, N32, N31, N30, 
        N29, N28, N27, N26}) );
  DFFSR \state_reg[3]  ( .D(nextState[3]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[3]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[5]  ( .D(nextState[5]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[5]) );
  DFFSR \state_reg[6]  ( .D(nextState[6]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[6]) );
  DFFSR \state_reg[4]  ( .D(nextState[4]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[4]) );
  DFFSR \state_reg[7]  ( .D(nextState[7]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[7]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        state[0]) );
  DFFSR STOP_RCVING_reg ( .D(n73), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        STOP_RCVING) );
  DFFSR \nextState_reg[3]  ( .D(n77), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[3]) );
  DFFSR \nextState_reg[2]  ( .D(n76), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[2]) );
  DFFSR \nextState_reg[0]  ( .D(n74), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[0]) );
  DFFSR \nextState_reg[4]  ( .D(n78), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[4]) );
  DFFSR \nextState_reg[1]  ( .D(n75), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[1]) );
  DFFSR \nextState_reg[5]  ( .D(n79), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[5]) );
  DFFSR \nextState_reg[6]  ( .D(n80), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[6]) );
  DFFSR \nextState_reg[7]  ( .D(n81), .CLK(CLK), .R(n18), .S(1'b1), .Q(
        nextState[7]) );
  INVX2 U20 ( .A(RST), .Y(n18) );
  INVX2 U22 ( .A(nextState[0]), .Y(n19) );
  INVX2 U23 ( .A(n101), .Y(n20) );
  INVX2 U24 ( .A(nextState[1]), .Y(n21) );
  INVX2 U25 ( .A(nextState[2]), .Y(n22) );
  INVX2 U26 ( .A(nextState[3]), .Y(n23) );
  INVX2 U27 ( .A(nextState[4]), .Y(n24) );
  INVX2 U28 ( .A(nextState[5]), .Y(n25) );
  INVX2 U29 ( .A(nextState[6]), .Y(n26) );
  INVX2 U30 ( .A(nextState[7]), .Y(n27) );
  INVX2 U31 ( .A(n87), .Y(n28) );
  INVX2 U32 ( .A(state[6]), .Y(n29) );
  INVX2 U33 ( .A(n85), .Y(n30) );
  INVX2 U34 ( .A(state[5]), .Y(n31) );
  INVX2 U35 ( .A(state[4]), .Y(n32) );
  INVX2 U36 ( .A(state[2]), .Y(n33) );
  INVX2 U37 ( .A(state[1]), .Y(n34) );
endmodule


module uart_rcv_block_0 ( CLK, RST, SERIAL_IN, KEY_ERROR, PROG_ERROR, PLAINKEY, 
        RBUF_FULL, PARITY_ERROR );
  output [63:0] PLAINKEY;
  input CLK, RST, SERIAL_IN;
  output KEY_ERROR, PROG_ERROR, RBUF_FULL, PARITY_ERROR;
  wire   START_BIT, CHK_ERROR, OE, SB_DETECT, STOP_RCVING, RBUF_LOAD, SBC_CLR,
         SBC_EN, SET_RBUF_FULL, TIMER_TRIG, CLR_RBUF, SBE, SHIFT_STROBE, n1,
         n2;
  wire   [7:0] LOAD_DATA;
  wire   [7:0] RCV_DATA;
  wire   [1:0] STOP_DATA;

  uart_edge_detector_0 U_0 ( .CLK(CLK), .RST(n1), .SERIAL_IN(SERIAL_IN), 
        .START_BIT(START_BIT) );
  uart_error_0 U_1 ( .RST(n1), .CLK(CLK), .RBUF_FULL(RBUF_FULL), .CHK_ERROR(
        CHK_ERROR), .OE(OE) );
  uart_rcu_0 U_2 ( .CLK(CLK), .RST(n1), .START_BIT(START_BIT), .STOP_RCVING(
        STOP_RCVING), .SB_DETECT(SB_DETECT), .RBUF_LOAD(RBUF_LOAD), 
        .TIMER_TRIG(TIMER_TRIG), .CHK_ERROR(CHK_ERROR), .SET_RBUF_FULL(
        SET_RBUF_FULL), .SBC_EN(SBC_EN), .SBC_CLR(SBC_CLR) );
  uart_rcv_buf_0 U_3 ( .CLK(CLK), .RST(n1), .LOAD_RBUF(RBUF_LOAD), .LOAD_DATA(
        LOAD_DATA), .RCV_DATA(RCV_DATA) );
  uart_rcv_buf_full_0 U_4 ( .CLK(CLK), .RST(n1), .CLR_RBUF(CLR_RBUF), 
        .SET_RBUF_FULL(SET_RBUF_FULL), .RBUF_FULL(RBUF_FULL) );
  uart_sb_check_0 U_5 ( .RST(n1), .CLK(CLK), .SBC_CLR(SBC_CLR), .SBC_EN(SBC_EN), .STOP_DATA(STOP_DATA), .SB_DETECT(SB_DETECT), .SBE(SBE) );
  uart_sr_10bit_0 U_6 ( .CLK(CLK), .RST(n1), .SHIFT_STROBE(SHIFT_STROBE), 
        .SERIAL_IN(SERIAL_IN), .LOAD_DATA(LOAD_DATA), .STOP_DATA(STOP_DATA) );
  keyreg_0 U_8 ( .CLK(CLK), .RST(n1), .SBE(SBE), .OE(OE), .RBUF_FULL(RBUF_FULL), .RCV_DATA(RCV_DATA), .PLAINKEY(PLAINKEY), .KEY_ERROR(KEY_ERROR), 
        .PROG_ERROR(PROG_ERROR), .CLR_RBUFF(CLR_RBUF), .PARITY_ERROR(
        PARITY_ERROR) );
  uart_timer_0 U_7 ( .CLK(CLK), .RST(n1), .TIMER_TRIG(TIMER_TRIG), 
        .STOP_RCVING(STOP_RCVING), .SHIFT_STROBE(SHIFT_STROBE) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module EDBlock_0 ( BYTE, BYTE_READY, CLK, OPCODE, RST, SERIAL_IN, DATA_IN, 
        KEY_ERROR, PARITY_ERROR, PDATA_READY, PROCESSED_DATA, PROG_ERROR, 
        RBUF_FULL, W_ENABLE, R_ENABLE, DATA, ADDR );
  input [7:0] BYTE;
  input [1:0] OPCODE;
  input [7:0] DATA_IN;
  output [7:0] PROCESSED_DATA;
  output [7:0] DATA;
  output [7:0] ADDR;
  input BYTE_READY, CLK, RST, SERIAL_IN;
  output KEY_ERROR, PARITY_ERROR, PDATA_READY, PROG_ERROR, RBUF_FULL, W_ENABLE,
         R_ENABLE;
  wire   n1, n2;
  wire   [63:0] PLAINKEY;

  KSA_0 U_0 ( .KEY(PLAINKEY), .CLK(CLK), .RST(n1), .KEY_ERROR(KEY_ERROR), 
        .BYTE_READY(BYTE_READY), .BYTE(BYTE), .OPCODE(OPCODE), .DATA_IN(
        DATA_IN), .PROCESSED_DATA(PROCESSED_DATA), .PDATA_READY(PDATA_READY), 
        .W_ENABLE(W_ENABLE), .R_ENABLE(R_ENABLE), .ADDR(ADDR), .DATA(DATA) );
  uart_rcv_block_0 U_1 ( .CLK(CLK), .RST(n1), .SERIAL_IN(SERIAL_IN), 
        .KEY_ERROR(KEY_ERROR), .PROG_ERROR(PROG_ERROR), .PLAINKEY(PLAINKEY), 
        .RBUF_FULL(RBUF_FULL), .PARITY_ERROR(PARITY_ERROR) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module RBUFFER_0 ( CLK, RST, NEXT_BYTE, DATA, OPCODE, BYTE_COUNT, EOP, B_READY, 
        R_ENABLE, PRGA_IN, PRGA_OPCODE );
  input [7:0] DATA;
  input [1:0] OPCODE;
  input [4:0] BYTE_COUNT;
  output [7:0] PRGA_IN;
  output [1:0] PRGA_OPCODE;
  input CLK, RST, NEXT_BYTE, EOP;
  output B_READY, R_ENABLE;
  wire   N39, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103;
  wire   [2:0] state;
  wire   [2:0] nextState;
  wire   [7:0] tempData;
  wire   [1:0] tempOpcode;
  assign N39 = BYTE_COUNT[4];

  DFFPOSX1 B_READY_reg ( .D(n92), .CLK(CLK), .Q(B_READY) );
  DFFPOSX1 \tempData_reg[7]  ( .D(n71), .CLK(CLK), .Q(tempData[7]) );
  DFFPOSX1 \tempData_reg[6]  ( .D(n72), .CLK(CLK), .Q(tempData[6]) );
  DFFPOSX1 \tempData_reg[5]  ( .D(n73), .CLK(CLK), .Q(tempData[5]) );
  DFFPOSX1 \tempData_reg[4]  ( .D(n74), .CLK(CLK), .Q(tempData[4]) );
  DFFPOSX1 \tempData_reg[3]  ( .D(n75), .CLK(CLK), .Q(tempData[3]) );
  DFFPOSX1 \tempData_reg[2]  ( .D(n86), .CLK(CLK), .Q(tempData[2]) );
  DFFPOSX1 \tempData_reg[1]  ( .D(n88), .CLK(CLK), .Q(tempData[1]) );
  DFFPOSX1 \tempData_reg[0]  ( .D(n89), .CLK(CLK), .Q(tempData[0]) );
  DFFPOSX1 \tempOpcode_reg[1]  ( .D(n90), .CLK(CLK), .Q(tempOpcode[1]) );
  DFFPOSX1 \PRGA_OPCODE_reg[1]  ( .D(n93), .CLK(CLK), .Q(PRGA_OPCODE[1]) );
  DFFPOSX1 \tempOpcode_reg[0]  ( .D(n91), .CLK(CLK), .Q(tempOpcode[0]) );
  DFFPOSX1 \PRGA_OPCODE_reg[0]  ( .D(n94), .CLK(CLK), .Q(PRGA_OPCODE[0]) );
  DFFPOSX1 R_ENABLE_reg ( .D(n95), .CLK(CLK), .Q(R_ENABLE) );
  DFFPOSX1 \PRGA_IN_reg[7]  ( .D(n96), .CLK(CLK), .Q(PRGA_IN[7]) );
  DFFPOSX1 \PRGA_IN_reg[6]  ( .D(n97), .CLK(CLK), .Q(PRGA_IN[6]) );
  DFFPOSX1 \PRGA_IN_reg[5]  ( .D(n98), .CLK(CLK), .Q(PRGA_IN[5]) );
  DFFPOSX1 \PRGA_IN_reg[4]  ( .D(n99), .CLK(CLK), .Q(PRGA_IN[4]) );
  DFFPOSX1 \PRGA_IN_reg[3]  ( .D(n100), .CLK(CLK), .Q(PRGA_IN[3]) );
  DFFPOSX1 \PRGA_IN_reg[2]  ( .D(n101), .CLK(CLK), .Q(PRGA_IN[2]) );
  DFFPOSX1 \PRGA_IN_reg[1]  ( .D(n102), .CLK(CLK), .Q(PRGA_IN[1]) );
  DFFPOSX1 \PRGA_IN_reg[0]  ( .D(n103), .CLK(CLK), .Q(PRGA_IN[0]) );
  DFFSR \state_reg[1]  ( .D(nextState[1]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[2]  ( .D(nextState[2]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[0]  ( .D(nextState[0]), .CLK(CLK), .R(n4), .S(1'b1), .Q(
        state[0]) );
  INVX2 U6 ( .A(n44), .Y(n31) );
  INVX2 U7 ( .A(RST), .Y(n4) );
  OR2X2 U8 ( .A(n42), .B(RST), .Y(n32) );
  AND2X2 U9 ( .A(n42), .B(n4), .Y(n47) );
  OAI21X1 U10 ( .A(n5), .B(n6), .C(n7), .Y(nextState[2]) );
  MUX2X1 U11 ( .B(n8), .A(n9), .S(state[0]), .Y(n7) );
  NOR2X1 U12 ( .A(state[2]), .B(n10), .Y(n9) );
  AND2X1 U13 ( .A(state[2]), .B(n11), .Y(n8) );
  OAI21X1 U14 ( .A(NEXT_BYTE), .B(n12), .C(state[1]), .Y(n11) );
  AND2X1 U15 ( .A(n13), .B(NEXT_BYTE), .Y(n5) );
  OAI21X1 U16 ( .A(state[2]), .B(n14), .C(n15), .Y(nextState[1]) );
  OAI21X1 U17 ( .A(n16), .B(n17), .C(n18), .Y(n15) );
  INVX1 U18 ( .A(n6), .Y(n17) );
  OAI21X1 U19 ( .A(state[2]), .B(n19), .C(n20), .Y(nextState[0]) );
  AOI22X1 U20 ( .A(n21), .B(n22), .C(NEXT_BYTE), .D(n23), .Y(n20) );
  OAI21X1 U21 ( .A(n13), .B(n6), .C(n24), .Y(n23) );
  INVX1 U22 ( .A(n16), .Y(n24) );
  NOR2X1 U23 ( .A(n19), .B(n12), .Y(n16) );
  NOR2X1 U24 ( .A(n25), .B(N39), .Y(n12) );
  NAND3X1 U25 ( .A(state[0]), .B(n10), .C(state[2]), .Y(n6) );
  AND2X1 U26 ( .A(OPCODE[1]), .B(OPCODE[0]), .Y(n13) );
  OAI21X1 U27 ( .A(n26), .B(n18), .C(n27), .Y(n22) );
  INVX1 U28 ( .A(NEXT_BYTE), .Y(n18) );
  AOI21X1 U29 ( .A(EOP), .B(n25), .C(N39), .Y(n26) );
  NAND2X1 U30 ( .A(n28), .B(n29), .Y(n25) );
  NOR2X1 U31 ( .A(BYTE_COUNT[3]), .B(BYTE_COUNT[2]), .Y(n29) );
  NOR2X1 U32 ( .A(BYTE_COUNT[1]), .B(BYTE_COUNT[0]), .Y(n28) );
  NOR2X1 U33 ( .A(state[1]), .B(state[0]), .Y(n21) );
  INVX1 U34 ( .A(n30), .Y(n71) );
  AOI22X1 U35 ( .A(n31), .B(DATA[7]), .C(n32), .D(tempData[7]), .Y(n30) );
  INVX1 U36 ( .A(n33), .Y(n72) );
  AOI22X1 U37 ( .A(n31), .B(DATA[6]), .C(n32), .D(tempData[6]), .Y(n33) );
  INVX1 U38 ( .A(n34), .Y(n73) );
  AOI22X1 U39 ( .A(n31), .B(DATA[5]), .C(n32), .D(tempData[5]), .Y(n34) );
  INVX1 U40 ( .A(n35), .Y(n74) );
  AOI22X1 U41 ( .A(n31), .B(DATA[4]), .C(n32), .D(tempData[4]), .Y(n35) );
  INVX1 U42 ( .A(n36), .Y(n75) );
  AOI22X1 U43 ( .A(n31), .B(DATA[3]), .C(n32), .D(tempData[3]), .Y(n36) );
  INVX1 U44 ( .A(n37), .Y(n86) );
  AOI22X1 U45 ( .A(n31), .B(DATA[2]), .C(n32), .D(tempData[2]), .Y(n37) );
  INVX1 U46 ( .A(n38), .Y(n88) );
  AOI22X1 U47 ( .A(n31), .B(DATA[1]), .C(n32), .D(tempData[1]), .Y(n38) );
  INVX1 U48 ( .A(n39), .Y(n89) );
  AOI22X1 U49 ( .A(n31), .B(DATA[0]), .C(n32), .D(tempData[0]), .Y(n39) );
  INVX1 U50 ( .A(n40), .Y(n90) );
  AOI22X1 U51 ( .A(OPCODE[1]), .B(n31), .C(n32), .D(tempOpcode[1]), .Y(n40) );
  INVX1 U52 ( .A(n41), .Y(n91) );
  AOI22X1 U53 ( .A(OPCODE[0]), .B(n31), .C(n32), .D(tempOpcode[0]), .Y(n41) );
  OAI21X1 U54 ( .A(n4), .B(n43), .C(n44), .Y(n92) );
  INVX1 U55 ( .A(B_READY), .Y(n43) );
  OAI21X1 U56 ( .A(n4), .B(n45), .C(n46), .Y(n93) );
  AOI22X1 U57 ( .A(n31), .B(OPCODE[1]), .C(n47), .D(tempOpcode[1]), .Y(n46) );
  INVX1 U58 ( .A(PRGA_OPCODE[1]), .Y(n45) );
  OAI21X1 U59 ( .A(n4), .B(n48), .C(n49), .Y(n94) );
  AOI22X1 U60 ( .A(n31), .B(OPCODE[0]), .C(n47), .D(tempOpcode[0]), .Y(n49) );
  INVX1 U61 ( .A(PRGA_OPCODE[0]), .Y(n48) );
  MUX2X1 U62 ( .B(n50), .A(n51), .S(RST), .Y(n95) );
  INVX1 U63 ( .A(R_ENABLE), .Y(n51) );
  NAND3X1 U64 ( .A(n10), .B(n27), .C(state[0]), .Y(n50) );
  OAI21X1 U65 ( .A(n4), .B(n52), .C(n53), .Y(n96) );
  AOI22X1 U66 ( .A(DATA[7]), .B(n31), .C(n47), .D(tempData[7]), .Y(n53) );
  INVX1 U67 ( .A(PRGA_IN[7]), .Y(n52) );
  OAI21X1 U68 ( .A(n4), .B(n54), .C(n55), .Y(n97) );
  AOI22X1 U69 ( .A(DATA[6]), .B(n31), .C(n47), .D(tempData[6]), .Y(n55) );
  INVX1 U70 ( .A(PRGA_IN[6]), .Y(n54) );
  OAI21X1 U71 ( .A(n4), .B(n56), .C(n57), .Y(n98) );
  AOI22X1 U72 ( .A(DATA[5]), .B(n31), .C(n47), .D(tempData[5]), .Y(n57) );
  INVX1 U73 ( .A(PRGA_IN[5]), .Y(n56) );
  OAI21X1 U74 ( .A(n4), .B(n58), .C(n59), .Y(n99) );
  AOI22X1 U75 ( .A(DATA[4]), .B(n31), .C(n47), .D(tempData[4]), .Y(n59) );
  INVX1 U76 ( .A(PRGA_IN[4]), .Y(n58) );
  OAI21X1 U77 ( .A(n4), .B(n60), .C(n61), .Y(n100) );
  AOI22X1 U78 ( .A(DATA[3]), .B(n31), .C(n47), .D(tempData[3]), .Y(n61) );
  INVX1 U79 ( .A(PRGA_IN[3]), .Y(n60) );
  OAI21X1 U80 ( .A(n4), .B(n62), .C(n63), .Y(n101) );
  AOI22X1 U81 ( .A(DATA[2]), .B(n31), .C(n47), .D(tempData[2]), .Y(n63) );
  INVX1 U82 ( .A(PRGA_IN[2]), .Y(n62) );
  OAI21X1 U83 ( .A(n4), .B(n64), .C(n65), .Y(n102) );
  AOI22X1 U84 ( .A(DATA[1]), .B(n31), .C(n47), .D(tempData[1]), .Y(n65) );
  INVX1 U85 ( .A(PRGA_IN[1]), .Y(n64) );
  OAI21X1 U86 ( .A(n4), .B(n66), .C(n67), .Y(n103) );
  AOI22X1 U87 ( .A(DATA[0]), .B(n31), .C(n47), .D(tempData[0]), .Y(n67) );
  NAND2X1 U88 ( .A(n14), .B(state[2]), .Y(n42) );
  INVX1 U89 ( .A(n68), .Y(n14) );
  OAI21X1 U90 ( .A(state[1]), .B(n69), .C(n19), .Y(n68) );
  NAND2X1 U91 ( .A(state[1]), .B(n69), .Y(n19) );
  NAND3X1 U92 ( .A(n69), .B(n10), .C(n70), .Y(n44) );
  NOR2X1 U93 ( .A(RST), .B(n27), .Y(n70) );
  INVX1 U94 ( .A(state[2]), .Y(n27) );
  INVX1 U95 ( .A(state[1]), .Y(n10) );
  INVX1 U96 ( .A(state[0]), .Y(n69) );
  INVX1 U97 ( .A(PRGA_IN[0]), .Y(n66) );
endmodule


module RFIFO_0 ( CLK, RST, W_ENABLE, R_ENABLE, RCV_DATA, RCV_OPCODE, DATA, 
        OUT_OPCODE, BYTE_COUNT, EMPTY, FULL );
  input [7:0] RCV_DATA;
  input [1:0] RCV_OPCODE;
  output [7:0] DATA;
  output [1:0] OUT_OPCODE;
  output [4:0] BYTE_COUNT;
  input CLK, RST, W_ENABLE, R_ENABLE;
  output EMPTY, FULL;
  wire   state, N32, N33, N34, N43, N44, N45, N46, \opcode[0][1] ,
         \opcode[0][0] , \opcode[1][1] , \opcode[1][0] , \opcode[2][1] ,
         \opcode[2][0] , \opcode[3][1] , \opcode[3][0] , \opcode[4][1] ,
         \opcode[4][0] , \opcode[5][1] , \opcode[5][0] , \opcode[6][1] ,
         \opcode[6][0] , \opcode[7][1] , \opcode[7][0] , \opcode[8][1] ,
         \opcode[8][0] , \opcode[9][1] , \opcode[9][0] , \opcode[10][1] ,
         \opcode[10][0] , \opcode[11][1] , \opcode[11][0] , \opcode[12][1] ,
         \opcode[12][0] , \opcode[13][1] , \opcode[13][0] , \opcode[14][1] ,
         \opcode[14][0] , \opcode[15][1] , \opcode[15][0] , \opcode[16][1] ,
         \opcode[16][0] , \opcode[17][1] , \opcode[17][0] , \opcode[18][1] ,
         \opcode[18][0] , \opcode[19][1] , \opcode[19][0] , \opcode[20][1] ,
         \opcode[20][0] , \opcode[21][1] , \opcode[21][0] , \opcode[22][1] ,
         \opcode[22][0] , \opcode[23][1] , \opcode[23][0] , \opcode[24][1] ,
         \opcode[24][0] , \opcode[25][1] , \opcode[25][0] , \opcode[26][1] ,
         \opcode[26][0] , \opcode[27][1] , \opcode[27][0] , \opcode[28][1] ,
         \opcode[28][0] , \opcode[29][1] , \opcode[29][0] , \opcode[30][1] ,
         \opcode[30][0] , \opcode[31][1] , \opcode[31][0] , \memory[0][7] ,
         \memory[0][6] , \memory[0][5] , \memory[0][4] , \memory[0][3] ,
         \memory[0][2] , \memory[0][1] , \memory[0][0] , \memory[1][7] ,
         \memory[1][6] , \memory[1][5] , \memory[1][4] , \memory[1][3] ,
         \memory[1][2] , \memory[1][1] , \memory[1][0] , \memory[2][7] ,
         \memory[2][6] , \memory[2][5] , \memory[2][4] , \memory[2][3] ,
         \memory[2][2] , \memory[2][1] , \memory[2][0] , \memory[3][7] ,
         \memory[3][6] , \memory[3][5] , \memory[3][4] , \memory[3][3] ,
         \memory[3][2] , \memory[3][1] , \memory[3][0] , \memory[4][7] ,
         \memory[4][6] , \memory[4][5] , \memory[4][4] , \memory[4][3] ,
         \memory[4][2] , \memory[4][1] , \memory[4][0] , \memory[5][7] ,
         \memory[5][6] , \memory[5][5] , \memory[5][4] , \memory[5][3] ,
         \memory[5][2] , \memory[5][1] , \memory[5][0] , \memory[6][7] ,
         \memory[6][6] , \memory[6][5] , \memory[6][4] , \memory[6][3] ,
         \memory[6][2] , \memory[6][1] , \memory[6][0] , \memory[7][7] ,
         \memory[7][6] , \memory[7][5] , \memory[7][4] , \memory[7][3] ,
         \memory[7][2] , \memory[7][1] , \memory[7][0] , \memory[8][7] ,
         \memory[8][6] , \memory[8][5] , \memory[8][4] , \memory[8][3] ,
         \memory[8][2] , \memory[8][1] , \memory[8][0] , \memory[9][7] ,
         \memory[9][6] , \memory[9][5] , \memory[9][4] , \memory[9][3] ,
         \memory[9][2] , \memory[9][1] , \memory[9][0] , \memory[10][7] ,
         \memory[10][6] , \memory[10][5] , \memory[10][4] , \memory[10][3] ,
         \memory[10][2] , \memory[10][1] , \memory[10][0] , \memory[11][7] ,
         \memory[11][6] , \memory[11][5] , \memory[11][4] , \memory[11][3] ,
         \memory[11][2] , \memory[11][1] , \memory[11][0] , \memory[12][7] ,
         \memory[12][6] , \memory[12][5] , \memory[12][4] , \memory[12][3] ,
         \memory[12][2] , \memory[12][1] , \memory[12][0] , \memory[13][7] ,
         \memory[13][6] , \memory[13][5] , \memory[13][4] , \memory[13][3] ,
         \memory[13][2] , \memory[13][1] , \memory[13][0] , \memory[14][7] ,
         \memory[14][6] , \memory[14][5] , \memory[14][4] , \memory[14][3] ,
         \memory[14][2] , \memory[14][1] , \memory[14][0] , \memory[15][7] ,
         \memory[15][6] , \memory[15][5] , \memory[15][4] , \memory[15][3] ,
         \memory[15][2] , \memory[15][1] , \memory[15][0] , \memory[16][7] ,
         \memory[16][6] , \memory[16][5] , \memory[16][4] , \memory[16][3] ,
         \memory[16][2] , \memory[16][1] , \memory[16][0] , \memory[17][7] ,
         \memory[17][6] , \memory[17][5] , \memory[17][4] , \memory[17][3] ,
         \memory[17][2] , \memory[17][1] , \memory[17][0] , \memory[18][7] ,
         \memory[18][6] , \memory[18][5] , \memory[18][4] , \memory[18][3] ,
         \memory[18][2] , \memory[18][1] , \memory[18][0] , \memory[19][7] ,
         \memory[19][6] , \memory[19][5] , \memory[19][4] , \memory[19][3] ,
         \memory[19][2] , \memory[19][1] , \memory[19][0] , \memory[20][7] ,
         \memory[20][6] , \memory[20][5] , \memory[20][4] , \memory[20][3] ,
         \memory[20][2] , \memory[20][1] , \memory[20][0] , \memory[21][7] ,
         \memory[21][6] , \memory[21][5] , \memory[21][4] , \memory[21][3] ,
         \memory[21][2] , \memory[21][1] , \memory[21][0] , \memory[22][7] ,
         \memory[22][6] , \memory[22][5] , \memory[22][4] , \memory[22][3] ,
         \memory[22][2] , \memory[22][1] , \memory[22][0] , \memory[23][7] ,
         \memory[23][6] , \memory[23][5] , \memory[23][4] , \memory[23][3] ,
         \memory[23][2] , \memory[23][1] , \memory[23][0] , \memory[24][7] ,
         \memory[24][6] , \memory[24][5] , \memory[24][4] , \memory[24][3] ,
         \memory[24][2] , \memory[24][1] , \memory[24][0] , \memory[25][7] ,
         \memory[25][6] , \memory[25][5] , \memory[25][4] , \memory[25][3] ,
         \memory[25][2] , \memory[25][1] , \memory[25][0] , \memory[26][7] ,
         \memory[26][6] , \memory[26][5] , \memory[26][4] , \memory[26][3] ,
         \memory[26][2] , \memory[26][1] , \memory[26][0] , \memory[27][7] ,
         \memory[27][6] , \memory[27][5] , \memory[27][4] , \memory[27][3] ,
         \memory[27][2] , \memory[27][1] , \memory[27][0] , \memory[28][7] ,
         \memory[28][6] , \memory[28][5] , \memory[28][4] , \memory[28][3] ,
         \memory[28][2] , \memory[28][1] , \memory[28][0] , \memory[29][7] ,
         \memory[29][6] , \memory[29][5] , \memory[29][4] , \memory[29][3] ,
         \memory[29][2] , \memory[29][1] , \memory[29][0] , \memory[30][7] ,
         \memory[30][6] , \memory[30][5] , \memory[30][4] , \memory[30][3] ,
         \memory[30][2] , \memory[30][1] , \memory[30][0] , \memory[31][7] ,
         \memory[31][6] , \memory[31][5] , \memory[31][4] , \memory[31][3] ,
         \memory[31][2] , \memory[31][1] , \memory[31][0] , N48, N49, N50, N51,
         N189, N190, N191, N192, N193, N195, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         \add_76_aco/carry[4] , \add_76_aco/carry[3] , \add_76_aco/carry[2] ,
         \add_76_aco/carry[1] , \sub_72/carry[4] , \sub_72/carry[3] ,
         \sub_72/carry[2] , \sub_72/carry[1] , \add_67/carry[4] ,
         \add_67/carry[3] , \add_67/carry[2] , \r83/carry[4] , \r83/carry[3] ,
         \r83/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n855, n857, n859, n861, n863,
         n864, n865, n866, n867, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1373, n1374,
         n1375, n1376, n1377;
  wire   [4:0] readptr;
  wire   [4:0] writeptr;

  DFFSR state_reg ( .D(1'b1), .CLK(CLK), .R(n98), .S(1'b1), .Q(state) );
  DFFPOSX1 FULL_reg ( .D(n1200), .CLK(CLK), .Q(FULL) );
  DFFPOSX1 \memory_reg[0][7]  ( .D(n1175), .CLK(CLK), .Q(\memory[0][7] ) );
  DFFPOSX1 \memory_reg[0][6]  ( .D(n1174), .CLK(CLK), .Q(\memory[0][6] ) );
  DFFPOSX1 \memory_reg[0][5]  ( .D(n1173), .CLK(CLK), .Q(\memory[0][5] ) );
  DFFPOSX1 \memory_reg[0][4]  ( .D(n1172), .CLK(CLK), .Q(\memory[0][4] ) );
  DFFPOSX1 \memory_reg[0][3]  ( .D(n1171), .CLK(CLK), .Q(\memory[0][3] ) );
  DFFPOSX1 \memory_reg[0][2]  ( .D(n1170), .CLK(CLK), .Q(\memory[0][2] ) );
  DFFPOSX1 \memory_reg[0][1]  ( .D(n1169), .CLK(CLK), .Q(\memory[0][1] ) );
  DFFPOSX1 \memory_reg[0][0]  ( .D(n1168), .CLK(CLK), .Q(\memory[0][0] ) );
  DFFPOSX1 \memory_reg[1][7]  ( .D(n1183), .CLK(CLK), .Q(\memory[1][7] ) );
  DFFPOSX1 \memory_reg[1][6]  ( .D(n1182), .CLK(CLK), .Q(\memory[1][6] ) );
  DFFPOSX1 \memory_reg[1][5]  ( .D(n1181), .CLK(CLK), .Q(\memory[1][5] ) );
  DFFPOSX1 \memory_reg[1][4]  ( .D(n1180), .CLK(CLK), .Q(\memory[1][4] ) );
  DFFPOSX1 \memory_reg[1][3]  ( .D(n1179), .CLK(CLK), .Q(\memory[1][3] ) );
  DFFPOSX1 \memory_reg[1][2]  ( .D(n1178), .CLK(CLK), .Q(\memory[1][2] ) );
  DFFPOSX1 \memory_reg[1][1]  ( .D(n1177), .CLK(CLK), .Q(\memory[1][1] ) );
  DFFPOSX1 \memory_reg[1][0]  ( .D(n1176), .CLK(CLK), .Q(\memory[1][0] ) );
  DFFPOSX1 \memory_reg[2][7]  ( .D(n1191), .CLK(CLK), .Q(\memory[2][7] ) );
  DFFPOSX1 \memory_reg[2][6]  ( .D(n1190), .CLK(CLK), .Q(\memory[2][6] ) );
  DFFPOSX1 \memory_reg[2][5]  ( .D(n1189), .CLK(CLK), .Q(\memory[2][5] ) );
  DFFPOSX1 \memory_reg[2][4]  ( .D(n1188), .CLK(CLK), .Q(\memory[2][4] ) );
  DFFPOSX1 \memory_reg[2][3]  ( .D(n1187), .CLK(CLK), .Q(\memory[2][3] ) );
  DFFPOSX1 \memory_reg[2][2]  ( .D(n1186), .CLK(CLK), .Q(\memory[2][2] ) );
  DFFPOSX1 \memory_reg[2][1]  ( .D(n1185), .CLK(CLK), .Q(\memory[2][1] ) );
  DFFPOSX1 \memory_reg[2][0]  ( .D(n1184), .CLK(CLK), .Q(\memory[2][0] ) );
  DFFPOSX1 \memory_reg[3][7]  ( .D(n1199), .CLK(CLK), .Q(\memory[3][7] ) );
  DFFPOSX1 \memory_reg[3][6]  ( .D(n1198), .CLK(CLK), .Q(\memory[3][6] ) );
  DFFPOSX1 \memory_reg[3][5]  ( .D(n1197), .CLK(CLK), .Q(\memory[3][5] ) );
  DFFPOSX1 \memory_reg[3][4]  ( .D(n1196), .CLK(CLK), .Q(\memory[3][4] ) );
  DFFPOSX1 \memory_reg[3][3]  ( .D(n1195), .CLK(CLK), .Q(\memory[3][3] ) );
  DFFPOSX1 \memory_reg[3][2]  ( .D(n1194), .CLK(CLK), .Q(\memory[3][2] ) );
  DFFPOSX1 \memory_reg[3][1]  ( .D(n1193), .CLK(CLK), .Q(\memory[3][1] ) );
  DFFPOSX1 \memory_reg[3][0]  ( .D(n1192), .CLK(CLK), .Q(\memory[3][0] ) );
  DFFPOSX1 \memory_reg[4][7]  ( .D(n1371), .CLK(CLK), .Q(\memory[4][7] ) );
  DFFPOSX1 \memory_reg[4][6]  ( .D(n1370), .CLK(CLK), .Q(\memory[4][6] ) );
  DFFPOSX1 \memory_reg[4][5]  ( .D(n1369), .CLK(CLK), .Q(\memory[4][5] ) );
  DFFPOSX1 \memory_reg[4][4]  ( .D(n1368), .CLK(CLK), .Q(\memory[4][4] ) );
  DFFPOSX1 \memory_reg[4][3]  ( .D(n1367), .CLK(CLK), .Q(\memory[4][3] ) );
  DFFPOSX1 \memory_reg[4][2]  ( .D(n1366), .CLK(CLK), .Q(\memory[4][2] ) );
  DFFPOSX1 \memory_reg[4][1]  ( .D(n1365), .CLK(CLK), .Q(\memory[4][1] ) );
  DFFPOSX1 \memory_reg[4][0]  ( .D(n1364), .CLK(CLK), .Q(\memory[4][0] ) );
  DFFPOSX1 \memory_reg[5][7]  ( .D(n1361), .CLK(CLK), .Q(\memory[5][7] ) );
  DFFPOSX1 \memory_reg[5][6]  ( .D(n1360), .CLK(CLK), .Q(\memory[5][6] ) );
  DFFPOSX1 \memory_reg[5][5]  ( .D(n1359), .CLK(CLK), .Q(\memory[5][5] ) );
  DFFPOSX1 \memory_reg[5][4]  ( .D(n1358), .CLK(CLK), .Q(\memory[5][4] ) );
  DFFPOSX1 \memory_reg[5][3]  ( .D(n1357), .CLK(CLK), .Q(\memory[5][3] ) );
  DFFPOSX1 \memory_reg[5][2]  ( .D(n1356), .CLK(CLK), .Q(\memory[5][2] ) );
  DFFPOSX1 \memory_reg[5][1]  ( .D(n1355), .CLK(CLK), .Q(\memory[5][1] ) );
  DFFPOSX1 \memory_reg[5][0]  ( .D(n1354), .CLK(CLK), .Q(\memory[5][0] ) );
  DFFPOSX1 \memory_reg[6][7]  ( .D(n1351), .CLK(CLK), .Q(\memory[6][7] ) );
  DFFPOSX1 \memory_reg[6][6]  ( .D(n1350), .CLK(CLK), .Q(\memory[6][6] ) );
  DFFPOSX1 \memory_reg[6][5]  ( .D(n1349), .CLK(CLK), .Q(\memory[6][5] ) );
  DFFPOSX1 \memory_reg[6][4]  ( .D(n1348), .CLK(CLK), .Q(\memory[6][4] ) );
  DFFPOSX1 \memory_reg[6][3]  ( .D(n1347), .CLK(CLK), .Q(\memory[6][3] ) );
  DFFPOSX1 \memory_reg[6][2]  ( .D(n1346), .CLK(CLK), .Q(\memory[6][2] ) );
  DFFPOSX1 \memory_reg[6][1]  ( .D(n1345), .CLK(CLK), .Q(\memory[6][1] ) );
  DFFPOSX1 \memory_reg[6][0]  ( .D(n1344), .CLK(CLK), .Q(\memory[6][0] ) );
  DFFPOSX1 \memory_reg[7][7]  ( .D(n1341), .CLK(CLK), .Q(\memory[7][7] ) );
  DFFPOSX1 \memory_reg[7][6]  ( .D(n1340), .CLK(CLK), .Q(\memory[7][6] ) );
  DFFPOSX1 \memory_reg[7][5]  ( .D(n1339), .CLK(CLK), .Q(\memory[7][5] ) );
  DFFPOSX1 \memory_reg[7][4]  ( .D(n1338), .CLK(CLK), .Q(\memory[7][4] ) );
  DFFPOSX1 \memory_reg[7][3]  ( .D(n1337), .CLK(CLK), .Q(\memory[7][3] ) );
  DFFPOSX1 \memory_reg[7][2]  ( .D(n1336), .CLK(CLK), .Q(\memory[7][2] ) );
  DFFPOSX1 \memory_reg[7][1]  ( .D(n1335), .CLK(CLK), .Q(\memory[7][1] ) );
  DFFPOSX1 \memory_reg[7][0]  ( .D(n1334), .CLK(CLK), .Q(\memory[7][0] ) );
  DFFPOSX1 \memory_reg[8][7]  ( .D(n1202), .CLK(CLK), .Q(\memory[8][7] ) );
  DFFPOSX1 \memory_reg[8][6]  ( .D(n1203), .CLK(CLK), .Q(\memory[8][6] ) );
  DFFPOSX1 \memory_reg[8][5]  ( .D(n1204), .CLK(CLK), .Q(\memory[8][5] ) );
  DFFPOSX1 \memory_reg[8][4]  ( .D(n1205), .CLK(CLK), .Q(\memory[8][4] ) );
  DFFPOSX1 \memory_reg[8][3]  ( .D(n1206), .CLK(CLK), .Q(\memory[8][3] ) );
  DFFPOSX1 \memory_reg[8][2]  ( .D(n1207), .CLK(CLK), .Q(\memory[8][2] ) );
  DFFPOSX1 \memory_reg[8][1]  ( .D(n1208), .CLK(CLK), .Q(\memory[8][1] ) );
  DFFPOSX1 \memory_reg[8][0]  ( .D(n1209), .CLK(CLK), .Q(\memory[8][0] ) );
  DFFPOSX1 \memory_reg[9][7]  ( .D(n1210), .CLK(CLK), .Q(\memory[9][7] ) );
  DFFPOSX1 \memory_reg[9][6]  ( .D(n1211), .CLK(CLK), .Q(\memory[9][6] ) );
  DFFPOSX1 \memory_reg[9][5]  ( .D(n1212), .CLK(CLK), .Q(\memory[9][5] ) );
  DFFPOSX1 \memory_reg[9][4]  ( .D(n1213), .CLK(CLK), .Q(\memory[9][4] ) );
  DFFPOSX1 \memory_reg[9][3]  ( .D(n1214), .CLK(CLK), .Q(\memory[9][3] ) );
  DFFPOSX1 \memory_reg[9][2]  ( .D(n1215), .CLK(CLK), .Q(\memory[9][2] ) );
  DFFPOSX1 \memory_reg[9][1]  ( .D(n1216), .CLK(CLK), .Q(\memory[9][1] ) );
  DFFPOSX1 \memory_reg[9][0]  ( .D(n1217), .CLK(CLK), .Q(\memory[9][0] ) );
  DFFPOSX1 \memory_reg[10][7]  ( .D(n1218), .CLK(CLK), .Q(\memory[10][7] ) );
  DFFPOSX1 \memory_reg[10][6]  ( .D(n1219), .CLK(CLK), .Q(\memory[10][6] ) );
  DFFPOSX1 \memory_reg[10][5]  ( .D(n1220), .CLK(CLK), .Q(\memory[10][5] ) );
  DFFPOSX1 \memory_reg[10][4]  ( .D(n1221), .CLK(CLK), .Q(\memory[10][4] ) );
  DFFPOSX1 \memory_reg[10][3]  ( .D(n1222), .CLK(CLK), .Q(\memory[10][3] ) );
  DFFPOSX1 \memory_reg[10][2]  ( .D(n1223), .CLK(CLK), .Q(\memory[10][2] ) );
  DFFPOSX1 \memory_reg[10][1]  ( .D(n1224), .CLK(CLK), .Q(\memory[10][1] ) );
  DFFPOSX1 \memory_reg[10][0]  ( .D(n1225), .CLK(CLK), .Q(\memory[10][0] ) );
  DFFPOSX1 \memory_reg[11][7]  ( .D(n1226), .CLK(CLK), .Q(\memory[11][7] ) );
  DFFPOSX1 \memory_reg[11][6]  ( .D(n1227), .CLK(CLK), .Q(\memory[11][6] ) );
  DFFPOSX1 \memory_reg[11][5]  ( .D(n1228), .CLK(CLK), .Q(\memory[11][5] ) );
  DFFPOSX1 \memory_reg[11][4]  ( .D(n1229), .CLK(CLK), .Q(\memory[11][4] ) );
  DFFPOSX1 \memory_reg[11][3]  ( .D(n1230), .CLK(CLK), .Q(\memory[11][3] ) );
  DFFPOSX1 \memory_reg[11][2]  ( .D(n1231), .CLK(CLK), .Q(\memory[11][2] ) );
  DFFPOSX1 \memory_reg[11][1]  ( .D(n1232), .CLK(CLK), .Q(\memory[11][1] ) );
  DFFPOSX1 \memory_reg[11][0]  ( .D(n1233), .CLK(CLK), .Q(\memory[11][0] ) );
  DFFPOSX1 \memory_reg[12][7]  ( .D(n1064), .CLK(CLK), .Q(\memory[12][7] ) );
  DFFPOSX1 \memory_reg[12][6]  ( .D(n1065), .CLK(CLK), .Q(\memory[12][6] ) );
  DFFPOSX1 \memory_reg[12][5]  ( .D(n1066), .CLK(CLK), .Q(\memory[12][5] ) );
  DFFPOSX1 \memory_reg[12][4]  ( .D(n1067), .CLK(CLK), .Q(\memory[12][4] ) );
  DFFPOSX1 \memory_reg[12][3]  ( .D(n1068), .CLK(CLK), .Q(\memory[12][3] ) );
  DFFPOSX1 \memory_reg[12][2]  ( .D(n1069), .CLK(CLK), .Q(\memory[12][2] ) );
  DFFPOSX1 \memory_reg[12][1]  ( .D(n1070), .CLK(CLK), .Q(\memory[12][1] ) );
  DFFPOSX1 \memory_reg[12][0]  ( .D(n1071), .CLK(CLK), .Q(\memory[12][0] ) );
  DFFPOSX1 \memory_reg[13][7]  ( .D(n1022), .CLK(CLK), .Q(\memory[13][7] ) );
  DFFPOSX1 \memory_reg[13][6]  ( .D(n1023), .CLK(CLK), .Q(\memory[13][6] ) );
  DFFPOSX1 \memory_reg[13][5]  ( .D(n1024), .CLK(CLK), .Q(\memory[13][5] ) );
  DFFPOSX1 \memory_reg[13][4]  ( .D(n1025), .CLK(CLK), .Q(\memory[13][4] ) );
  DFFPOSX1 \memory_reg[13][3]  ( .D(n1026), .CLK(CLK), .Q(\memory[13][3] ) );
  DFFPOSX1 \memory_reg[13][2]  ( .D(n1027), .CLK(CLK), .Q(\memory[13][2] ) );
  DFFPOSX1 \memory_reg[13][1]  ( .D(n1028), .CLK(CLK), .Q(\memory[13][1] ) );
  DFFPOSX1 \memory_reg[13][0]  ( .D(n1029), .CLK(CLK), .Q(\memory[13][0] ) );
  DFFPOSX1 \memory_reg[14][7]  ( .D(n1014), .CLK(CLK), .Q(\memory[14][7] ) );
  DFFPOSX1 \memory_reg[14][6]  ( .D(n1015), .CLK(CLK), .Q(\memory[14][6] ) );
  DFFPOSX1 \memory_reg[14][5]  ( .D(n1016), .CLK(CLK), .Q(\memory[14][5] ) );
  DFFPOSX1 \memory_reg[14][4]  ( .D(n1017), .CLK(CLK), .Q(\memory[14][4] ) );
  DFFPOSX1 \memory_reg[14][3]  ( .D(n1018), .CLK(CLK), .Q(\memory[14][3] ) );
  DFFPOSX1 \memory_reg[14][2]  ( .D(n1019), .CLK(CLK), .Q(\memory[14][2] ) );
  DFFPOSX1 \memory_reg[14][1]  ( .D(n1020), .CLK(CLK), .Q(\memory[14][1] ) );
  DFFPOSX1 \memory_reg[14][0]  ( .D(n1021), .CLK(CLK), .Q(\memory[14][0] ) );
  DFFPOSX1 \memory_reg[15][7]  ( .D(n1006), .CLK(CLK), .Q(\memory[15][7] ) );
  DFFPOSX1 \memory_reg[15][6]  ( .D(n1007), .CLK(CLK), .Q(\memory[15][6] ) );
  DFFPOSX1 \memory_reg[15][5]  ( .D(n1008), .CLK(CLK), .Q(\memory[15][5] ) );
  DFFPOSX1 \memory_reg[15][4]  ( .D(n1009), .CLK(CLK), .Q(\memory[15][4] ) );
  DFFPOSX1 \memory_reg[15][3]  ( .D(n1010), .CLK(CLK), .Q(\memory[15][3] ) );
  DFFPOSX1 \memory_reg[15][2]  ( .D(n1011), .CLK(CLK), .Q(\memory[15][2] ) );
  DFFPOSX1 \memory_reg[15][1]  ( .D(n1012), .CLK(CLK), .Q(\memory[15][1] ) );
  DFFPOSX1 \memory_reg[15][0]  ( .D(n1013), .CLK(CLK), .Q(\memory[15][0] ) );
  DFFPOSX1 \memory_reg[16][7]  ( .D(n1234), .CLK(CLK), .Q(\memory[16][7] ) );
  DFFPOSX1 \memory_reg[16][6]  ( .D(n1235), .CLK(CLK), .Q(\memory[16][6] ) );
  DFFPOSX1 \memory_reg[16][5]  ( .D(n1236), .CLK(CLK), .Q(\memory[16][5] ) );
  DFFPOSX1 \memory_reg[16][4]  ( .D(n1237), .CLK(CLK), .Q(\memory[16][4] ) );
  DFFPOSX1 \memory_reg[16][3]  ( .D(n1238), .CLK(CLK), .Q(\memory[16][3] ) );
  DFFPOSX1 \memory_reg[16][2]  ( .D(n1239), .CLK(CLK), .Q(\memory[16][2] ) );
  DFFPOSX1 \memory_reg[16][1]  ( .D(n1240), .CLK(CLK), .Q(\memory[16][1] ) );
  DFFPOSX1 \memory_reg[16][0]  ( .D(n1241), .CLK(CLK), .Q(\memory[16][0] ) );
  DFFPOSX1 \memory_reg[17][7]  ( .D(n1242), .CLK(CLK), .Q(\memory[17][7] ) );
  DFFPOSX1 \memory_reg[17][6]  ( .D(n1243), .CLK(CLK), .Q(\memory[17][6] ) );
  DFFPOSX1 \memory_reg[17][5]  ( .D(n1244), .CLK(CLK), .Q(\memory[17][5] ) );
  DFFPOSX1 \memory_reg[17][4]  ( .D(n1245), .CLK(CLK), .Q(\memory[17][4] ) );
  DFFPOSX1 \memory_reg[17][3]  ( .D(n1246), .CLK(CLK), .Q(\memory[17][3] ) );
  DFFPOSX1 \memory_reg[17][2]  ( .D(n1247), .CLK(CLK), .Q(\memory[17][2] ) );
  DFFPOSX1 \memory_reg[17][1]  ( .D(n1248), .CLK(CLK), .Q(\memory[17][1] ) );
  DFFPOSX1 \memory_reg[17][0]  ( .D(n1249), .CLK(CLK), .Q(\memory[17][0] ) );
  DFFPOSX1 \memory_reg[18][7]  ( .D(n1250), .CLK(CLK), .Q(\memory[18][7] ) );
  DFFPOSX1 \memory_reg[18][6]  ( .D(n1251), .CLK(CLK), .Q(\memory[18][6] ) );
  DFFPOSX1 \memory_reg[18][5]  ( .D(n1252), .CLK(CLK), .Q(\memory[18][5] ) );
  DFFPOSX1 \memory_reg[18][4]  ( .D(n1253), .CLK(CLK), .Q(\memory[18][4] ) );
  DFFPOSX1 \memory_reg[18][3]  ( .D(n1254), .CLK(CLK), .Q(\memory[18][3] ) );
  DFFPOSX1 \memory_reg[18][2]  ( .D(n1255), .CLK(CLK), .Q(\memory[18][2] ) );
  DFFPOSX1 \memory_reg[18][1]  ( .D(n1256), .CLK(CLK), .Q(\memory[18][1] ) );
  DFFPOSX1 \memory_reg[18][0]  ( .D(n1257), .CLK(CLK), .Q(\memory[18][0] ) );
  DFFPOSX1 \memory_reg[19][7]  ( .D(n1258), .CLK(CLK), .Q(\memory[19][7] ) );
  DFFPOSX1 \memory_reg[19][6]  ( .D(n1259), .CLK(CLK), .Q(\memory[19][6] ) );
  DFFPOSX1 \memory_reg[19][5]  ( .D(n1260), .CLK(CLK), .Q(\memory[19][5] ) );
  DFFPOSX1 \memory_reg[19][4]  ( .D(n1261), .CLK(CLK), .Q(\memory[19][4] ) );
  DFFPOSX1 \memory_reg[19][3]  ( .D(n1262), .CLK(CLK), .Q(\memory[19][3] ) );
  DFFPOSX1 \memory_reg[19][2]  ( .D(n1263), .CLK(CLK), .Q(\memory[19][2] ) );
  DFFPOSX1 \memory_reg[19][1]  ( .D(n1264), .CLK(CLK), .Q(\memory[19][1] ) );
  DFFPOSX1 \memory_reg[19][0]  ( .D(n1265), .CLK(CLK), .Q(\memory[19][0] ) );
  DFFPOSX1 \memory_reg[20][7]  ( .D(n998), .CLK(CLK), .Q(\memory[20][7] ) );
  DFFPOSX1 \memory_reg[20][6]  ( .D(n999), .CLK(CLK), .Q(\memory[20][6] ) );
  DFFPOSX1 \memory_reg[20][5]  ( .D(n1000), .CLK(CLK), .Q(\memory[20][5] ) );
  DFFPOSX1 \memory_reg[20][4]  ( .D(n1001), .CLK(CLK), .Q(\memory[20][4] ) );
  DFFPOSX1 \memory_reg[20][3]  ( .D(n1002), .CLK(CLK), .Q(\memory[20][3] ) );
  DFFPOSX1 \memory_reg[20][2]  ( .D(n1003), .CLK(CLK), .Q(\memory[20][2] ) );
  DFFPOSX1 \memory_reg[20][1]  ( .D(n1004), .CLK(CLK), .Q(\memory[20][1] ) );
  DFFPOSX1 \memory_reg[20][0]  ( .D(n1005), .CLK(CLK), .Q(\memory[20][0] ) );
  DFFPOSX1 \memory_reg[21][7]  ( .D(n990), .CLK(CLK), .Q(\memory[21][7] ) );
  DFFPOSX1 \memory_reg[21][6]  ( .D(n991), .CLK(CLK), .Q(\memory[21][6] ) );
  DFFPOSX1 \memory_reg[21][5]  ( .D(n992), .CLK(CLK), .Q(\memory[21][5] ) );
  DFFPOSX1 \memory_reg[21][4]  ( .D(n993), .CLK(CLK), .Q(\memory[21][4] ) );
  DFFPOSX1 \memory_reg[21][3]  ( .D(n994), .CLK(CLK), .Q(\memory[21][3] ) );
  DFFPOSX1 \memory_reg[21][2]  ( .D(n995), .CLK(CLK), .Q(\memory[21][2] ) );
  DFFPOSX1 \memory_reg[21][1]  ( .D(n996), .CLK(CLK), .Q(\memory[21][1] ) );
  DFFPOSX1 \memory_reg[21][0]  ( .D(n997), .CLK(CLK), .Q(\memory[21][0] ) );
  DFFPOSX1 \memory_reg[22][7]  ( .D(n982), .CLK(CLK), .Q(\memory[22][7] ) );
  DFFPOSX1 \memory_reg[22][6]  ( .D(n983), .CLK(CLK), .Q(\memory[22][6] ) );
  DFFPOSX1 \memory_reg[22][5]  ( .D(n984), .CLK(CLK), .Q(\memory[22][5] ) );
  DFFPOSX1 \memory_reg[22][4]  ( .D(n985), .CLK(CLK), .Q(\memory[22][4] ) );
  DFFPOSX1 \memory_reg[22][3]  ( .D(n986), .CLK(CLK), .Q(\memory[22][3] ) );
  DFFPOSX1 \memory_reg[22][2]  ( .D(n987), .CLK(CLK), .Q(\memory[22][2] ) );
  DFFPOSX1 \memory_reg[22][1]  ( .D(n988), .CLK(CLK), .Q(\memory[22][1] ) );
  DFFPOSX1 \memory_reg[22][0]  ( .D(n989), .CLK(CLK), .Q(\memory[22][0] ) );
  DFFPOSX1 \memory_reg[23][7]  ( .D(n974), .CLK(CLK), .Q(\memory[23][7] ) );
  DFFPOSX1 \memory_reg[23][6]  ( .D(n975), .CLK(CLK), .Q(\memory[23][6] ) );
  DFFPOSX1 \memory_reg[23][5]  ( .D(n976), .CLK(CLK), .Q(\memory[23][5] ) );
  DFFPOSX1 \memory_reg[23][4]  ( .D(n977), .CLK(CLK), .Q(\memory[23][4] ) );
  DFFPOSX1 \memory_reg[23][3]  ( .D(n978), .CLK(CLK), .Q(\memory[23][3] ) );
  DFFPOSX1 \memory_reg[23][2]  ( .D(n979), .CLK(CLK), .Q(\memory[23][2] ) );
  DFFPOSX1 \memory_reg[23][1]  ( .D(n980), .CLK(CLK), .Q(\memory[23][1] ) );
  DFFPOSX1 \memory_reg[23][0]  ( .D(n981), .CLK(CLK), .Q(\memory[23][0] ) );
  DFFPOSX1 \memory_reg[24][7]  ( .D(n966), .CLK(CLK), .Q(\memory[24][7] ) );
  DFFPOSX1 \memory_reg[24][6]  ( .D(n967), .CLK(CLK), .Q(\memory[24][6] ) );
  DFFPOSX1 \memory_reg[24][5]  ( .D(n968), .CLK(CLK), .Q(\memory[24][5] ) );
  DFFPOSX1 \memory_reg[24][4]  ( .D(n969), .CLK(CLK), .Q(\memory[24][4] ) );
  DFFPOSX1 \memory_reg[24][3]  ( .D(n970), .CLK(CLK), .Q(\memory[24][3] ) );
  DFFPOSX1 \memory_reg[24][2]  ( .D(n971), .CLK(CLK), .Q(\memory[24][2] ) );
  DFFPOSX1 \memory_reg[24][1]  ( .D(n972), .CLK(CLK), .Q(\memory[24][1] ) );
  DFFPOSX1 \memory_reg[24][0]  ( .D(n973), .CLK(CLK), .Q(\memory[24][0] ) );
  DFFPOSX1 \memory_reg[25][7]  ( .D(n958), .CLK(CLK), .Q(\memory[25][7] ) );
  DFFPOSX1 \memory_reg[25][6]  ( .D(n959), .CLK(CLK), .Q(\memory[25][6] ) );
  DFFPOSX1 \memory_reg[25][5]  ( .D(n960), .CLK(CLK), .Q(\memory[25][5] ) );
  DFFPOSX1 \memory_reg[25][4]  ( .D(n961), .CLK(CLK), .Q(\memory[25][4] ) );
  DFFPOSX1 \memory_reg[25][3]  ( .D(n962), .CLK(CLK), .Q(\memory[25][3] ) );
  DFFPOSX1 \memory_reg[25][2]  ( .D(n963), .CLK(CLK), .Q(\memory[25][2] ) );
  DFFPOSX1 \memory_reg[25][1]  ( .D(n964), .CLK(CLK), .Q(\memory[25][1] ) );
  DFFPOSX1 \memory_reg[25][0]  ( .D(n965), .CLK(CLK), .Q(\memory[25][0] ) );
  DFFPOSX1 \memory_reg[26][7]  ( .D(n950), .CLK(CLK), .Q(\memory[26][7] ) );
  DFFPOSX1 \memory_reg[26][6]  ( .D(n951), .CLK(CLK), .Q(\memory[26][6] ) );
  DFFPOSX1 \memory_reg[26][5]  ( .D(n952), .CLK(CLK), .Q(\memory[26][5] ) );
  DFFPOSX1 \memory_reg[26][4]  ( .D(n953), .CLK(CLK), .Q(\memory[26][4] ) );
  DFFPOSX1 \memory_reg[26][3]  ( .D(n954), .CLK(CLK), .Q(\memory[26][3] ) );
  DFFPOSX1 \memory_reg[26][2]  ( .D(n955), .CLK(CLK), .Q(\memory[26][2] ) );
  DFFPOSX1 \memory_reg[26][1]  ( .D(n956), .CLK(CLK), .Q(\memory[26][1] ) );
  DFFPOSX1 \memory_reg[26][0]  ( .D(n957), .CLK(CLK), .Q(\memory[26][0] ) );
  DFFPOSX1 \memory_reg[27][7]  ( .D(n942), .CLK(CLK), .Q(\memory[27][7] ) );
  DFFPOSX1 \memory_reg[27][6]  ( .D(n943), .CLK(CLK), .Q(\memory[27][6] ) );
  DFFPOSX1 \memory_reg[27][5]  ( .D(n944), .CLK(CLK), .Q(\memory[27][5] ) );
  DFFPOSX1 \memory_reg[27][4]  ( .D(n945), .CLK(CLK), .Q(\memory[27][4] ) );
  DFFPOSX1 \memory_reg[27][3]  ( .D(n946), .CLK(CLK), .Q(\memory[27][3] ) );
  DFFPOSX1 \memory_reg[27][2]  ( .D(n947), .CLK(CLK), .Q(\memory[27][2] ) );
  DFFPOSX1 \memory_reg[27][1]  ( .D(n948), .CLK(CLK), .Q(\memory[27][1] ) );
  DFFPOSX1 \memory_reg[27][0]  ( .D(n949), .CLK(CLK), .Q(\memory[27][0] ) );
  DFFPOSX1 \memory_reg[28][7]  ( .D(n1266), .CLK(CLK), .Q(\memory[28][7] ) );
  DFFPOSX1 \memory_reg[28][6]  ( .D(n1267), .CLK(CLK), .Q(\memory[28][6] ) );
  DFFPOSX1 \memory_reg[28][5]  ( .D(n1268), .CLK(CLK), .Q(\memory[28][5] ) );
  DFFPOSX1 \memory_reg[28][4]  ( .D(n1269), .CLK(CLK), .Q(\memory[28][4] ) );
  DFFPOSX1 \memory_reg[28][3]  ( .D(n1270), .CLK(CLK), .Q(\memory[28][3] ) );
  DFFPOSX1 \memory_reg[28][2]  ( .D(n1271), .CLK(CLK), .Q(\memory[28][2] ) );
  DFFPOSX1 \memory_reg[28][1]  ( .D(n1272), .CLK(CLK), .Q(\memory[28][1] ) );
  DFFPOSX1 \memory_reg[28][0]  ( .D(n1273), .CLK(CLK), .Q(\memory[28][0] ) );
  DFFPOSX1 \memory_reg[29][7]  ( .D(n1274), .CLK(CLK), .Q(\memory[29][7] ) );
  DFFPOSX1 \memory_reg[29][6]  ( .D(n1275), .CLK(CLK), .Q(\memory[29][6] ) );
  DFFPOSX1 \memory_reg[29][5]  ( .D(n1276), .CLK(CLK), .Q(\memory[29][5] ) );
  DFFPOSX1 \memory_reg[29][4]  ( .D(n1277), .CLK(CLK), .Q(\memory[29][4] ) );
  DFFPOSX1 \memory_reg[29][3]  ( .D(n1278), .CLK(CLK), .Q(\memory[29][3] ) );
  DFFPOSX1 \memory_reg[29][2]  ( .D(n1279), .CLK(CLK), .Q(\memory[29][2] ) );
  DFFPOSX1 \memory_reg[29][1]  ( .D(n1280), .CLK(CLK), .Q(\memory[29][1] ) );
  DFFPOSX1 \memory_reg[29][0]  ( .D(n1281), .CLK(CLK), .Q(\memory[29][0] ) );
  DFFPOSX1 \memory_reg[30][7]  ( .D(n1282), .CLK(CLK), .Q(\memory[30][7] ) );
  DFFPOSX1 \memory_reg[30][6]  ( .D(n1283), .CLK(CLK), .Q(\memory[30][6] ) );
  DFFPOSX1 \memory_reg[30][5]  ( .D(n1284), .CLK(CLK), .Q(\memory[30][5] ) );
  DFFPOSX1 \memory_reg[30][4]  ( .D(n1285), .CLK(CLK), .Q(\memory[30][4] ) );
  DFFPOSX1 \memory_reg[30][3]  ( .D(n1286), .CLK(CLK), .Q(\memory[30][3] ) );
  DFFPOSX1 \memory_reg[30][2]  ( .D(n1287), .CLK(CLK), .Q(\memory[30][2] ) );
  DFFPOSX1 \memory_reg[30][1]  ( .D(n1288), .CLK(CLK), .Q(\memory[30][1] ) );
  DFFPOSX1 \memory_reg[30][0]  ( .D(n1289), .CLK(CLK), .Q(\memory[30][0] ) );
  DFFPOSX1 \memory_reg[31][7]  ( .D(n1290), .CLK(CLK), .Q(\memory[31][7] ) );
  DFFPOSX1 \memory_reg[31][6]  ( .D(n1291), .CLK(CLK), .Q(\memory[31][6] ) );
  DFFPOSX1 \memory_reg[31][5]  ( .D(n1292), .CLK(CLK), .Q(\memory[31][5] ) );
  DFFPOSX1 \memory_reg[31][4]  ( .D(n1293), .CLK(CLK), .Q(\memory[31][4] ) );
  DFFPOSX1 \memory_reg[31][3]  ( .D(n1294), .CLK(CLK), .Q(\memory[31][3] ) );
  DFFPOSX1 \memory_reg[31][2]  ( .D(n1295), .CLK(CLK), .Q(\memory[31][2] ) );
  DFFPOSX1 \memory_reg[31][1]  ( .D(n1296), .CLK(CLK), .Q(\memory[31][1] ) );
  DFFPOSX1 \memory_reg[31][0]  ( .D(n1297), .CLK(CLK), .Q(\memory[31][0] ) );
  DFFPOSX1 \opcode_reg[0][1]  ( .D(n935), .CLK(CLK), .Q(\opcode[0][1] ) );
  DFFPOSX1 \opcode_reg[0][0]  ( .D(n934), .CLK(CLK), .Q(\opcode[0][0] ) );
  DFFPOSX1 \opcode_reg[1][1]  ( .D(n937), .CLK(CLK), .Q(\opcode[1][1] ) );
  DFFPOSX1 \opcode_reg[1][0]  ( .D(n936), .CLK(CLK), .Q(\opcode[1][0] ) );
  DFFPOSX1 \opcode_reg[2][1]  ( .D(n939), .CLK(CLK), .Q(\opcode[2][1] ) );
  DFFPOSX1 \opcode_reg[2][0]  ( .D(n938), .CLK(CLK), .Q(\opcode[2][0] ) );
  DFFPOSX1 \opcode_reg[3][1]  ( .D(n941), .CLK(CLK), .Q(\opcode[3][1] ) );
  DFFPOSX1 \opcode_reg[3][0]  ( .D(n940), .CLK(CLK), .Q(\opcode[3][0] ) );
  DFFPOSX1 \opcode_reg[4][1]  ( .D(n1363), .CLK(CLK), .Q(\opcode[4][1] ) );
  DFFPOSX1 \opcode_reg[4][0]  ( .D(n1362), .CLK(CLK), .Q(\opcode[4][0] ) );
  DFFPOSX1 \opcode_reg[5][1]  ( .D(n1353), .CLK(CLK), .Q(\opcode[5][1] ) );
  DFFPOSX1 \opcode_reg[5][0]  ( .D(n1352), .CLK(CLK), .Q(\opcode[5][0] ) );
  DFFPOSX1 \opcode_reg[6][1]  ( .D(n1343), .CLK(CLK), .Q(\opcode[6][1] ) );
  DFFPOSX1 \opcode_reg[6][0]  ( .D(n1342), .CLK(CLK), .Q(\opcode[6][0] ) );
  DFFPOSX1 \opcode_reg[7][1]  ( .D(n1333), .CLK(CLK), .Q(\opcode[7][1] ) );
  DFFPOSX1 \opcode_reg[7][0]  ( .D(n1332), .CLK(CLK), .Q(\opcode[7][0] ) );
  DFFPOSX1 \opcode_reg[8][1]  ( .D(n1298), .CLK(CLK), .Q(\opcode[8][1] ) );
  DFFPOSX1 \opcode_reg[8][0]  ( .D(n1299), .CLK(CLK), .Q(\opcode[8][0] ) );
  DFFPOSX1 \opcode_reg[9][1]  ( .D(n1300), .CLK(CLK), .Q(\opcode[9][1] ) );
  DFFPOSX1 \opcode_reg[9][0]  ( .D(n1301), .CLK(CLK), .Q(\opcode[9][0] ) );
  DFFPOSX1 \opcode_reg[10][1]  ( .D(n1302), .CLK(CLK), .Q(\opcode[10][1] ) );
  DFFPOSX1 \opcode_reg[10][0]  ( .D(n1303), .CLK(CLK), .Q(\opcode[10][0] ) );
  DFFPOSX1 \opcode_reg[11][1]  ( .D(n1304), .CLK(CLK), .Q(\opcode[11][1] ) );
  DFFPOSX1 \opcode_reg[11][0]  ( .D(n1305), .CLK(CLK), .Q(\opcode[11][0] ) );
  DFFPOSX1 \opcode_reg[12][1]  ( .D(n932), .CLK(CLK), .Q(\opcode[12][1] ) );
  DFFPOSX1 \opcode_reg[12][0]  ( .D(n933), .CLK(CLK), .Q(\opcode[12][0] ) );
  DFFPOSX1 \opcode_reg[13][1]  ( .D(n930), .CLK(CLK), .Q(\opcode[13][1] ) );
  DFFPOSX1 \opcode_reg[13][0]  ( .D(n931), .CLK(CLK), .Q(\opcode[13][0] ) );
  DFFPOSX1 \opcode_reg[14][1]  ( .D(n928), .CLK(CLK), .Q(\opcode[14][1] ) );
  DFFPOSX1 \opcode_reg[14][0]  ( .D(n929), .CLK(CLK), .Q(\opcode[14][0] ) );
  DFFPOSX1 \opcode_reg[15][1]  ( .D(n926), .CLK(CLK), .Q(\opcode[15][1] ) );
  DFFPOSX1 \opcode_reg[15][0]  ( .D(n927), .CLK(CLK), .Q(\opcode[15][0] ) );
  DFFPOSX1 \opcode_reg[16][1]  ( .D(n1306), .CLK(CLK), .Q(\opcode[16][1] ) );
  DFFPOSX1 \opcode_reg[16][0]  ( .D(n1307), .CLK(CLK), .Q(\opcode[16][0] ) );
  DFFPOSX1 \opcode_reg[17][1]  ( .D(n1308), .CLK(CLK), .Q(\opcode[17][1] ) );
  DFFPOSX1 \opcode_reg[17][0]  ( .D(n1309), .CLK(CLK), .Q(\opcode[17][0] ) );
  DFFPOSX1 \opcode_reg[18][1]  ( .D(n1310), .CLK(CLK), .Q(\opcode[18][1] ) );
  DFFPOSX1 \opcode_reg[18][0]  ( .D(n1311), .CLK(CLK), .Q(\opcode[18][0] ) );
  DFFPOSX1 \opcode_reg[19][1]  ( .D(n1312), .CLK(CLK), .Q(\opcode[19][1] ) );
  DFFPOSX1 \opcode_reg[19][0]  ( .D(n1313), .CLK(CLK), .Q(\opcode[19][0] ) );
  DFFPOSX1 \opcode_reg[20][1]  ( .D(n924), .CLK(CLK), .Q(\opcode[20][1] ) );
  DFFPOSX1 \opcode_reg[20][0]  ( .D(n925), .CLK(CLK), .Q(\opcode[20][0] ) );
  DFFPOSX1 \opcode_reg[21][1]  ( .D(n922), .CLK(CLK), .Q(\opcode[21][1] ) );
  DFFPOSX1 \opcode_reg[21][0]  ( .D(n923), .CLK(CLK), .Q(\opcode[21][0] ) );
  DFFPOSX1 \opcode_reg[22][1]  ( .D(n920), .CLK(CLK), .Q(\opcode[22][1] ) );
  DFFPOSX1 \opcode_reg[22][0]  ( .D(n921), .CLK(CLK), .Q(\opcode[22][0] ) );
  DFFPOSX1 \opcode_reg[23][1]  ( .D(n918), .CLK(CLK), .Q(\opcode[23][1] ) );
  DFFPOSX1 \opcode_reg[23][0]  ( .D(n919), .CLK(CLK), .Q(\opcode[23][0] ) );
  DFFPOSX1 \opcode_reg[24][1]  ( .D(n916), .CLK(CLK), .Q(\opcode[24][1] ) );
  DFFPOSX1 \opcode_reg[24][0]  ( .D(n917), .CLK(CLK), .Q(\opcode[24][0] ) );
  DFFPOSX1 \opcode_reg[25][1]  ( .D(n914), .CLK(CLK), .Q(\opcode[25][1] ) );
  DFFPOSX1 \opcode_reg[25][0]  ( .D(n915), .CLK(CLK), .Q(\opcode[25][0] ) );
  DFFPOSX1 \opcode_reg[26][1]  ( .D(n912), .CLK(CLK), .Q(\opcode[26][1] ) );
  DFFPOSX1 \opcode_reg[26][0]  ( .D(n913), .CLK(CLK), .Q(\opcode[26][0] ) );
  DFFPOSX1 \opcode_reg[27][1]  ( .D(n910), .CLK(CLK), .Q(\opcode[27][1] ) );
  DFFPOSX1 \opcode_reg[27][0]  ( .D(n911), .CLK(CLK), .Q(\opcode[27][0] ) );
  DFFPOSX1 \opcode_reg[28][1]  ( .D(n1314), .CLK(CLK), .Q(\opcode[28][1] ) );
  DFFPOSX1 \opcode_reg[28][0]  ( .D(n1315), .CLK(CLK), .Q(\opcode[28][0] ) );
  DFFPOSX1 \opcode_reg[29][1]  ( .D(n1316), .CLK(CLK), .Q(\opcode[29][1] ) );
  DFFPOSX1 \opcode_reg[29][0]  ( .D(n1317), .CLK(CLK), .Q(\opcode[29][0] ) );
  DFFPOSX1 \opcode_reg[30][1]  ( .D(n1318), .CLK(CLK), .Q(\opcode[30][1] ) );
  DFFPOSX1 \opcode_reg[30][0]  ( .D(n1319), .CLK(CLK), .Q(\opcode[30][0] ) );
  DFFPOSX1 \opcode_reg[31][1]  ( .D(n1320), .CLK(CLK), .Q(\opcode[31][1] ) );
  DFFPOSX1 \opcode_reg[31][0]  ( .D(n1321), .CLK(CLK), .Q(\opcode[31][0] ) );
  DFFPOSX1 \DATA_reg[7]  ( .D(n1322), .CLK(CLK), .Q(DATA[7]) );
  DFFPOSX1 \DATA_reg[6]  ( .D(n1323), .CLK(CLK), .Q(DATA[6]) );
  DFFPOSX1 \DATA_reg[5]  ( .D(n1324), .CLK(CLK), .Q(DATA[5]) );
  DFFPOSX1 \DATA_reg[4]  ( .D(n1325), .CLK(CLK), .Q(DATA[4]) );
  DFFPOSX1 \DATA_reg[3]  ( .D(n1326), .CLK(CLK), .Q(DATA[3]) );
  DFFPOSX1 \DATA_reg[2]  ( .D(n1327), .CLK(CLK), .Q(DATA[2]) );
  DFFPOSX1 \DATA_reg[1]  ( .D(n1328), .CLK(CLK), .Q(DATA[1]) );
  DFFPOSX1 \DATA_reg[0]  ( .D(n1329), .CLK(CLK), .Q(DATA[0]) );
  DFFPOSX1 \OUT_OPCODE_reg[1]  ( .D(n1330), .CLK(CLK), .Q(OUT_OPCODE[1]) );
  DFFPOSX1 \OUT_OPCODE_reg[0]  ( .D(n1331), .CLK(CLK), .Q(OUT_OPCODE[0]) );
  DFFPOSX1 EMPTY_reg ( .D(n1201), .CLK(CLK), .Q(EMPTY) );
  FAX1 \sub_72/U2_1  ( .A(n78), .B(n517), .C(\sub_72/carry[1] ), .YC(
        \sub_72/carry[2] ), .YS(N190) );
  FAX1 \sub_72/U2_2  ( .A(n76), .B(n855), .C(\sub_72/carry[2] ), .YC(
        \sub_72/carry[3] ), .YS(N191) );
  FAX1 \sub_72/U2_3  ( .A(n83), .B(n824), .C(\sub_72/carry[3] ), .YC(
        \sub_72/carry[4] ), .YS(N192) );
  FAX1 \sub_72/U2_4  ( .A(writeptr[4]), .B(n845), .C(\sub_72/carry[4] ), .YS(
        N193) );
  HAX1 \add_67/U1_1_1  ( .A(n79), .B(n81), .YC(\add_67/carry[2] ), .YS(N48) );
  HAX1 \add_67/U1_1_2  ( .A(n76), .B(\add_67/carry[2] ), .YC(\add_67/carry[3] ), .YS(N49) );
  HAX1 \add_67/U1_1_3  ( .A(n83), .B(\add_67/carry[3] ), .YC(\add_67/carry[4] ), .YS(N50) );
  HAX1 \r83/U1_1_1  ( .A(n78), .B(writeptr[0]), .YC(\r83/carry[2] ), .YS(N32)
         );
  HAX1 \r83/U1_1_2  ( .A(writeptr[2]), .B(\r83/carry[2] ), .YC(\r83/carry[3] ), 
        .YS(N33) );
  HAX1 \r83/U1_1_3  ( .A(writeptr[3]), .B(\r83/carry[3] ), .YC(\r83/carry[4] ), 
        .YS(N34) );
  DFFSR \BYTE_COUNT_reg[0]  ( .D(N338), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        BYTE_COUNT[0]) );
  DFFSR \BYTE_COUNT_reg[1]  ( .D(N339), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        BYTE_COUNT[1]) );
  DFFSR \BYTE_COUNT_reg[2]  ( .D(N340), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        BYTE_COUNT[2]) );
  DFFSR \readptr_reg[0]  ( .D(N343), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        readptr[0]) );
  DFFSR \readptr_reg[1]  ( .D(N344), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        readptr[1]) );
  DFFSR \BYTE_COUNT_reg[3]  ( .D(N341), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        BYTE_COUNT[3]) );
  DFFSR \readptr_reg[2]  ( .D(N345), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        readptr[2]) );
  DFFSR \BYTE_COUNT_reg[4]  ( .D(N342), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        BYTE_COUNT[4]) );
  DFFSR \readptr_reg[3]  ( .D(N346), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        readptr[3]) );
  DFFSR \writeptr_reg[4]  ( .D(n1373), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        writeptr[4]) );
  DFFSR \writeptr_reg[3]  ( .D(n1374), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        writeptr[3]) );
  DFFSR \writeptr_reg[2]  ( .D(n1377), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        writeptr[2]) );
  DFFSR \writeptr_reg[1]  ( .D(n1376), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        writeptr[1]) );
  DFFSR \writeptr_reg[0]  ( .D(n1375), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        writeptr[0]) );
  DFFSR \readptr_reg[4]  ( .D(N347), .CLK(CLK), .R(n98), .S(1'b1), .Q(
        readptr[4]) );
  INVX4 U3 ( .A(n55), .Y(n124) );
  OR2X1 U4 ( .A(n152), .B(n43), .Y(n55) );
  INVX4 U5 ( .A(n50), .Y(n119) );
  OR2X1 U6 ( .A(n147), .B(n43), .Y(n50) );
  INVX4 U7 ( .A(n56), .Y(n114) );
  OR2X1 U8 ( .A(n193), .B(n43), .Y(n56) );
  INVX4 U9 ( .A(n49), .Y(n435) );
  OR2X1 U10 ( .A(n244), .B(n43), .Y(n49) );
  INVX4 U11 ( .A(n57), .Y(n461) );
  OR2X1 U12 ( .A(n156), .B(n43), .Y(n57) );
  BUFX2 U13 ( .A(n218), .Y(n1) );
  INVX2 U14 ( .A(n77), .Y(n78) );
  INVX2 U15 ( .A(n503), .Y(n109) );
  BUFX2 U16 ( .A(n452), .Y(n74) );
  INVX2 U17 ( .A(n23), .Y(n73) );
  INVX2 U18 ( .A(n6), .Y(n58) );
  INVX2 U19 ( .A(n11), .Y(n59) );
  INVX2 U20 ( .A(n12), .Y(n60) );
  INVX2 U21 ( .A(n14), .Y(n72) );
  INVX2 U22 ( .A(n3), .Y(n71) );
  INVX2 U23 ( .A(n4), .Y(n70) );
  INVX2 U24 ( .A(n13), .Y(n69) );
  INVX2 U25 ( .A(n24), .Y(n65) );
  INVX2 U26 ( .A(n10), .Y(n66) );
  INVX2 U27 ( .A(n15), .Y(n67) );
  INVX2 U28 ( .A(n25), .Y(n68) );
  INVX2 U29 ( .A(n7), .Y(n64) );
  INVX2 U30 ( .A(n9), .Y(n63) );
  INVX2 U31 ( .A(n26), .Y(n62) );
  INVX2 U32 ( .A(n8), .Y(n61) );
  AND2X2 U33 ( .A(n483), .B(n361), .Y(n2) );
  OR2X2 U34 ( .A(n1), .B(n193), .Y(n3) );
  OR2X2 U35 ( .A(n1), .B(n147), .Y(n4) );
  AND2X2 U36 ( .A(n496), .B(n82), .Y(n5) );
  OR2X2 U37 ( .A(n43), .B(n184), .Y(n6) );
  OR2X2 U38 ( .A(n44), .B(n184), .Y(n7) );
  OR2X2 U39 ( .A(n45), .B(n152), .Y(n8) );
  OR2X2 U40 ( .A(n44), .B(n193), .Y(n9) );
  OR2X2 U41 ( .A(n46), .B(n161), .Y(n10) );
  OR2X2 U42 ( .A(n1), .B(n235), .Y(n11) );
  OR2X2 U43 ( .A(n1), .B(n244), .Y(n12) );
  OR2X2 U44 ( .A(n1), .B(n152), .Y(n13) );
  OR2X2 U45 ( .A(n1), .B(n184), .Y(n14) );
  OR2X2 U46 ( .A(n46), .B(n235), .Y(n15) );
  NAND2X1 U47 ( .A(n253), .B(n128), .Y(n16) );
  NAND2X1 U48 ( .A(n253), .B(n138), .Y(n17) );
  NAND2X1 U49 ( .A(n253), .B(n143), .Y(n18) );
  NAND2X1 U50 ( .A(n253), .B(n123), .Y(n19) );
  NAND2X1 U51 ( .A(n253), .B(n108), .Y(n20) );
  NAND2X1 U52 ( .A(n253), .B(n133), .Y(n21) );
  NAND2X1 U53 ( .A(n253), .B(n113), .Y(n22) );
  OR2X2 U54 ( .A(n43), .B(n235), .Y(n23) );
  OR2X2 U55 ( .A(n45), .B(n156), .Y(n24) );
  OR2X2 U56 ( .A(n44), .B(n244), .Y(n25) );
  OR2X2 U57 ( .A(n45), .B(n147), .Y(n26) );
  AND2X2 U58 ( .A(n496), .B(n83), .Y(n27) );
  INVX2 U59 ( .A(n106), .Y(n89) );
  BUFX2 U75 ( .A(n183), .Y(n43) );
  NAND2X1 U76 ( .A(n47), .B(n27), .Y(n183) );
  NAND2X1 U77 ( .A(n47), .B(n5), .Y(n218) );
  OR2X2 U78 ( .A(n156), .B(n1), .Y(n48) );
  INVX2 U79 ( .A(n148), .Y(n139) );
  INVX2 U80 ( .A(n510), .Y(n361) );
  INVX2 U81 ( .A(n511), .Y(n165) );
  BUFX2 U82 ( .A(n286), .Y(n44) );
  BUFX2 U83 ( .A(n286), .Y(n45) );
  BUFX2 U84 ( .A(n286), .Y(n46) );
  NOR2X1 U85 ( .A(n510), .B(n483), .Y(n47) );
  INVX2 U86 ( .A(writeptr[2]), .Y(n75) );
  INVX2 U87 ( .A(n89), .Y(n88) );
  INVX4 U88 ( .A(n48), .Y(n129) );
  INVX4 U89 ( .A(n54), .Y(n134) );
  XNOR2X1 U90 ( .A(readptr[0]), .B(n81), .Y(n519) );
  INVX2 U91 ( .A(RST), .Y(n98) );
  INVX2 U92 ( .A(n82), .Y(n83) );
  INVX2 U93 ( .A(n75), .Y(n76) );
  INVX2 U94 ( .A(RCV_DATA[7]), .Y(n90) );
  INVX2 U95 ( .A(RCV_DATA[1]), .Y(n96) );
  INVX2 U96 ( .A(RCV_DATA[3]), .Y(n94) );
  INVX2 U97 ( .A(RCV_DATA[5]), .Y(n92) );
  INVX2 U98 ( .A(RCV_DATA[0]), .Y(n97) );
  INVX2 U99 ( .A(RCV_DATA[2]), .Y(n95) );
  INVX2 U100 ( .A(RCV_DATA[4]), .Y(n93) );
  INVX2 U101 ( .A(RCV_DATA[6]), .Y(n91) );
  XNOR2X1 U102 ( .A(readptr[4]), .B(n51), .Y(n516) );
  XNOR2X1 U103 ( .A(\r83/carry[4] ), .B(writeptr[4]), .Y(n51) );
  INVX2 U104 ( .A(writeptr[3]), .Y(n82) );
  BUFX2 U105 ( .A(state), .Y(n84) );
  INVX1 U106 ( .A(n80), .Y(n81) );
  INVX2 U107 ( .A(writeptr[0]), .Y(n80) );
  INVX1 U108 ( .A(n47), .Y(n52) );
  INVX2 U109 ( .A(n52), .Y(n53) );
  INVX1 U110 ( .A(n77), .Y(n79) );
  INVX1 U111 ( .A(writeptr[1]), .Y(n77) );
  OR2X2 U112 ( .A(n161), .B(n1), .Y(n54) );
  INVX1 U113 ( .A(RCV_OPCODE[0]), .Y(n106) );
  AND2X2 U114 ( .A(RCV_OPCODE[1]), .B(n89), .Y(n483) );
  INVX1 U115 ( .A(RCV_OPCODE[1]), .Y(n87) );
  INVX1 U116 ( .A(RCV_OPCODE[1]), .Y(n86) );
  INVX1 U117 ( .A(RCV_OPCODE[1]), .Y(n85) );
  AND2X2 U118 ( .A(n478), .B(n47), .Y(n253) );
  AND2X2 U119 ( .A(n253), .B(n118), .Y(n394) );
  AND2X2 U120 ( .A(n818), .B(n820), .Y(n537) );
  AND2X2 U121 ( .A(n816), .B(n820), .Y(n536) );
  AND2X2 U122 ( .A(n818), .B(n821), .Y(n539) );
  AND2X2 U123 ( .A(n816), .B(n821), .Y(n538) );
  AND2X2 U124 ( .A(n832), .B(n820), .Y(n550) );
  AND2X2 U125 ( .A(n820), .B(n831), .Y(n549) );
  AND2X2 U126 ( .A(n821), .B(n832), .Y(n552) );
  AND2X2 U127 ( .A(n821), .B(n831), .Y(n551) );
  AND2X2 U128 ( .A(n843), .B(n821), .Y(n565) );
  AND2X2 U129 ( .A(n842), .B(n821), .Y(n564) );
  AND2X2 U130 ( .A(n843), .B(n820), .Y(n567) );
  AND2X2 U131 ( .A(n842), .B(n820), .Y(n566) );
  AND2X2 U132 ( .A(n853), .B(n820), .Y(n578) );
  AND2X2 U133 ( .A(n852), .B(n820), .Y(n577) );
  AND2X2 U134 ( .A(n853), .B(n821), .Y(n580) );
  AND2X2 U135 ( .A(n852), .B(n821), .Y(n579) );
  OR2X1 U136 ( .A(n823), .B(n81), .Y(\sub_72/carry[1] ) );
  XNOR2X1 U137 ( .A(writeptr[0]), .B(n823), .Y(N189) );
  XOR2X1 U138 ( .A(readptr[4]), .B(\add_76_aco/carry[4] ), .Y(N337) );
  AND2X1 U139 ( .A(readptr[3]), .B(\add_76_aco/carry[3] ), .Y(
        \add_76_aco/carry[4] ) );
  XOR2X1 U140 ( .A(\add_76_aco/carry[3] ), .B(readptr[3]), .Y(N336) );
  AND2X1 U141 ( .A(readptr[2]), .B(\add_76_aco/carry[2] ), .Y(
        \add_76_aco/carry[3] ) );
  XOR2X1 U142 ( .A(\add_76_aco/carry[2] ), .B(readptr[2]), .Y(N335) );
  AND2X1 U143 ( .A(readptr[1]), .B(\add_76_aco/carry[1] ), .Y(
        \add_76_aco/carry[2] ) );
  XOR2X1 U144 ( .A(\add_76_aco/carry[1] ), .B(readptr[1]), .Y(N334) );
  AND2X1 U145 ( .A(readptr[0]), .B(N195), .Y(\add_76_aco/carry[1] ) );
  XOR2X1 U146 ( .A(N195), .B(readptr[0]), .Y(N333) );
  NOR2X1 U147 ( .A(n79), .B(n81), .Y(n100) );
  AOI21X1 U148 ( .A(n81), .B(n79), .C(n100), .Y(n99) );
  NAND2X1 U149 ( .A(n100), .B(n75), .Y(n101) );
  OAI21X1 U150 ( .A(n100), .B(n75), .C(n101), .Y(N44) );
  XNOR2X1 U151 ( .A(n83), .B(n101), .Y(N45) );
  NOR2X1 U152 ( .A(n83), .B(n101), .Y(n102) );
  XOR2X1 U153 ( .A(writeptr[4]), .B(n102), .Y(N46) );
  INVX2 U154 ( .A(n99), .Y(N43) );
  XOR2X1 U155 ( .A(\add_67/carry[4] ), .B(writeptr[4]), .Y(N51) );
  MUX2X1 U156 ( .B(n86), .A(n104), .S(n105), .Y(n910) );
  MUX2X1 U157 ( .B(n88), .A(n107), .S(n105), .Y(n911) );
  AOI21X1 U158 ( .A(n108), .B(n109), .C(n58), .Y(n105) );
  MUX2X1 U159 ( .B(n85), .A(n110), .S(n111), .Y(n912) );
  MUX2X1 U160 ( .B(n88), .A(n112), .S(n111), .Y(n913) );
  AOI21X1 U161 ( .A(n109), .B(n113), .C(n114), .Y(n111) );
  MUX2X1 U162 ( .B(n85), .A(n115), .S(n116), .Y(n914) );
  MUX2X1 U163 ( .B(n88), .A(n117), .S(n116), .Y(n915) );
  AOI21X1 U164 ( .A(n109), .B(n118), .C(n119), .Y(n116) );
  MUX2X1 U165 ( .B(n85), .A(n120), .S(n121), .Y(n916) );
  MUX2X1 U166 ( .B(n88), .A(n122), .S(n121), .Y(n917) );
  AOI21X1 U167 ( .A(n109), .B(n123), .C(n124), .Y(n121) );
  MUX2X1 U168 ( .B(n85), .A(n125), .S(n126), .Y(n918) );
  INVX1 U169 ( .A(\opcode[23][1] ), .Y(n125) );
  MUX2X1 U170 ( .B(n88), .A(n127), .S(n126), .Y(n919) );
  AOI21X1 U171 ( .A(n109), .B(n128), .C(n129), .Y(n126) );
  INVX1 U172 ( .A(\opcode[23][0] ), .Y(n127) );
  MUX2X1 U173 ( .B(n85), .A(n130), .S(n131), .Y(n920) );
  INVX1 U174 ( .A(\opcode[22][1] ), .Y(n130) );
  MUX2X1 U175 ( .B(n88), .A(n132), .S(n131), .Y(n921) );
  AOI21X1 U176 ( .A(n109), .B(n133), .C(n134), .Y(n131) );
  INVX1 U177 ( .A(\opcode[22][0] ), .Y(n132) );
  MUX2X1 U178 ( .B(n85), .A(n135), .S(n136), .Y(n922) );
  INVX1 U179 ( .A(\opcode[21][1] ), .Y(n135) );
  MUX2X1 U180 ( .B(n88), .A(n137), .S(n136), .Y(n923) );
  AOI21X1 U181 ( .A(n138), .B(n139), .C(n59), .Y(n136) );
  INVX1 U182 ( .A(\opcode[21][0] ), .Y(n137) );
  MUX2X1 U183 ( .B(n85), .A(n140), .S(n141), .Y(n924) );
  INVX1 U184 ( .A(\opcode[20][1] ), .Y(n140) );
  MUX2X1 U185 ( .B(n88), .A(n142), .S(n141), .Y(n925) );
  AOI21X1 U186 ( .A(n143), .B(n139), .C(n60), .Y(n141) );
  INVX1 U187 ( .A(\opcode[20][0] ), .Y(n142) );
  INVX1 U188 ( .A(n144), .Y(n926) );
  MUX2X1 U189 ( .B(\opcode[15][1] ), .A(RCV_OPCODE[1]), .S(n145), .Y(n144) );
  INVX1 U190 ( .A(n146), .Y(n927) );
  MUX2X1 U191 ( .B(\opcode[15][0] ), .A(RCV_OPCODE[0]), .S(n145), .Y(n146) );
  OAI21X1 U192 ( .A(n147), .B(n148), .C(n17), .Y(n145) );
  INVX1 U193 ( .A(n149), .Y(n928) );
  MUX2X1 U194 ( .B(\opcode[14][1] ), .A(RCV_OPCODE[1]), .S(n150), .Y(n149) );
  INVX1 U195 ( .A(n151), .Y(n929) );
  MUX2X1 U196 ( .B(\opcode[14][0] ), .A(RCV_OPCODE[0]), .S(n150), .Y(n151) );
  OAI21X1 U197 ( .A(n152), .B(n148), .C(n18), .Y(n150) );
  MUX2X1 U198 ( .B(n153), .A(n87), .S(n154), .Y(n930) );
  INVX1 U199 ( .A(\opcode[13][1] ), .Y(n153) );
  MUX2X1 U200 ( .B(n155), .A(n88), .S(n154), .Y(n931) );
  OAI21X1 U201 ( .A(n156), .B(n157), .C(n20), .Y(n154) );
  INVX1 U202 ( .A(\opcode[13][0] ), .Y(n155) );
  MUX2X1 U203 ( .B(n158), .A(n87), .S(n159), .Y(n932) );
  INVX1 U204 ( .A(\opcode[12][1] ), .Y(n158) );
  MUX2X1 U205 ( .B(n160), .A(n88), .S(n159), .Y(n933) );
  OAI21X1 U206 ( .A(n161), .B(n157), .C(n22), .Y(n159) );
  INVX1 U207 ( .A(\opcode[12][0] ), .Y(n160) );
  MUX2X1 U208 ( .B(n88), .A(n162), .S(n163), .Y(n934) );
  MUX2X1 U209 ( .B(n85), .A(n164), .S(n163), .Y(n935) );
  AOI21X1 U210 ( .A(n123), .B(n165), .C(n61), .Y(n163) );
  MUX2X1 U211 ( .B(n88), .A(n166), .S(n167), .Y(n936) );
  MUX2X1 U212 ( .B(n85), .A(n168), .S(n167), .Y(n937) );
  AOI21X1 U213 ( .A(n118), .B(n165), .C(n62), .Y(n167) );
  MUX2X1 U214 ( .B(n88), .A(n169), .S(n170), .Y(n938) );
  MUX2X1 U215 ( .B(n85), .A(n171), .S(n170), .Y(n939) );
  AOI21X1 U216 ( .A(n113), .B(n165), .C(n63), .Y(n170) );
  MUX2X1 U217 ( .B(n88), .A(n172), .S(n173), .Y(n940) );
  MUX2X1 U218 ( .B(n85), .A(n174), .S(n173), .Y(n941) );
  AOI21X1 U219 ( .A(n108), .B(n165), .C(n64), .Y(n173) );
  MUX2X1 U220 ( .B(n175), .A(n90), .S(n58), .Y(n942) );
  MUX2X1 U221 ( .B(n176), .A(n91), .S(n58), .Y(n943) );
  MUX2X1 U222 ( .B(n177), .A(n92), .S(n58), .Y(n944) );
  MUX2X1 U223 ( .B(n178), .A(n93), .S(n58), .Y(n945) );
  MUX2X1 U224 ( .B(n179), .A(n94), .S(n58), .Y(n946) );
  MUX2X1 U225 ( .B(n180), .A(n95), .S(n58), .Y(n947) );
  MUX2X1 U226 ( .B(n181), .A(n96), .S(n58), .Y(n948) );
  MUX2X1 U227 ( .B(n182), .A(n97), .S(n58), .Y(n949) );
  MUX2X1 U228 ( .B(n185), .A(n90), .S(n114), .Y(n950) );
  MUX2X1 U229 ( .B(n186), .A(n91), .S(n114), .Y(n951) );
  MUX2X1 U230 ( .B(n187), .A(n92), .S(n114), .Y(n952) );
  MUX2X1 U231 ( .B(n188), .A(n93), .S(n114), .Y(n953) );
  MUX2X1 U232 ( .B(n189), .A(n94), .S(n114), .Y(n954) );
  MUX2X1 U233 ( .B(n190), .A(n95), .S(n114), .Y(n955) );
  MUX2X1 U234 ( .B(n191), .A(n96), .S(n114), .Y(n956) );
  MUX2X1 U235 ( .B(n192), .A(n97), .S(n114), .Y(n957) );
  MUX2X1 U236 ( .B(n194), .A(n90), .S(n119), .Y(n958) );
  MUX2X1 U237 ( .B(n195), .A(n91), .S(n119), .Y(n959) );
  MUX2X1 U238 ( .B(n196), .A(n92), .S(n119), .Y(n960) );
  MUX2X1 U239 ( .B(n197), .A(n93), .S(n119), .Y(n961) );
  MUX2X1 U240 ( .B(n198), .A(n94), .S(n119), .Y(n962) );
  MUX2X1 U241 ( .B(n199), .A(n95), .S(n119), .Y(n963) );
  MUX2X1 U242 ( .B(n200), .A(n96), .S(n119), .Y(n964) );
  MUX2X1 U243 ( .B(n201), .A(n97), .S(n119), .Y(n965) );
  MUX2X1 U244 ( .B(n202), .A(n90), .S(n124), .Y(n966) );
  MUX2X1 U245 ( .B(n203), .A(n91), .S(n124), .Y(n967) );
  MUX2X1 U246 ( .B(n204), .A(n92), .S(n124), .Y(n968) );
  MUX2X1 U247 ( .B(n205), .A(n93), .S(n124), .Y(n969) );
  MUX2X1 U248 ( .B(n206), .A(n94), .S(n124), .Y(n970) );
  MUX2X1 U249 ( .B(n207), .A(n95), .S(n124), .Y(n971) );
  MUX2X1 U250 ( .B(n208), .A(n96), .S(n124), .Y(n972) );
  MUX2X1 U251 ( .B(n209), .A(n97), .S(n124), .Y(n973) );
  MUX2X1 U252 ( .B(n210), .A(n90), .S(n129), .Y(n974) );
  INVX1 U253 ( .A(\memory[23][7] ), .Y(n210) );
  MUX2X1 U254 ( .B(n211), .A(n91), .S(n129), .Y(n975) );
  INVX1 U255 ( .A(\memory[23][6] ), .Y(n211) );
  MUX2X1 U256 ( .B(n212), .A(n92), .S(n129), .Y(n976) );
  INVX1 U257 ( .A(\memory[23][5] ), .Y(n212) );
  MUX2X1 U258 ( .B(n213), .A(n93), .S(n129), .Y(n977) );
  INVX1 U259 ( .A(\memory[23][4] ), .Y(n213) );
  MUX2X1 U260 ( .B(n214), .A(n94), .S(n129), .Y(n978) );
  INVX1 U261 ( .A(\memory[23][3] ), .Y(n214) );
  MUX2X1 U262 ( .B(n215), .A(n95), .S(n129), .Y(n979) );
  INVX1 U263 ( .A(\memory[23][2] ), .Y(n215) );
  MUX2X1 U264 ( .B(n216), .A(n96), .S(n129), .Y(n980) );
  INVX1 U265 ( .A(\memory[23][1] ), .Y(n216) );
  MUX2X1 U266 ( .B(n217), .A(n97), .S(n129), .Y(n981) );
  INVX1 U267 ( .A(\memory[23][0] ), .Y(n217) );
  MUX2X1 U268 ( .B(n219), .A(n90), .S(n134), .Y(n982) );
  INVX1 U269 ( .A(\memory[22][7] ), .Y(n219) );
  MUX2X1 U270 ( .B(n220), .A(n91), .S(n134), .Y(n983) );
  INVX1 U271 ( .A(\memory[22][6] ), .Y(n220) );
  MUX2X1 U272 ( .B(n221), .A(n92), .S(n134), .Y(n984) );
  INVX1 U273 ( .A(\memory[22][5] ), .Y(n221) );
  MUX2X1 U274 ( .B(n222), .A(n93), .S(n134), .Y(n985) );
  INVX1 U275 ( .A(\memory[22][4] ), .Y(n222) );
  MUX2X1 U276 ( .B(n223), .A(n94), .S(n134), .Y(n986) );
  INVX1 U277 ( .A(\memory[22][3] ), .Y(n223) );
  MUX2X1 U278 ( .B(n224), .A(n95), .S(n134), .Y(n987) );
  INVX1 U279 ( .A(\memory[22][2] ), .Y(n224) );
  MUX2X1 U280 ( .B(n225), .A(n96), .S(n134), .Y(n988) );
  INVX1 U281 ( .A(\memory[22][1] ), .Y(n225) );
  MUX2X1 U282 ( .B(n226), .A(n97), .S(n134), .Y(n989) );
  INVX1 U283 ( .A(\memory[22][0] ), .Y(n226) );
  MUX2X1 U284 ( .B(n227), .A(n90), .S(n59), .Y(n990) );
  INVX1 U285 ( .A(\memory[21][7] ), .Y(n227) );
  MUX2X1 U286 ( .B(n228), .A(n91), .S(n59), .Y(n991) );
  INVX1 U287 ( .A(\memory[21][6] ), .Y(n228) );
  MUX2X1 U288 ( .B(n229), .A(n92), .S(n59), .Y(n992) );
  INVX1 U289 ( .A(\memory[21][5] ), .Y(n229) );
  MUX2X1 U290 ( .B(n230), .A(n93), .S(n59), .Y(n993) );
  INVX1 U291 ( .A(\memory[21][4] ), .Y(n230) );
  MUX2X1 U292 ( .B(n231), .A(n94), .S(n59), .Y(n994) );
  INVX1 U293 ( .A(\memory[21][3] ), .Y(n231) );
  MUX2X1 U294 ( .B(n232), .A(n95), .S(n59), .Y(n995) );
  INVX1 U295 ( .A(\memory[21][2] ), .Y(n232) );
  MUX2X1 U296 ( .B(n233), .A(n96), .S(n59), .Y(n996) );
  INVX1 U297 ( .A(\memory[21][1] ), .Y(n233) );
  MUX2X1 U298 ( .B(n234), .A(n97), .S(n59), .Y(n997) );
  INVX1 U299 ( .A(\memory[21][0] ), .Y(n234) );
  MUX2X1 U300 ( .B(n236), .A(n90), .S(n60), .Y(n998) );
  INVX1 U301 ( .A(\memory[20][7] ), .Y(n236) );
  MUX2X1 U302 ( .B(n237), .A(n91), .S(n60), .Y(n999) );
  INVX1 U303 ( .A(\memory[20][6] ), .Y(n237) );
  MUX2X1 U304 ( .B(n238), .A(n92), .S(n60), .Y(n1000) );
  INVX1 U305 ( .A(\memory[20][5] ), .Y(n238) );
  MUX2X1 U306 ( .B(n239), .A(n93), .S(n60), .Y(n1001) );
  INVX1 U307 ( .A(\memory[20][4] ), .Y(n239) );
  MUX2X1 U308 ( .B(n240), .A(n94), .S(n60), .Y(n1002) );
  INVX1 U309 ( .A(\memory[20][3] ), .Y(n240) );
  MUX2X1 U310 ( .B(n241), .A(n95), .S(n60), .Y(n1003) );
  INVX1 U311 ( .A(\memory[20][2] ), .Y(n241) );
  MUX2X1 U312 ( .B(n242), .A(n96), .S(n60), .Y(n1004) );
  INVX1 U313 ( .A(\memory[20][1] ), .Y(n242) );
  MUX2X1 U314 ( .B(n243), .A(n97), .S(n60), .Y(n1005) );
  INVX1 U315 ( .A(\memory[20][0] ), .Y(n243) );
  MUX2X1 U316 ( .B(n90), .A(n245), .S(n17), .Y(n1006) );
  INVX1 U317 ( .A(\memory[15][7] ), .Y(n245) );
  MUX2X1 U318 ( .B(n91), .A(n246), .S(n17), .Y(n1007) );
  INVX1 U319 ( .A(\memory[15][6] ), .Y(n246) );
  MUX2X1 U320 ( .B(n92), .A(n247), .S(n17), .Y(n1008) );
  INVX1 U321 ( .A(\memory[15][5] ), .Y(n247) );
  MUX2X1 U322 ( .B(n93), .A(n248), .S(n17), .Y(n1009) );
  INVX1 U323 ( .A(\memory[15][4] ), .Y(n248) );
  MUX2X1 U324 ( .B(n94), .A(n249), .S(n17), .Y(n1010) );
  INVX1 U325 ( .A(\memory[15][3] ), .Y(n249) );
  MUX2X1 U326 ( .B(n95), .A(n250), .S(n17), .Y(n1011) );
  INVX1 U327 ( .A(\memory[15][2] ), .Y(n250) );
  MUX2X1 U328 ( .B(n96), .A(n251), .S(n17), .Y(n1012) );
  INVX1 U329 ( .A(\memory[15][1] ), .Y(n251) );
  MUX2X1 U330 ( .B(n97), .A(n252), .S(n17), .Y(n1013) );
  INVX1 U331 ( .A(\memory[15][0] ), .Y(n252) );
  MUX2X1 U332 ( .B(n90), .A(n254), .S(n18), .Y(n1014) );
  INVX1 U333 ( .A(\memory[14][7] ), .Y(n254) );
  MUX2X1 U334 ( .B(n91), .A(n255), .S(n18), .Y(n1015) );
  INVX1 U335 ( .A(\memory[14][6] ), .Y(n255) );
  MUX2X1 U336 ( .B(n92), .A(n256), .S(n18), .Y(n1016) );
  INVX1 U337 ( .A(\memory[14][5] ), .Y(n256) );
  MUX2X1 U338 ( .B(n93), .A(n257), .S(n18), .Y(n1017) );
  INVX1 U339 ( .A(\memory[14][4] ), .Y(n257) );
  MUX2X1 U340 ( .B(n94), .A(n258), .S(n18), .Y(n1018) );
  INVX1 U341 ( .A(\memory[14][3] ), .Y(n258) );
  MUX2X1 U342 ( .B(n95), .A(n259), .S(n18), .Y(n1019) );
  INVX1 U343 ( .A(\memory[14][2] ), .Y(n259) );
  MUX2X1 U344 ( .B(n96), .A(n260), .S(n18), .Y(n1020) );
  INVX1 U345 ( .A(\memory[14][1] ), .Y(n260) );
  MUX2X1 U346 ( .B(n97), .A(n261), .S(n18), .Y(n1021) );
  INVX1 U347 ( .A(\memory[14][0] ), .Y(n261) );
  MUX2X1 U348 ( .B(n90), .A(n262), .S(n20), .Y(n1022) );
  INVX1 U349 ( .A(\memory[13][7] ), .Y(n262) );
  MUX2X1 U350 ( .B(n91), .A(n263), .S(n20), .Y(n1023) );
  INVX1 U351 ( .A(\memory[13][6] ), .Y(n263) );
  MUX2X1 U352 ( .B(n92), .A(n264), .S(n20), .Y(n1024) );
  INVX1 U353 ( .A(\memory[13][5] ), .Y(n264) );
  MUX2X1 U354 ( .B(n93), .A(n265), .S(n20), .Y(n1025) );
  INVX1 U355 ( .A(\memory[13][4] ), .Y(n265) );
  MUX2X1 U356 ( .B(n94), .A(n266), .S(n20), .Y(n1026) );
  INVX1 U357 ( .A(\memory[13][3] ), .Y(n266) );
  MUX2X1 U358 ( .B(n95), .A(n267), .S(n20), .Y(n1027) );
  INVX1 U359 ( .A(\memory[13][2] ), .Y(n267) );
  MUX2X1 U360 ( .B(n96), .A(n268), .S(n20), .Y(n1028) );
  INVX1 U361 ( .A(\memory[13][1] ), .Y(n268) );
  MUX2X1 U362 ( .B(n97), .A(n269), .S(n20), .Y(n1029) );
  INVX1 U363 ( .A(\memory[13][0] ), .Y(n269) );
  MUX2X1 U364 ( .B(n90), .A(n270), .S(n22), .Y(n1064) );
  INVX1 U365 ( .A(\memory[12][7] ), .Y(n270) );
  MUX2X1 U366 ( .B(n91), .A(n271), .S(n22), .Y(n1065) );
  INVX1 U367 ( .A(\memory[12][6] ), .Y(n271) );
  MUX2X1 U368 ( .B(n92), .A(n272), .S(n22), .Y(n1066) );
  INVX1 U369 ( .A(\memory[12][5] ), .Y(n272) );
  MUX2X1 U370 ( .B(n93), .A(n273), .S(n22), .Y(n1067) );
  INVX1 U371 ( .A(\memory[12][4] ), .Y(n273) );
  MUX2X1 U372 ( .B(n94), .A(n274), .S(n22), .Y(n1068) );
  INVX1 U373 ( .A(\memory[12][3] ), .Y(n274) );
  MUX2X1 U374 ( .B(n95), .A(n275), .S(n22), .Y(n1069) );
  INVX1 U375 ( .A(\memory[12][2] ), .Y(n275) );
  MUX2X1 U376 ( .B(n96), .A(n276), .S(n22), .Y(n1070) );
  INVX1 U377 ( .A(\memory[12][1] ), .Y(n276) );
  MUX2X1 U378 ( .B(n97), .A(n277), .S(n22), .Y(n1071) );
  INVX1 U379 ( .A(\memory[12][0] ), .Y(n277) );
  MUX2X1 U380 ( .B(n278), .A(n97), .S(n61), .Y(n1168) );
  MUX2X1 U381 ( .B(n279), .A(n96), .S(n61), .Y(n1169) );
  MUX2X1 U382 ( .B(n280), .A(n95), .S(n61), .Y(n1170) );
  MUX2X1 U383 ( .B(n281), .A(n94), .S(n61), .Y(n1171) );
  MUX2X1 U384 ( .B(n282), .A(n93), .S(n61), .Y(n1172) );
  MUX2X1 U385 ( .B(n283), .A(n92), .S(n61), .Y(n1173) );
  MUX2X1 U386 ( .B(n284), .A(n91), .S(n61), .Y(n1174) );
  MUX2X1 U387 ( .B(n285), .A(n90), .S(n61), .Y(n1175) );
  MUX2X1 U388 ( .B(n287), .A(n97), .S(n62), .Y(n1176) );
  MUX2X1 U389 ( .B(n288), .A(n96), .S(n62), .Y(n1177) );
  MUX2X1 U390 ( .B(n289), .A(n95), .S(n62), .Y(n1178) );
  MUX2X1 U391 ( .B(n290), .A(n94), .S(n62), .Y(n1179) );
  MUX2X1 U392 ( .B(n291), .A(n93), .S(n62), .Y(n1180) );
  MUX2X1 U393 ( .B(n292), .A(n92), .S(n62), .Y(n1181) );
  MUX2X1 U394 ( .B(n293), .A(n91), .S(n62), .Y(n1182) );
  MUX2X1 U395 ( .B(n294), .A(n90), .S(n62), .Y(n1183) );
  MUX2X1 U396 ( .B(n295), .A(n97), .S(n63), .Y(n1184) );
  MUX2X1 U397 ( .B(n296), .A(n96), .S(n63), .Y(n1185) );
  MUX2X1 U398 ( .B(n297), .A(n95), .S(n63), .Y(n1186) );
  MUX2X1 U399 ( .B(n298), .A(n94), .S(n63), .Y(n1187) );
  MUX2X1 U400 ( .B(n299), .A(n93), .S(n63), .Y(n1188) );
  MUX2X1 U401 ( .B(n300), .A(n92), .S(n63), .Y(n1189) );
  MUX2X1 U402 ( .B(n301), .A(n91), .S(n63), .Y(n1190) );
  MUX2X1 U403 ( .B(n302), .A(n90), .S(n63), .Y(n1191) );
  MUX2X1 U404 ( .B(n303), .A(n97), .S(n64), .Y(n1192) );
  MUX2X1 U405 ( .B(n304), .A(n96), .S(n64), .Y(n1193) );
  MUX2X1 U406 ( .B(n305), .A(n95), .S(n64), .Y(n1194) );
  MUX2X1 U407 ( .B(n306), .A(n94), .S(n64), .Y(n1195) );
  MUX2X1 U408 ( .B(n307), .A(n93), .S(n64), .Y(n1196) );
  MUX2X1 U409 ( .B(n308), .A(n92), .S(n64), .Y(n1197) );
  MUX2X1 U410 ( .B(n309), .A(n91), .S(n64), .Y(n1198) );
  MUX2X1 U411 ( .B(n310), .A(n90), .S(n64), .Y(n1199) );
  MUX2X1 U412 ( .B(n311), .A(n312), .S(RST), .Y(n1200) );
  INVX1 U413 ( .A(FULL), .Y(n312) );
  MUX2X1 U414 ( .B(n313), .A(n314), .S(RST), .Y(n1201) );
  INVX1 U415 ( .A(EMPTY), .Y(n314) );
  MUX2X1 U416 ( .B(n88), .A(n315), .S(n316), .Y(n1332) );
  INVX1 U417 ( .A(\opcode[7][0] ), .Y(n315) );
  MUX2X1 U418 ( .B(n85), .A(n317), .S(n316), .Y(n1333) );
  AOI21X1 U419 ( .A(n128), .B(n318), .C(n65), .Y(n316) );
  INVX1 U420 ( .A(\opcode[7][1] ), .Y(n317) );
  MUX2X1 U421 ( .B(n319), .A(n97), .S(n65), .Y(n1334) );
  INVX1 U422 ( .A(\memory[7][0] ), .Y(n319) );
  MUX2X1 U423 ( .B(n320), .A(n96), .S(n65), .Y(n1335) );
  INVX1 U424 ( .A(\memory[7][1] ), .Y(n320) );
  MUX2X1 U425 ( .B(n321), .A(n95), .S(n65), .Y(n1336) );
  INVX1 U426 ( .A(\memory[7][2] ), .Y(n321) );
  MUX2X1 U427 ( .B(n322), .A(n94), .S(n65), .Y(n1337) );
  INVX1 U428 ( .A(\memory[7][3] ), .Y(n322) );
  MUX2X1 U429 ( .B(n323), .A(n93), .S(n65), .Y(n1338) );
  INVX1 U430 ( .A(\memory[7][4] ), .Y(n323) );
  MUX2X1 U431 ( .B(n324), .A(n92), .S(n65), .Y(n1339) );
  INVX1 U432 ( .A(\memory[7][5] ), .Y(n324) );
  MUX2X1 U433 ( .B(n325), .A(n91), .S(n65), .Y(n1340) );
  INVX1 U434 ( .A(\memory[7][6] ), .Y(n325) );
  MUX2X1 U435 ( .B(n326), .A(n90), .S(n65), .Y(n1341) );
  INVX1 U436 ( .A(\memory[7][7] ), .Y(n326) );
  MUX2X1 U437 ( .B(n88), .A(n327), .S(n328), .Y(n1342) );
  INVX1 U438 ( .A(\opcode[6][0] ), .Y(n327) );
  MUX2X1 U439 ( .B(n86), .A(n329), .S(n328), .Y(n1343) );
  AOI21X1 U440 ( .A(n133), .B(n318), .C(n66), .Y(n328) );
  INVX1 U441 ( .A(n157), .Y(n318) );
  INVX1 U442 ( .A(\opcode[6][1] ), .Y(n329) );
  MUX2X1 U443 ( .B(n330), .A(n97), .S(n66), .Y(n1344) );
  INVX1 U444 ( .A(\memory[6][0] ), .Y(n330) );
  MUX2X1 U445 ( .B(n331), .A(n96), .S(n66), .Y(n1345) );
  INVX1 U446 ( .A(\memory[6][1] ), .Y(n331) );
  MUX2X1 U447 ( .B(n332), .A(n95), .S(n66), .Y(n1346) );
  INVX1 U448 ( .A(\memory[6][2] ), .Y(n332) );
  MUX2X1 U449 ( .B(n333), .A(n94), .S(n66), .Y(n1347) );
  INVX1 U450 ( .A(\memory[6][3] ), .Y(n333) );
  MUX2X1 U451 ( .B(n334), .A(n93), .S(n66), .Y(n1348) );
  INVX1 U452 ( .A(\memory[6][4] ), .Y(n334) );
  MUX2X1 U453 ( .B(n335), .A(n92), .S(n66), .Y(n1349) );
  INVX1 U454 ( .A(\memory[6][5] ), .Y(n335) );
  MUX2X1 U455 ( .B(n336), .A(n91), .S(n66), .Y(n1350) );
  INVX1 U456 ( .A(\memory[6][6] ), .Y(n336) );
  MUX2X1 U457 ( .B(n337), .A(n90), .S(n66), .Y(n1351) );
  INVX1 U458 ( .A(\memory[6][7] ), .Y(n337) );
  MUX2X1 U459 ( .B(n106), .A(n338), .S(n339), .Y(n1352) );
  INVX1 U460 ( .A(\opcode[5][0] ), .Y(n338) );
  MUX2X1 U461 ( .B(n86), .A(n340), .S(n339), .Y(n1353) );
  AOI21X1 U462 ( .A(n138), .B(n165), .C(n67), .Y(n339) );
  INVX1 U463 ( .A(\opcode[5][1] ), .Y(n340) );
  MUX2X1 U464 ( .B(n341), .A(n97), .S(n67), .Y(n1354) );
  INVX1 U465 ( .A(\memory[5][0] ), .Y(n341) );
  MUX2X1 U466 ( .B(n342), .A(n96), .S(n67), .Y(n1355) );
  INVX1 U467 ( .A(\memory[5][1] ), .Y(n342) );
  MUX2X1 U468 ( .B(n343), .A(n95), .S(n67), .Y(n1356) );
  INVX1 U469 ( .A(\memory[5][2] ), .Y(n343) );
  MUX2X1 U470 ( .B(n344), .A(n94), .S(n67), .Y(n1357) );
  INVX1 U471 ( .A(\memory[5][3] ), .Y(n344) );
  MUX2X1 U472 ( .B(n345), .A(n93), .S(n67), .Y(n1358) );
  INVX1 U473 ( .A(\memory[5][4] ), .Y(n345) );
  MUX2X1 U474 ( .B(n346), .A(n92), .S(n67), .Y(n1359) );
  INVX1 U475 ( .A(\memory[5][5] ), .Y(n346) );
  MUX2X1 U476 ( .B(n347), .A(n91), .S(n67), .Y(n1360) );
  INVX1 U477 ( .A(\memory[5][6] ), .Y(n347) );
  MUX2X1 U478 ( .B(n348), .A(n90), .S(n67), .Y(n1361) );
  INVX1 U479 ( .A(\memory[5][7] ), .Y(n348) );
  MUX2X1 U480 ( .B(n88), .A(n349), .S(n350), .Y(n1362) );
  INVX1 U481 ( .A(\opcode[4][0] ), .Y(n349) );
  MUX2X1 U482 ( .B(n86), .A(n351), .S(n350), .Y(n1363) );
  AOI21X1 U483 ( .A(n143), .B(n165), .C(n68), .Y(n350) );
  INVX1 U484 ( .A(\opcode[4][1] ), .Y(n351) );
  MUX2X1 U485 ( .B(n352), .A(n97), .S(n68), .Y(n1364) );
  INVX1 U486 ( .A(\memory[4][0] ), .Y(n352) );
  MUX2X1 U487 ( .B(n353), .A(n96), .S(n68), .Y(n1365) );
  INVX1 U488 ( .A(\memory[4][1] ), .Y(n353) );
  MUX2X1 U489 ( .B(n354), .A(n95), .S(n68), .Y(n1366) );
  INVX1 U490 ( .A(\memory[4][2] ), .Y(n354) );
  MUX2X1 U491 ( .B(n355), .A(n94), .S(n68), .Y(n1367) );
  INVX1 U492 ( .A(\memory[4][3] ), .Y(n355) );
  MUX2X1 U493 ( .B(n356), .A(n93), .S(n68), .Y(n1368) );
  INVX1 U494 ( .A(\memory[4][4] ), .Y(n356) );
  MUX2X1 U495 ( .B(n357), .A(n92), .S(n68), .Y(n1369) );
  INVX1 U496 ( .A(\memory[4][5] ), .Y(n357) );
  MUX2X1 U497 ( .B(n358), .A(n91), .S(n68), .Y(n1370) );
  INVX1 U498 ( .A(\memory[4][6] ), .Y(n358) );
  MUX2X1 U499 ( .B(n359), .A(n90), .S(n68), .Y(n1371) );
  NAND3X1 U500 ( .A(n47), .B(n82), .C(n360), .Y(n286) );
  INVX1 U501 ( .A(\memory[4][7] ), .Y(n359) );
  OAI21X1 U502 ( .A(n361), .B(n362), .C(n363), .Y(n1373) );
  AOI22X1 U503 ( .A(N51), .B(n53), .C(N46), .D(n2), .Y(n363) );
  OAI21X1 U504 ( .A(n361), .B(n82), .C(n364), .Y(n1374) );
  AOI22X1 U505 ( .A(N50), .B(n53), .C(N45), .D(n2), .Y(n364) );
  OAI21X1 U506 ( .A(n361), .B(n80), .C(n365), .Y(n1375) );
  AOI22X1 U507 ( .A(n80), .B(n53), .C(n80), .D(n2), .Y(n365) );
  OAI21X1 U508 ( .A(n361), .B(n366), .C(n367), .Y(n1376) );
  AOI22X1 U509 ( .A(N48), .B(n53), .C(N43), .D(n2), .Y(n367) );
  OAI21X1 U510 ( .A(n361), .B(n75), .C(n368), .Y(n1377) );
  AOI22X1 U511 ( .A(N49), .B(n53), .C(N44), .D(n2), .Y(n368) );
  MUX2X1 U512 ( .B(n90), .A(n369), .S(n21), .Y(n1202) );
  MUX2X1 U513 ( .B(n91), .A(n370), .S(n21), .Y(n1203) );
  MUX2X1 U514 ( .B(n92), .A(n371), .S(n21), .Y(n1204) );
  MUX2X1 U515 ( .B(n93), .A(n372), .S(n21), .Y(n1205) );
  MUX2X1 U516 ( .B(n94), .A(n373), .S(n21), .Y(n1206) );
  MUX2X1 U517 ( .B(n95), .A(n374), .S(n21), .Y(n1207) );
  MUX2X1 U518 ( .B(n96), .A(n375), .S(n21), .Y(n1208) );
  MUX2X1 U519 ( .B(n97), .A(n376), .S(n21), .Y(n1209) );
  MUX2X1 U520 ( .B(n90), .A(n377), .S(n16), .Y(n1210) );
  MUX2X1 U521 ( .B(n91), .A(n378), .S(n16), .Y(n1211) );
  MUX2X1 U522 ( .B(n92), .A(n379), .S(n16), .Y(n1212) );
  MUX2X1 U523 ( .B(n93), .A(n380), .S(n16), .Y(n1213) );
  MUX2X1 U524 ( .B(n94), .A(n381), .S(n16), .Y(n1214) );
  MUX2X1 U525 ( .B(n95), .A(n382), .S(n16), .Y(n1215) );
  MUX2X1 U526 ( .B(n96), .A(n383), .S(n16), .Y(n1216) );
  MUX2X1 U527 ( .B(n97), .A(n384), .S(n16), .Y(n1217) );
  MUX2X1 U528 ( .B(n90), .A(n385), .S(n19), .Y(n1218) );
  MUX2X1 U529 ( .B(n91), .A(n386), .S(n19), .Y(n1219) );
  MUX2X1 U530 ( .B(n92), .A(n387), .S(n19), .Y(n1220) );
  MUX2X1 U531 ( .B(n93), .A(n388), .S(n19), .Y(n1221) );
  MUX2X1 U532 ( .B(n94), .A(n389), .S(n19), .Y(n1222) );
  MUX2X1 U533 ( .B(n95), .A(n390), .S(n19), .Y(n1223) );
  MUX2X1 U534 ( .B(n96), .A(n391), .S(n19), .Y(n1224) );
  MUX2X1 U535 ( .B(n97), .A(n392), .S(n19), .Y(n1225) );
  MUX2X1 U536 ( .B(n393), .A(n90), .S(n394), .Y(n1226) );
  MUX2X1 U537 ( .B(n395), .A(n91), .S(n394), .Y(n1227) );
  MUX2X1 U538 ( .B(n396), .A(n92), .S(n394), .Y(n1228) );
  MUX2X1 U539 ( .B(n397), .A(n93), .S(n394), .Y(n1229) );
  MUX2X1 U540 ( .B(n398), .A(n94), .S(n394), .Y(n1230) );
  MUX2X1 U541 ( .B(n399), .A(n95), .S(n394), .Y(n1231) );
  MUX2X1 U542 ( .B(n400), .A(n96), .S(n394), .Y(n1232) );
  MUX2X1 U543 ( .B(n401), .A(n97), .S(n394), .Y(n1233) );
  MUX2X1 U544 ( .B(n402), .A(n90), .S(n69), .Y(n1234) );
  MUX2X1 U545 ( .B(n403), .A(n91), .S(n69), .Y(n1235) );
  MUX2X1 U546 ( .B(n404), .A(n92), .S(n69), .Y(n1236) );
  MUX2X1 U547 ( .B(n405), .A(n93), .S(n69), .Y(n1237) );
  MUX2X1 U548 ( .B(n406), .A(n94), .S(n69), .Y(n1238) );
  MUX2X1 U549 ( .B(n407), .A(n95), .S(n69), .Y(n1239) );
  MUX2X1 U550 ( .B(n408), .A(n96), .S(n69), .Y(n1240) );
  MUX2X1 U551 ( .B(n409), .A(n97), .S(n69), .Y(n1241) );
  MUX2X1 U552 ( .B(n410), .A(n90), .S(n70), .Y(n1242) );
  MUX2X1 U553 ( .B(n411), .A(n91), .S(n70), .Y(n1243) );
  MUX2X1 U554 ( .B(n412), .A(n92), .S(n70), .Y(n1244) );
  MUX2X1 U555 ( .B(n413), .A(n93), .S(n70), .Y(n1245) );
  MUX2X1 U556 ( .B(n414), .A(n94), .S(n70), .Y(n1246) );
  MUX2X1 U557 ( .B(n415), .A(n95), .S(n70), .Y(n1247) );
  MUX2X1 U558 ( .B(n416), .A(n96), .S(n70), .Y(n1248) );
  MUX2X1 U559 ( .B(n417), .A(n97), .S(n70), .Y(n1249) );
  MUX2X1 U560 ( .B(n418), .A(n90), .S(n71), .Y(n1250) );
  MUX2X1 U561 ( .B(n419), .A(n91), .S(n71), .Y(n1251) );
  MUX2X1 U562 ( .B(n420), .A(n92), .S(n71), .Y(n1252) );
  MUX2X1 U563 ( .B(n421), .A(n93), .S(n71), .Y(n1253) );
  MUX2X1 U564 ( .B(n422), .A(n94), .S(n71), .Y(n1254) );
  MUX2X1 U565 ( .B(n423), .A(n95), .S(n71), .Y(n1255) );
  MUX2X1 U566 ( .B(n424), .A(n96), .S(n71), .Y(n1256) );
  MUX2X1 U567 ( .B(n425), .A(n97), .S(n71), .Y(n1257) );
  MUX2X1 U568 ( .B(n426), .A(n90), .S(n72), .Y(n1258) );
  MUX2X1 U569 ( .B(n427), .A(n91), .S(n72), .Y(n1259) );
  MUX2X1 U570 ( .B(n428), .A(n92), .S(n72), .Y(n1260) );
  MUX2X1 U571 ( .B(n429), .A(n93), .S(n72), .Y(n1261) );
  MUX2X1 U572 ( .B(n430), .A(n94), .S(n72), .Y(n1262) );
  MUX2X1 U573 ( .B(n431), .A(n95), .S(n72), .Y(n1263) );
  MUX2X1 U574 ( .B(n432), .A(n96), .S(n72), .Y(n1264) );
  MUX2X1 U575 ( .B(n433), .A(n97), .S(n72), .Y(n1265) );
  INVX1 U576 ( .A(n434), .Y(n1266) );
  MUX2X1 U577 ( .B(\memory[28][7] ), .A(RCV_DATA[7]), .S(n435), .Y(n434) );
  INVX1 U578 ( .A(n436), .Y(n1267) );
  MUX2X1 U579 ( .B(\memory[28][6] ), .A(RCV_DATA[6]), .S(n435), .Y(n436) );
  INVX1 U580 ( .A(n437), .Y(n1268) );
  MUX2X1 U581 ( .B(\memory[28][5] ), .A(RCV_DATA[5]), .S(n435), .Y(n437) );
  INVX1 U582 ( .A(n438), .Y(n1269) );
  MUX2X1 U583 ( .B(\memory[28][4] ), .A(RCV_DATA[4]), .S(n435), .Y(n438) );
  INVX1 U584 ( .A(n439), .Y(n1270) );
  MUX2X1 U585 ( .B(\memory[28][3] ), .A(RCV_DATA[3]), .S(n435), .Y(n439) );
  INVX1 U586 ( .A(n440), .Y(n1271) );
  MUX2X1 U587 ( .B(\memory[28][2] ), .A(RCV_DATA[2]), .S(n435), .Y(n440) );
  INVX1 U588 ( .A(n441), .Y(n1272) );
  MUX2X1 U589 ( .B(\memory[28][1] ), .A(RCV_DATA[1]), .S(n435), .Y(n441) );
  INVX1 U590 ( .A(n442), .Y(n1273) );
  MUX2X1 U591 ( .B(\memory[28][0] ), .A(RCV_DATA[0]), .S(n435), .Y(n442) );
  INVX1 U592 ( .A(n443), .Y(n1274) );
  MUX2X1 U593 ( .B(\memory[29][7] ), .A(RCV_DATA[7]), .S(n73), .Y(n443) );
  INVX1 U594 ( .A(n444), .Y(n1275) );
  MUX2X1 U595 ( .B(\memory[29][6] ), .A(RCV_DATA[6]), .S(n73), .Y(n444) );
  INVX1 U596 ( .A(n445), .Y(n1276) );
  MUX2X1 U597 ( .B(\memory[29][5] ), .A(RCV_DATA[5]), .S(n73), .Y(n445) );
  INVX1 U598 ( .A(n446), .Y(n1277) );
  MUX2X1 U599 ( .B(\memory[29][4] ), .A(RCV_DATA[4]), .S(n73), .Y(n446) );
  INVX1 U600 ( .A(n447), .Y(n1278) );
  MUX2X1 U601 ( .B(\memory[29][3] ), .A(RCV_DATA[3]), .S(n73), .Y(n447) );
  INVX1 U602 ( .A(n448), .Y(n1279) );
  MUX2X1 U603 ( .B(\memory[29][2] ), .A(RCV_DATA[2]), .S(n73), .Y(n448) );
  INVX1 U604 ( .A(n449), .Y(n1280) );
  MUX2X1 U605 ( .B(\memory[29][1] ), .A(RCV_DATA[1]), .S(n73), .Y(n449) );
  INVX1 U606 ( .A(n450), .Y(n1281) );
  MUX2X1 U607 ( .B(\memory[29][0] ), .A(RCV_DATA[0]), .S(n73), .Y(n450) );
  INVX1 U608 ( .A(n451), .Y(n1282) );
  MUX2X1 U609 ( .B(\memory[30][7] ), .A(RCV_DATA[7]), .S(n74), .Y(n451) );
  INVX1 U610 ( .A(n453), .Y(n1283) );
  MUX2X1 U611 ( .B(\memory[30][6] ), .A(RCV_DATA[6]), .S(n74), .Y(n453) );
  INVX1 U612 ( .A(n454), .Y(n1284) );
  MUX2X1 U613 ( .B(\memory[30][5] ), .A(RCV_DATA[5]), .S(n74), .Y(n454) );
  INVX1 U614 ( .A(n455), .Y(n1285) );
  MUX2X1 U615 ( .B(\memory[30][4] ), .A(RCV_DATA[4]), .S(n74), .Y(n455) );
  INVX1 U616 ( .A(n456), .Y(n1286) );
  MUX2X1 U617 ( .B(\memory[30][3] ), .A(RCV_DATA[3]), .S(n74), .Y(n456) );
  INVX1 U618 ( .A(n457), .Y(n1287) );
  MUX2X1 U619 ( .B(\memory[30][2] ), .A(RCV_DATA[2]), .S(n74), .Y(n457) );
  INVX1 U620 ( .A(n458), .Y(n1288) );
  MUX2X1 U621 ( .B(\memory[30][1] ), .A(RCV_DATA[1]), .S(n74), .Y(n458) );
  INVX1 U622 ( .A(n459), .Y(n1289) );
  MUX2X1 U623 ( .B(\memory[30][0] ), .A(RCV_DATA[0]), .S(n74), .Y(n459) );
  INVX1 U624 ( .A(n460), .Y(n1290) );
  MUX2X1 U625 ( .B(\memory[31][7] ), .A(RCV_DATA[7]), .S(n461), .Y(n460) );
  INVX1 U626 ( .A(n462), .Y(n1291) );
  MUX2X1 U627 ( .B(\memory[31][6] ), .A(RCV_DATA[6]), .S(n461), .Y(n462) );
  INVX1 U628 ( .A(n463), .Y(n1292) );
  MUX2X1 U629 ( .B(\memory[31][5] ), .A(RCV_DATA[5]), .S(n461), .Y(n463) );
  INVX1 U630 ( .A(n464), .Y(n1293) );
  MUX2X1 U631 ( .B(\memory[31][4] ), .A(RCV_DATA[4]), .S(n461), .Y(n464) );
  INVX1 U632 ( .A(n465), .Y(n1294) );
  MUX2X1 U633 ( .B(\memory[31][3] ), .A(RCV_DATA[3]), .S(n461), .Y(n465) );
  INVX1 U634 ( .A(n466), .Y(n1295) );
  MUX2X1 U635 ( .B(\memory[31][2] ), .A(RCV_DATA[2]), .S(n461), .Y(n466) );
  INVX1 U636 ( .A(n467), .Y(n1296) );
  MUX2X1 U637 ( .B(\memory[31][1] ), .A(RCV_DATA[1]), .S(n461), .Y(n467) );
  INVX1 U638 ( .A(n468), .Y(n1297) );
  MUX2X1 U639 ( .B(\memory[31][0] ), .A(RCV_DATA[0]), .S(n461), .Y(n468) );
  MUX2X1 U640 ( .B(n469), .A(n87), .S(n470), .Y(n1298) );
  MUX2X1 U641 ( .B(n471), .A(n88), .S(n470), .Y(n1299) );
  OAI21X1 U642 ( .A(n193), .B(n157), .C(n21), .Y(n470) );
  MUX2X1 U643 ( .B(n472), .A(n87), .S(n473), .Y(n1300) );
  MUX2X1 U644 ( .B(n474), .A(n88), .S(n473), .Y(n1301) );
  OAI21X1 U645 ( .A(n184), .B(n157), .C(n16), .Y(n473) );
  MUX2X1 U646 ( .B(n475), .A(n87), .S(n476), .Y(n1302) );
  MUX2X1 U647 ( .B(n477), .A(n88), .S(n476), .Y(n1303) );
  OAI21X1 U648 ( .A(n244), .B(n157), .C(n19), .Y(n476) );
  NAND2X1 U649 ( .A(n478), .B(n2), .Y(n157) );
  MUX2X1 U650 ( .B(n86), .A(n479), .S(n480), .Y(n1304) );
  MUX2X1 U651 ( .B(n88), .A(n481), .S(n480), .Y(n1305) );
  NAND3X1 U652 ( .A(n478), .B(n361), .C(n482), .Y(n480) );
  MUX2X1 U653 ( .B(n184), .A(n235), .S(n483), .Y(n482) );
  AND2X1 U654 ( .A(n360), .B(n83), .Y(n478) );
  MUX2X1 U655 ( .B(n86), .A(n484), .S(n485), .Y(n1306) );
  MUX2X1 U656 ( .B(n88), .A(n486), .S(n485), .Y(n1307) );
  AOI21X1 U657 ( .A(n123), .B(n139), .C(n69), .Y(n485) );
  INVX1 U658 ( .A(n193), .Y(n123) );
  MUX2X1 U659 ( .B(n86), .A(n487), .S(n488), .Y(n1308) );
  MUX2X1 U660 ( .B(n88), .A(n489), .S(n488), .Y(n1309) );
  AOI21X1 U661 ( .A(n118), .B(n139), .C(n70), .Y(n488) );
  INVX1 U662 ( .A(n184), .Y(n118) );
  MUX2X1 U663 ( .B(n86), .A(n490), .S(n491), .Y(n1310) );
  MUX2X1 U664 ( .B(n88), .A(n492), .S(n491), .Y(n1311) );
  AOI21X1 U665 ( .A(n113), .B(n139), .C(n71), .Y(n491) );
  NAND3X1 U666 ( .A(n80), .B(n75), .C(n79), .Y(n193) );
  INVX1 U667 ( .A(n244), .Y(n113) );
  MUX2X1 U668 ( .B(n86), .A(n493), .S(n494), .Y(n1312) );
  MUX2X1 U669 ( .B(n88), .A(n495), .S(n494), .Y(n1313) );
  AOI21X1 U670 ( .A(n108), .B(n139), .C(n72), .Y(n494) );
  NAND3X1 U671 ( .A(n81), .B(n75), .C(n79), .Y(n184) );
  NAND3X1 U672 ( .A(n496), .B(n82), .C(n2), .Y(n148) );
  INVX1 U673 ( .A(n235), .Y(n108) );
  MUX2X1 U674 ( .B(n86), .A(n497), .S(n498), .Y(n1314) );
  INVX1 U675 ( .A(\opcode[28][1] ), .Y(n497) );
  MUX2X1 U676 ( .B(n88), .A(n499), .S(n498), .Y(n1315) );
  AOI21X1 U677 ( .A(n109), .B(n143), .C(n435), .Y(n498) );
  NAND3X1 U678 ( .A(n80), .B(n366), .C(n76), .Y(n244) );
  INVX1 U679 ( .A(n161), .Y(n143) );
  INVX1 U680 ( .A(\opcode[28][0] ), .Y(n499) );
  MUX2X1 U681 ( .B(n86), .A(n500), .S(n501), .Y(n1316) );
  INVX1 U682 ( .A(\opcode[29][1] ), .Y(n500) );
  MUX2X1 U683 ( .B(n88), .A(n502), .S(n501), .Y(n1317) );
  AOI21X1 U684 ( .A(n109), .B(n138), .C(n73), .Y(n501) );
  NAND3X1 U685 ( .A(n81), .B(n366), .C(n76), .Y(n235) );
  INVX1 U686 ( .A(n156), .Y(n138) );
  NAND3X1 U687 ( .A(n2), .B(n496), .C(n83), .Y(n503) );
  INVX1 U688 ( .A(\opcode[29][0] ), .Y(n502) );
  MUX2X1 U689 ( .B(n86), .A(n504), .S(n505), .Y(n1318) );
  INVX1 U690 ( .A(\opcode[30][1] ), .Y(n504) );
  MUX2X1 U691 ( .B(n88), .A(n506), .S(n505), .Y(n1319) );
  AOI21X1 U692 ( .A(n133), .B(n165), .C(n74), .Y(n505) );
  NOR2X1 U693 ( .A(n161), .B(n43), .Y(n452) );
  NAND3X1 U694 ( .A(n76), .B(n80), .C(n79), .Y(n161) );
  INVX1 U695 ( .A(n152), .Y(n133) );
  NAND3X1 U696 ( .A(n366), .B(n75), .C(n80), .Y(n152) );
  INVX1 U697 ( .A(\opcode[30][0] ), .Y(n506) );
  MUX2X1 U698 ( .B(n87), .A(n507), .S(n508), .Y(n1320) );
  INVX1 U699 ( .A(\opcode[31][1] ), .Y(n507) );
  MUX2X1 U700 ( .B(n106), .A(n509), .S(n508), .Y(n1321) );
  AOI21X1 U701 ( .A(n128), .B(n165), .C(n461), .Y(n508) );
  NOR2X1 U702 ( .A(n362), .B(RST), .Y(n496) );
  INVX1 U703 ( .A(writeptr[4]), .Y(n362) );
  NAND3X1 U704 ( .A(n76), .B(n81), .C(n79), .Y(n156) );
  NAND3X1 U705 ( .A(n2), .B(n82), .C(n360), .Y(n511) );
  NOR2X1 U706 ( .A(writeptr[4]), .B(RST), .Y(n360) );
  NAND2X1 U707 ( .A(W_ENABLE), .B(n311), .Y(n510) );
  NAND3X1 U708 ( .A(n512), .B(n513), .C(n514), .Y(n311) );
  NOR2X1 U709 ( .A(n515), .B(n516), .Y(n514) );
  XOR2X1 U710 ( .A(readptr[3]), .B(N34), .Y(n515) );
  XOR2X1 U711 ( .A(n517), .B(N32), .Y(n513) );
  NOR2X1 U712 ( .A(n518), .B(n519), .Y(n512) );
  XOR2X1 U713 ( .A(readptr[2]), .B(N33), .Y(n518) );
  INVX1 U714 ( .A(n147), .Y(n128) );
  NAND3X1 U715 ( .A(n366), .B(n75), .C(n81), .Y(n147) );
  INVX1 U716 ( .A(n79), .Y(n366) );
  INVX1 U717 ( .A(\opcode[31][0] ), .Y(n509) );
  INVX1 U718 ( .A(n520), .Y(n1322) );
  MUX2X1 U719 ( .B(n521), .A(DATA[7]), .S(n522), .Y(n520) );
  NAND2X1 U720 ( .A(n523), .B(n524), .Y(n521) );
  NOR2X1 U721 ( .A(n525), .B(n526), .Y(n524) );
  NAND3X1 U722 ( .A(n527), .B(n528), .C(n529), .Y(n526) );
  NOR2X1 U723 ( .A(n530), .B(n531), .Y(n529) );
  OAI22X1 U724 ( .A(n402), .B(n532), .C(n410), .D(n533), .Y(n531) );
  INVX1 U725 ( .A(\memory[17][7] ), .Y(n410) );
  INVX1 U726 ( .A(\memory[16][7] ), .Y(n402) );
  OAI22X1 U727 ( .A(n418), .B(n534), .C(n426), .D(n535), .Y(n530) );
  INVX1 U728 ( .A(\memory[19][7] ), .Y(n426) );
  INVX1 U729 ( .A(\memory[18][7] ), .Y(n418) );
  AOI22X1 U730 ( .A(n536), .B(\memory[23][7] ), .C(n537), .D(\memory[22][7] ), 
        .Y(n528) );
  AOI22X1 U731 ( .A(n538), .B(\memory[21][7] ), .C(n539), .D(\memory[20][7] ), 
        .Y(n527) );
  NAND3X1 U732 ( .A(n540), .B(n541), .C(n542), .Y(n525) );
  NOR2X1 U733 ( .A(n543), .B(n544), .Y(n542) );
  OAI22X1 U734 ( .A(n202), .B(n545), .C(n194), .D(n546), .Y(n544) );
  INVX1 U735 ( .A(\memory[25][7] ), .Y(n194) );
  INVX1 U736 ( .A(\memory[24][7] ), .Y(n202) );
  OAI22X1 U737 ( .A(n185), .B(n547), .C(n175), .D(n548), .Y(n543) );
  INVX1 U738 ( .A(\memory[27][7] ), .Y(n175) );
  INVX1 U739 ( .A(\memory[26][7] ), .Y(n185) );
  AOI22X1 U740 ( .A(n549), .B(\memory[31][7] ), .C(n550), .D(\memory[30][7] ), 
        .Y(n541) );
  AOI22X1 U741 ( .A(n551), .B(\memory[29][7] ), .C(n552), .D(\memory[28][7] ), 
        .Y(n540) );
  NOR2X1 U742 ( .A(n553), .B(n554), .Y(n523) );
  NAND3X1 U743 ( .A(n555), .B(n556), .C(n557), .Y(n554) );
  NOR2X1 U744 ( .A(n558), .B(n559), .Y(n557) );
  OAI22X1 U745 ( .A(n310), .B(n560), .C(n302), .D(n561), .Y(n559) );
  INVX1 U746 ( .A(\memory[2][7] ), .Y(n302) );
  INVX1 U747 ( .A(\memory[3][7] ), .Y(n310) );
  OAI22X1 U748 ( .A(n294), .B(n562), .C(n285), .D(n563), .Y(n558) );
  INVX1 U749 ( .A(\memory[0][7] ), .Y(n285) );
  INVX1 U750 ( .A(\memory[1][7] ), .Y(n294) );
  AOI22X1 U751 ( .A(n564), .B(\memory[4][7] ), .C(n565), .D(\memory[5][7] ), 
        .Y(n556) );
  AOI22X1 U752 ( .A(n566), .B(\memory[6][7] ), .C(n567), .D(\memory[7][7] ), 
        .Y(n555) );
  NAND3X1 U753 ( .A(n568), .B(n569), .C(n570), .Y(n553) );
  NOR2X1 U754 ( .A(n571), .B(n572), .Y(n570) );
  OAI22X1 U755 ( .A(n369), .B(n573), .C(n377), .D(n574), .Y(n572) );
  INVX1 U756 ( .A(\memory[9][7] ), .Y(n377) );
  INVX1 U757 ( .A(\memory[8][7] ), .Y(n369) );
  OAI22X1 U758 ( .A(n385), .B(n575), .C(n393), .D(n576), .Y(n571) );
  INVX1 U759 ( .A(\memory[11][7] ), .Y(n393) );
  INVX1 U760 ( .A(\memory[10][7] ), .Y(n385) );
  AOI22X1 U761 ( .A(n577), .B(\memory[15][7] ), .C(n578), .D(\memory[14][7] ), 
        .Y(n569) );
  AOI22X1 U762 ( .A(n579), .B(\memory[13][7] ), .C(n580), .D(\memory[12][7] ), 
        .Y(n568) );
  INVX1 U763 ( .A(n581), .Y(n1323) );
  MUX2X1 U764 ( .B(n582), .A(DATA[6]), .S(n522), .Y(n581) );
  NAND2X1 U765 ( .A(n583), .B(n584), .Y(n582) );
  NOR2X1 U766 ( .A(n585), .B(n586), .Y(n584) );
  NAND3X1 U767 ( .A(n587), .B(n588), .C(n589), .Y(n586) );
  NOR2X1 U768 ( .A(n590), .B(n591), .Y(n589) );
  OAI22X1 U769 ( .A(n403), .B(n532), .C(n411), .D(n533), .Y(n591) );
  INVX1 U770 ( .A(\memory[17][6] ), .Y(n411) );
  INVX1 U771 ( .A(\memory[16][6] ), .Y(n403) );
  OAI22X1 U772 ( .A(n419), .B(n534), .C(n427), .D(n535), .Y(n590) );
  INVX1 U773 ( .A(\memory[19][6] ), .Y(n427) );
  INVX1 U774 ( .A(\memory[18][6] ), .Y(n419) );
  AOI22X1 U775 ( .A(n536), .B(\memory[23][6] ), .C(n537), .D(\memory[22][6] ), 
        .Y(n588) );
  AOI22X1 U776 ( .A(n538), .B(\memory[21][6] ), .C(n539), .D(\memory[20][6] ), 
        .Y(n587) );
  NAND3X1 U777 ( .A(n592), .B(n593), .C(n594), .Y(n585) );
  NOR2X1 U778 ( .A(n595), .B(n596), .Y(n594) );
  OAI22X1 U779 ( .A(n203), .B(n545), .C(n195), .D(n546), .Y(n596) );
  INVX1 U780 ( .A(\memory[25][6] ), .Y(n195) );
  INVX1 U781 ( .A(\memory[24][6] ), .Y(n203) );
  OAI22X1 U782 ( .A(n186), .B(n547), .C(n176), .D(n548), .Y(n595) );
  INVX1 U783 ( .A(\memory[27][6] ), .Y(n176) );
  INVX1 U784 ( .A(\memory[26][6] ), .Y(n186) );
  AOI22X1 U785 ( .A(n549), .B(\memory[31][6] ), .C(n550), .D(\memory[30][6] ), 
        .Y(n593) );
  AOI22X1 U786 ( .A(n551), .B(\memory[29][6] ), .C(n552), .D(\memory[28][6] ), 
        .Y(n592) );
  NOR2X1 U787 ( .A(n597), .B(n598), .Y(n583) );
  NAND3X1 U788 ( .A(n599), .B(n600), .C(n601), .Y(n598) );
  NOR2X1 U789 ( .A(n602), .B(n603), .Y(n601) );
  OAI22X1 U790 ( .A(n309), .B(n560), .C(n301), .D(n561), .Y(n603) );
  INVX1 U791 ( .A(\memory[2][6] ), .Y(n301) );
  INVX1 U792 ( .A(\memory[3][6] ), .Y(n309) );
  OAI22X1 U793 ( .A(n293), .B(n562), .C(n284), .D(n563), .Y(n602) );
  INVX1 U794 ( .A(\memory[0][6] ), .Y(n284) );
  INVX1 U795 ( .A(\memory[1][6] ), .Y(n293) );
  AOI22X1 U796 ( .A(n564), .B(\memory[4][6] ), .C(n565), .D(\memory[5][6] ), 
        .Y(n600) );
  AOI22X1 U797 ( .A(n566), .B(\memory[6][6] ), .C(n567), .D(\memory[7][6] ), 
        .Y(n599) );
  NAND3X1 U798 ( .A(n604), .B(n605), .C(n606), .Y(n597) );
  NOR2X1 U799 ( .A(n607), .B(n608), .Y(n606) );
  OAI22X1 U800 ( .A(n370), .B(n573), .C(n378), .D(n574), .Y(n608) );
  INVX1 U801 ( .A(\memory[9][6] ), .Y(n378) );
  INVX1 U802 ( .A(\memory[8][6] ), .Y(n370) );
  OAI22X1 U803 ( .A(n386), .B(n575), .C(n395), .D(n576), .Y(n607) );
  INVX1 U804 ( .A(\memory[11][6] ), .Y(n395) );
  INVX1 U805 ( .A(\memory[10][6] ), .Y(n386) );
  AOI22X1 U806 ( .A(n577), .B(\memory[15][6] ), .C(n578), .D(\memory[14][6] ), 
        .Y(n605) );
  AOI22X1 U807 ( .A(n579), .B(\memory[13][6] ), .C(n580), .D(\memory[12][6] ), 
        .Y(n604) );
  INVX1 U808 ( .A(n609), .Y(n1324) );
  MUX2X1 U809 ( .B(n610), .A(DATA[5]), .S(n522), .Y(n609) );
  NAND2X1 U810 ( .A(n611), .B(n612), .Y(n610) );
  NOR2X1 U811 ( .A(n613), .B(n614), .Y(n612) );
  NAND3X1 U812 ( .A(n615), .B(n616), .C(n617), .Y(n614) );
  NOR2X1 U813 ( .A(n618), .B(n619), .Y(n617) );
  OAI22X1 U814 ( .A(n404), .B(n532), .C(n412), .D(n533), .Y(n619) );
  INVX1 U815 ( .A(\memory[17][5] ), .Y(n412) );
  INVX1 U816 ( .A(\memory[16][5] ), .Y(n404) );
  OAI22X1 U817 ( .A(n420), .B(n534), .C(n428), .D(n535), .Y(n618) );
  INVX1 U818 ( .A(\memory[19][5] ), .Y(n428) );
  INVX1 U819 ( .A(\memory[18][5] ), .Y(n420) );
  AOI22X1 U820 ( .A(n536), .B(\memory[23][5] ), .C(n537), .D(\memory[22][5] ), 
        .Y(n616) );
  AOI22X1 U821 ( .A(n538), .B(\memory[21][5] ), .C(n539), .D(\memory[20][5] ), 
        .Y(n615) );
  NAND3X1 U822 ( .A(n620), .B(n621), .C(n622), .Y(n613) );
  NOR2X1 U823 ( .A(n623), .B(n624), .Y(n622) );
  OAI22X1 U824 ( .A(n204), .B(n545), .C(n196), .D(n546), .Y(n624) );
  INVX1 U825 ( .A(\memory[25][5] ), .Y(n196) );
  INVX1 U826 ( .A(\memory[24][5] ), .Y(n204) );
  OAI22X1 U827 ( .A(n187), .B(n547), .C(n177), .D(n548), .Y(n623) );
  INVX1 U828 ( .A(\memory[27][5] ), .Y(n177) );
  INVX1 U829 ( .A(\memory[26][5] ), .Y(n187) );
  AOI22X1 U830 ( .A(n549), .B(\memory[31][5] ), .C(n550), .D(\memory[30][5] ), 
        .Y(n621) );
  AOI22X1 U831 ( .A(n551), .B(\memory[29][5] ), .C(n552), .D(\memory[28][5] ), 
        .Y(n620) );
  NOR2X1 U832 ( .A(n625), .B(n626), .Y(n611) );
  NAND3X1 U833 ( .A(n627), .B(n628), .C(n629), .Y(n626) );
  NOR2X1 U834 ( .A(n630), .B(n631), .Y(n629) );
  OAI22X1 U835 ( .A(n308), .B(n560), .C(n300), .D(n561), .Y(n631) );
  INVX1 U836 ( .A(\memory[2][5] ), .Y(n300) );
  INVX1 U837 ( .A(\memory[3][5] ), .Y(n308) );
  OAI22X1 U838 ( .A(n292), .B(n562), .C(n283), .D(n563), .Y(n630) );
  INVX1 U839 ( .A(\memory[0][5] ), .Y(n283) );
  INVX1 U840 ( .A(\memory[1][5] ), .Y(n292) );
  AOI22X1 U841 ( .A(n564), .B(\memory[4][5] ), .C(n565), .D(\memory[5][5] ), 
        .Y(n628) );
  AOI22X1 U842 ( .A(n566), .B(\memory[6][5] ), .C(n567), .D(\memory[7][5] ), 
        .Y(n627) );
  NAND3X1 U843 ( .A(n632), .B(n633), .C(n634), .Y(n625) );
  NOR2X1 U844 ( .A(n635), .B(n636), .Y(n634) );
  OAI22X1 U845 ( .A(n371), .B(n573), .C(n379), .D(n574), .Y(n636) );
  INVX1 U846 ( .A(\memory[9][5] ), .Y(n379) );
  INVX1 U847 ( .A(\memory[8][5] ), .Y(n371) );
  OAI22X1 U848 ( .A(n387), .B(n575), .C(n396), .D(n576), .Y(n635) );
  INVX1 U849 ( .A(\memory[11][5] ), .Y(n396) );
  INVX1 U850 ( .A(\memory[10][5] ), .Y(n387) );
  AOI22X1 U851 ( .A(n577), .B(\memory[15][5] ), .C(n578), .D(\memory[14][5] ), 
        .Y(n633) );
  AOI22X1 U852 ( .A(n579), .B(\memory[13][5] ), .C(n580), .D(\memory[12][5] ), 
        .Y(n632) );
  INVX1 U853 ( .A(n637), .Y(n1325) );
  MUX2X1 U854 ( .B(n638), .A(DATA[4]), .S(n522), .Y(n637) );
  NAND2X1 U855 ( .A(n639), .B(n640), .Y(n638) );
  NOR2X1 U856 ( .A(n641), .B(n642), .Y(n640) );
  NAND3X1 U857 ( .A(n643), .B(n644), .C(n645), .Y(n642) );
  NOR2X1 U858 ( .A(n646), .B(n647), .Y(n645) );
  OAI22X1 U859 ( .A(n405), .B(n532), .C(n413), .D(n533), .Y(n647) );
  INVX1 U860 ( .A(\memory[17][4] ), .Y(n413) );
  INVX1 U861 ( .A(\memory[16][4] ), .Y(n405) );
  OAI22X1 U862 ( .A(n421), .B(n534), .C(n429), .D(n535), .Y(n646) );
  INVX1 U863 ( .A(\memory[19][4] ), .Y(n429) );
  INVX1 U864 ( .A(\memory[18][4] ), .Y(n421) );
  AOI22X1 U865 ( .A(n536), .B(\memory[23][4] ), .C(n537), .D(\memory[22][4] ), 
        .Y(n644) );
  AOI22X1 U866 ( .A(n538), .B(\memory[21][4] ), .C(n539), .D(\memory[20][4] ), 
        .Y(n643) );
  NAND3X1 U867 ( .A(n648), .B(n649), .C(n650), .Y(n641) );
  NOR2X1 U868 ( .A(n651), .B(n652), .Y(n650) );
  OAI22X1 U869 ( .A(n205), .B(n545), .C(n197), .D(n546), .Y(n652) );
  INVX1 U870 ( .A(\memory[25][4] ), .Y(n197) );
  INVX1 U871 ( .A(\memory[24][4] ), .Y(n205) );
  OAI22X1 U872 ( .A(n188), .B(n547), .C(n178), .D(n548), .Y(n651) );
  INVX1 U873 ( .A(\memory[27][4] ), .Y(n178) );
  INVX1 U874 ( .A(\memory[26][4] ), .Y(n188) );
  AOI22X1 U875 ( .A(n549), .B(\memory[31][4] ), .C(n550), .D(\memory[30][4] ), 
        .Y(n649) );
  AOI22X1 U876 ( .A(n551), .B(\memory[29][4] ), .C(n552), .D(\memory[28][4] ), 
        .Y(n648) );
  NOR2X1 U877 ( .A(n653), .B(n654), .Y(n639) );
  NAND3X1 U878 ( .A(n655), .B(n656), .C(n657), .Y(n654) );
  NOR2X1 U879 ( .A(n658), .B(n659), .Y(n657) );
  OAI22X1 U880 ( .A(n307), .B(n560), .C(n299), .D(n561), .Y(n659) );
  INVX1 U881 ( .A(\memory[2][4] ), .Y(n299) );
  INVX1 U882 ( .A(\memory[3][4] ), .Y(n307) );
  OAI22X1 U883 ( .A(n291), .B(n562), .C(n282), .D(n563), .Y(n658) );
  INVX1 U884 ( .A(\memory[0][4] ), .Y(n282) );
  INVX1 U885 ( .A(\memory[1][4] ), .Y(n291) );
  AOI22X1 U886 ( .A(n564), .B(\memory[4][4] ), .C(n565), .D(\memory[5][4] ), 
        .Y(n656) );
  AOI22X1 U887 ( .A(n566), .B(\memory[6][4] ), .C(n567), .D(\memory[7][4] ), 
        .Y(n655) );
  NAND3X1 U888 ( .A(n660), .B(n661), .C(n662), .Y(n653) );
  NOR2X1 U889 ( .A(n663), .B(n664), .Y(n662) );
  OAI22X1 U890 ( .A(n372), .B(n573), .C(n380), .D(n574), .Y(n664) );
  INVX1 U891 ( .A(\memory[9][4] ), .Y(n380) );
  INVX1 U892 ( .A(\memory[8][4] ), .Y(n372) );
  OAI22X1 U893 ( .A(n388), .B(n575), .C(n397), .D(n576), .Y(n663) );
  INVX1 U894 ( .A(\memory[11][4] ), .Y(n397) );
  INVX1 U895 ( .A(\memory[10][4] ), .Y(n388) );
  AOI22X1 U896 ( .A(n577), .B(\memory[15][4] ), .C(n578), .D(\memory[14][4] ), 
        .Y(n661) );
  AOI22X1 U897 ( .A(n579), .B(\memory[13][4] ), .C(n580), .D(\memory[12][4] ), 
        .Y(n660) );
  INVX1 U898 ( .A(n665), .Y(n1326) );
  MUX2X1 U899 ( .B(n666), .A(DATA[3]), .S(n522), .Y(n665) );
  NAND2X1 U900 ( .A(n667), .B(n668), .Y(n666) );
  NOR2X1 U901 ( .A(n669), .B(n670), .Y(n668) );
  NAND3X1 U902 ( .A(n671), .B(n672), .C(n673), .Y(n670) );
  NOR2X1 U903 ( .A(n674), .B(n675), .Y(n673) );
  OAI22X1 U904 ( .A(n406), .B(n532), .C(n414), .D(n533), .Y(n675) );
  INVX1 U905 ( .A(\memory[17][3] ), .Y(n414) );
  INVX1 U906 ( .A(\memory[16][3] ), .Y(n406) );
  OAI22X1 U907 ( .A(n422), .B(n534), .C(n430), .D(n535), .Y(n674) );
  INVX1 U908 ( .A(\memory[19][3] ), .Y(n430) );
  INVX1 U909 ( .A(\memory[18][3] ), .Y(n422) );
  AOI22X1 U910 ( .A(n536), .B(\memory[23][3] ), .C(n537), .D(\memory[22][3] ), 
        .Y(n672) );
  AOI22X1 U911 ( .A(n538), .B(\memory[21][3] ), .C(n539), .D(\memory[20][3] ), 
        .Y(n671) );
  NAND3X1 U912 ( .A(n676), .B(n677), .C(n678), .Y(n669) );
  NOR2X1 U913 ( .A(n679), .B(n680), .Y(n678) );
  OAI22X1 U914 ( .A(n206), .B(n545), .C(n198), .D(n546), .Y(n680) );
  INVX1 U915 ( .A(\memory[25][3] ), .Y(n198) );
  INVX1 U916 ( .A(\memory[24][3] ), .Y(n206) );
  OAI22X1 U917 ( .A(n189), .B(n547), .C(n179), .D(n548), .Y(n679) );
  INVX1 U918 ( .A(\memory[27][3] ), .Y(n179) );
  INVX1 U919 ( .A(\memory[26][3] ), .Y(n189) );
  AOI22X1 U920 ( .A(n549), .B(\memory[31][3] ), .C(n550), .D(\memory[30][3] ), 
        .Y(n677) );
  AOI22X1 U921 ( .A(n551), .B(\memory[29][3] ), .C(n552), .D(\memory[28][3] ), 
        .Y(n676) );
  NOR2X1 U922 ( .A(n681), .B(n682), .Y(n667) );
  NAND3X1 U923 ( .A(n683), .B(n684), .C(n685), .Y(n682) );
  NOR2X1 U924 ( .A(n686), .B(n687), .Y(n685) );
  OAI22X1 U925 ( .A(n306), .B(n560), .C(n298), .D(n561), .Y(n687) );
  INVX1 U926 ( .A(\memory[2][3] ), .Y(n298) );
  INVX1 U927 ( .A(\memory[3][3] ), .Y(n306) );
  OAI22X1 U928 ( .A(n290), .B(n562), .C(n281), .D(n563), .Y(n686) );
  INVX1 U929 ( .A(\memory[0][3] ), .Y(n281) );
  INVX1 U930 ( .A(\memory[1][3] ), .Y(n290) );
  AOI22X1 U931 ( .A(n564), .B(\memory[4][3] ), .C(n565), .D(\memory[5][3] ), 
        .Y(n684) );
  AOI22X1 U932 ( .A(n566), .B(\memory[6][3] ), .C(n567), .D(\memory[7][3] ), 
        .Y(n683) );
  NAND3X1 U933 ( .A(n688), .B(n689), .C(n690), .Y(n681) );
  NOR2X1 U934 ( .A(n691), .B(n692), .Y(n690) );
  OAI22X1 U935 ( .A(n373), .B(n573), .C(n381), .D(n574), .Y(n692) );
  INVX1 U936 ( .A(\memory[9][3] ), .Y(n381) );
  INVX1 U937 ( .A(\memory[8][3] ), .Y(n373) );
  OAI22X1 U938 ( .A(n389), .B(n575), .C(n398), .D(n576), .Y(n691) );
  INVX1 U939 ( .A(\memory[11][3] ), .Y(n398) );
  INVX1 U940 ( .A(\memory[10][3] ), .Y(n389) );
  AOI22X1 U941 ( .A(n577), .B(\memory[15][3] ), .C(n578), .D(\memory[14][3] ), 
        .Y(n689) );
  AOI22X1 U942 ( .A(n579), .B(\memory[13][3] ), .C(n580), .D(\memory[12][3] ), 
        .Y(n688) );
  INVX1 U943 ( .A(n693), .Y(n1327) );
  MUX2X1 U944 ( .B(n694), .A(DATA[2]), .S(n522), .Y(n693) );
  NAND2X1 U945 ( .A(n695), .B(n696), .Y(n694) );
  NOR2X1 U946 ( .A(n697), .B(n698), .Y(n696) );
  NAND3X1 U947 ( .A(n699), .B(n700), .C(n701), .Y(n698) );
  NOR2X1 U948 ( .A(n702), .B(n703), .Y(n701) );
  OAI22X1 U949 ( .A(n407), .B(n532), .C(n415), .D(n533), .Y(n703) );
  INVX1 U950 ( .A(\memory[17][2] ), .Y(n415) );
  INVX1 U951 ( .A(\memory[16][2] ), .Y(n407) );
  OAI22X1 U952 ( .A(n423), .B(n534), .C(n431), .D(n535), .Y(n702) );
  INVX1 U953 ( .A(\memory[19][2] ), .Y(n431) );
  INVX1 U954 ( .A(\memory[18][2] ), .Y(n423) );
  AOI22X1 U955 ( .A(n536), .B(\memory[23][2] ), .C(n537), .D(\memory[22][2] ), 
        .Y(n700) );
  AOI22X1 U956 ( .A(n538), .B(\memory[21][2] ), .C(n539), .D(\memory[20][2] ), 
        .Y(n699) );
  NAND3X1 U957 ( .A(n704), .B(n705), .C(n706), .Y(n697) );
  NOR2X1 U958 ( .A(n707), .B(n708), .Y(n706) );
  OAI22X1 U959 ( .A(n207), .B(n545), .C(n199), .D(n546), .Y(n708) );
  INVX1 U960 ( .A(\memory[25][2] ), .Y(n199) );
  INVX1 U961 ( .A(\memory[24][2] ), .Y(n207) );
  OAI22X1 U962 ( .A(n190), .B(n547), .C(n180), .D(n548), .Y(n707) );
  INVX1 U963 ( .A(\memory[27][2] ), .Y(n180) );
  INVX1 U964 ( .A(\memory[26][2] ), .Y(n190) );
  AOI22X1 U965 ( .A(n549), .B(\memory[31][2] ), .C(n550), .D(\memory[30][2] ), 
        .Y(n705) );
  AOI22X1 U966 ( .A(n551), .B(\memory[29][2] ), .C(n552), .D(\memory[28][2] ), 
        .Y(n704) );
  NOR2X1 U967 ( .A(n709), .B(n710), .Y(n695) );
  NAND3X1 U968 ( .A(n711), .B(n712), .C(n713), .Y(n710) );
  NOR2X1 U969 ( .A(n714), .B(n715), .Y(n713) );
  OAI22X1 U970 ( .A(n305), .B(n560), .C(n297), .D(n561), .Y(n715) );
  INVX1 U971 ( .A(\memory[2][2] ), .Y(n297) );
  INVX1 U972 ( .A(\memory[3][2] ), .Y(n305) );
  OAI22X1 U973 ( .A(n289), .B(n562), .C(n280), .D(n563), .Y(n714) );
  INVX1 U974 ( .A(\memory[0][2] ), .Y(n280) );
  INVX1 U975 ( .A(\memory[1][2] ), .Y(n289) );
  AOI22X1 U976 ( .A(n564), .B(\memory[4][2] ), .C(n565), .D(\memory[5][2] ), 
        .Y(n712) );
  AOI22X1 U977 ( .A(n566), .B(\memory[6][2] ), .C(n567), .D(\memory[7][2] ), 
        .Y(n711) );
  NAND3X1 U978 ( .A(n716), .B(n717), .C(n718), .Y(n709) );
  NOR2X1 U979 ( .A(n719), .B(n720), .Y(n718) );
  OAI22X1 U980 ( .A(n374), .B(n573), .C(n382), .D(n574), .Y(n720) );
  INVX1 U981 ( .A(\memory[9][2] ), .Y(n382) );
  INVX1 U982 ( .A(\memory[8][2] ), .Y(n374) );
  OAI22X1 U983 ( .A(n390), .B(n575), .C(n399), .D(n576), .Y(n719) );
  INVX1 U984 ( .A(\memory[11][2] ), .Y(n399) );
  INVX1 U985 ( .A(\memory[10][2] ), .Y(n390) );
  AOI22X1 U986 ( .A(n577), .B(\memory[15][2] ), .C(n578), .D(\memory[14][2] ), 
        .Y(n717) );
  AOI22X1 U987 ( .A(n579), .B(\memory[13][2] ), .C(n580), .D(\memory[12][2] ), 
        .Y(n716) );
  INVX1 U988 ( .A(n721), .Y(n1328) );
  MUX2X1 U989 ( .B(n722), .A(DATA[1]), .S(n522), .Y(n721) );
  NAND2X1 U990 ( .A(n723), .B(n724), .Y(n722) );
  NOR2X1 U991 ( .A(n725), .B(n726), .Y(n724) );
  NAND3X1 U992 ( .A(n727), .B(n728), .C(n729), .Y(n726) );
  NOR2X1 U993 ( .A(n730), .B(n731), .Y(n729) );
  OAI22X1 U994 ( .A(n408), .B(n532), .C(n416), .D(n533), .Y(n731) );
  INVX1 U995 ( .A(\memory[17][1] ), .Y(n416) );
  INVX1 U996 ( .A(\memory[16][1] ), .Y(n408) );
  OAI22X1 U997 ( .A(n424), .B(n534), .C(n432), .D(n535), .Y(n730) );
  INVX1 U998 ( .A(\memory[19][1] ), .Y(n432) );
  INVX1 U999 ( .A(\memory[18][1] ), .Y(n424) );
  AOI22X1 U1000 ( .A(n536), .B(\memory[23][1] ), .C(n537), .D(\memory[22][1] ), 
        .Y(n728) );
  AOI22X1 U1001 ( .A(n538), .B(\memory[21][1] ), .C(n539), .D(\memory[20][1] ), 
        .Y(n727) );
  NAND3X1 U1002 ( .A(n732), .B(n733), .C(n734), .Y(n725) );
  NOR2X1 U1003 ( .A(n735), .B(n736), .Y(n734) );
  OAI22X1 U1004 ( .A(n208), .B(n545), .C(n200), .D(n546), .Y(n736) );
  INVX1 U1005 ( .A(\memory[25][1] ), .Y(n200) );
  INVX1 U1006 ( .A(\memory[24][1] ), .Y(n208) );
  OAI22X1 U1007 ( .A(n191), .B(n547), .C(n181), .D(n548), .Y(n735) );
  INVX1 U1008 ( .A(\memory[27][1] ), .Y(n181) );
  INVX1 U1009 ( .A(\memory[26][1] ), .Y(n191) );
  AOI22X1 U1010 ( .A(n549), .B(\memory[31][1] ), .C(n550), .D(\memory[30][1] ), 
        .Y(n733) );
  AOI22X1 U1011 ( .A(n551), .B(\memory[29][1] ), .C(n552), .D(\memory[28][1] ), 
        .Y(n732) );
  NOR2X1 U1012 ( .A(n737), .B(n738), .Y(n723) );
  NAND3X1 U1013 ( .A(n739), .B(n740), .C(n741), .Y(n738) );
  NOR2X1 U1014 ( .A(n742), .B(n743), .Y(n741) );
  OAI22X1 U1015 ( .A(n304), .B(n560), .C(n296), .D(n561), .Y(n743) );
  INVX1 U1016 ( .A(\memory[2][1] ), .Y(n296) );
  INVX1 U1017 ( .A(\memory[3][1] ), .Y(n304) );
  OAI22X1 U1018 ( .A(n288), .B(n562), .C(n279), .D(n563), .Y(n742) );
  INVX1 U1019 ( .A(\memory[0][1] ), .Y(n279) );
  INVX1 U1020 ( .A(\memory[1][1] ), .Y(n288) );
  AOI22X1 U1021 ( .A(n564), .B(\memory[4][1] ), .C(n565), .D(\memory[5][1] ), 
        .Y(n740) );
  AOI22X1 U1022 ( .A(n566), .B(\memory[6][1] ), .C(n567), .D(\memory[7][1] ), 
        .Y(n739) );
  NAND3X1 U1023 ( .A(n744), .B(n745), .C(n746), .Y(n737) );
  NOR2X1 U1024 ( .A(n747), .B(n748), .Y(n746) );
  OAI22X1 U1025 ( .A(n375), .B(n573), .C(n383), .D(n574), .Y(n748) );
  INVX1 U1026 ( .A(\memory[9][1] ), .Y(n383) );
  INVX1 U1027 ( .A(\memory[8][1] ), .Y(n375) );
  OAI22X1 U1028 ( .A(n391), .B(n575), .C(n400), .D(n576), .Y(n747) );
  INVX1 U1029 ( .A(\memory[11][1] ), .Y(n400) );
  INVX1 U1030 ( .A(\memory[10][1] ), .Y(n391) );
  AOI22X1 U1031 ( .A(n577), .B(\memory[15][1] ), .C(n578), .D(\memory[14][1] ), 
        .Y(n745) );
  AOI22X1 U1032 ( .A(n579), .B(\memory[13][1] ), .C(n580), .D(\memory[12][1] ), 
        .Y(n744) );
  INVX1 U1033 ( .A(n749), .Y(n1329) );
  MUX2X1 U1034 ( .B(n750), .A(DATA[0]), .S(n522), .Y(n749) );
  NAND2X1 U1035 ( .A(n751), .B(n752), .Y(n750) );
  NOR2X1 U1036 ( .A(n753), .B(n754), .Y(n752) );
  NAND3X1 U1037 ( .A(n755), .B(n756), .C(n757), .Y(n754) );
  NOR2X1 U1038 ( .A(n758), .B(n759), .Y(n757) );
  OAI22X1 U1039 ( .A(n409), .B(n532), .C(n417), .D(n533), .Y(n759) );
  INVX1 U1040 ( .A(\memory[17][0] ), .Y(n417) );
  INVX1 U1041 ( .A(\memory[16][0] ), .Y(n409) );
  OAI22X1 U1042 ( .A(n425), .B(n534), .C(n433), .D(n535), .Y(n758) );
  INVX1 U1043 ( .A(\memory[19][0] ), .Y(n433) );
  INVX1 U1044 ( .A(\memory[18][0] ), .Y(n425) );
  AOI22X1 U1045 ( .A(n536), .B(\memory[23][0] ), .C(n537), .D(\memory[22][0] ), 
        .Y(n756) );
  AOI22X1 U1046 ( .A(n538), .B(\memory[21][0] ), .C(n539), .D(\memory[20][0] ), 
        .Y(n755) );
  NAND3X1 U1047 ( .A(n760), .B(n761), .C(n762), .Y(n753) );
  NOR2X1 U1048 ( .A(n763), .B(n764), .Y(n762) );
  OAI22X1 U1049 ( .A(n209), .B(n545), .C(n201), .D(n546), .Y(n764) );
  INVX1 U1050 ( .A(\memory[25][0] ), .Y(n201) );
  INVX1 U1051 ( .A(\memory[24][0] ), .Y(n209) );
  OAI22X1 U1052 ( .A(n192), .B(n547), .C(n182), .D(n548), .Y(n763) );
  INVX1 U1053 ( .A(\memory[27][0] ), .Y(n182) );
  INVX1 U1054 ( .A(\memory[26][0] ), .Y(n192) );
  AOI22X1 U1055 ( .A(n549), .B(\memory[31][0] ), .C(n550), .D(\memory[30][0] ), 
        .Y(n761) );
  AOI22X1 U1056 ( .A(n551), .B(\memory[29][0] ), .C(n552), .D(\memory[28][0] ), 
        .Y(n760) );
  NOR2X1 U1057 ( .A(n765), .B(n766), .Y(n751) );
  NAND3X1 U1058 ( .A(n767), .B(n768), .C(n769), .Y(n766) );
  NOR2X1 U1059 ( .A(n770), .B(n771), .Y(n769) );
  OAI22X1 U1060 ( .A(n303), .B(n560), .C(n295), .D(n561), .Y(n771) );
  INVX1 U1061 ( .A(\memory[2][0] ), .Y(n295) );
  INVX1 U1062 ( .A(\memory[3][0] ), .Y(n303) );
  OAI22X1 U1063 ( .A(n287), .B(n562), .C(n278), .D(n563), .Y(n770) );
  INVX1 U1064 ( .A(\memory[0][0] ), .Y(n278) );
  INVX1 U1065 ( .A(\memory[1][0] ), .Y(n287) );
  AOI22X1 U1066 ( .A(n564), .B(\memory[4][0] ), .C(n565), .D(\memory[5][0] ), 
        .Y(n768) );
  AOI22X1 U1067 ( .A(n566), .B(\memory[6][0] ), .C(n567), .D(\memory[7][0] ), 
        .Y(n767) );
  NAND3X1 U1068 ( .A(n772), .B(n773), .C(n774), .Y(n765) );
  NOR2X1 U1069 ( .A(n775), .B(n776), .Y(n774) );
  OAI22X1 U1070 ( .A(n376), .B(n573), .C(n384), .D(n574), .Y(n776) );
  INVX1 U1071 ( .A(\memory[9][0] ), .Y(n384) );
  INVX1 U1072 ( .A(\memory[8][0] ), .Y(n376) );
  OAI22X1 U1073 ( .A(n392), .B(n575), .C(n401), .D(n576), .Y(n775) );
  INVX1 U1074 ( .A(\memory[11][0] ), .Y(n401) );
  INVX1 U1075 ( .A(\memory[10][0] ), .Y(n392) );
  AOI22X1 U1076 ( .A(n577), .B(\memory[15][0] ), .C(n578), .D(\memory[14][0] ), 
        .Y(n773) );
  AOI22X1 U1077 ( .A(n579), .B(\memory[13][0] ), .C(n580), .D(\memory[12][0] ), 
        .Y(n772) );
  INVX1 U1078 ( .A(n777), .Y(n1330) );
  MUX2X1 U1079 ( .B(n778), .A(OUT_OPCODE[1]), .S(n522), .Y(n777) );
  NAND2X1 U1080 ( .A(n779), .B(n780), .Y(n778) );
  NOR2X1 U1081 ( .A(n781), .B(n782), .Y(n780) );
  NAND3X1 U1082 ( .A(n783), .B(n784), .C(n785), .Y(n782) );
  NOR2X1 U1083 ( .A(n786), .B(n787), .Y(n785) );
  OAI22X1 U1084 ( .A(n484), .B(n532), .C(n487), .D(n533), .Y(n787) );
  INVX1 U1085 ( .A(\opcode[17][1] ), .Y(n487) );
  INVX1 U1086 ( .A(\opcode[16][1] ), .Y(n484) );
  OAI22X1 U1087 ( .A(n490), .B(n534), .C(n493), .D(n535), .Y(n786) );
  INVX1 U1088 ( .A(\opcode[19][1] ), .Y(n493) );
  INVX1 U1089 ( .A(\opcode[18][1] ), .Y(n490) );
  AOI22X1 U1090 ( .A(n536), .B(\opcode[23][1] ), .C(n537), .D(\opcode[22][1] ), 
        .Y(n784) );
  AOI22X1 U1091 ( .A(n538), .B(\opcode[21][1] ), .C(n539), .D(\opcode[20][1] ), 
        .Y(n783) );
  NAND3X1 U1092 ( .A(n788), .B(n789), .C(n790), .Y(n781) );
  NOR2X1 U1093 ( .A(n791), .B(n792), .Y(n790) );
  OAI22X1 U1094 ( .A(n120), .B(n545), .C(n115), .D(n546), .Y(n792) );
  INVX1 U1095 ( .A(\opcode[25][1] ), .Y(n115) );
  INVX1 U1096 ( .A(\opcode[24][1] ), .Y(n120) );
  OAI22X1 U1097 ( .A(n110), .B(n547), .C(n104), .D(n548), .Y(n791) );
  INVX1 U1098 ( .A(\opcode[27][1] ), .Y(n104) );
  INVX1 U1099 ( .A(\opcode[26][1] ), .Y(n110) );
  AOI22X1 U1100 ( .A(n549), .B(\opcode[31][1] ), .C(n550), .D(\opcode[30][1] ), 
        .Y(n789) );
  AOI22X1 U1101 ( .A(n551), .B(\opcode[29][1] ), .C(n552), .D(\opcode[28][1] ), 
        .Y(n788) );
  NOR2X1 U1102 ( .A(n793), .B(n794), .Y(n779) );
  NAND3X1 U1103 ( .A(n795), .B(n796), .C(n797), .Y(n794) );
  NOR2X1 U1104 ( .A(n798), .B(n799), .Y(n797) );
  OAI22X1 U1105 ( .A(n174), .B(n560), .C(n171), .D(n561), .Y(n799) );
  INVX1 U1106 ( .A(\opcode[2][1] ), .Y(n171) );
  INVX1 U1107 ( .A(\opcode[3][1] ), .Y(n174) );
  OAI22X1 U1108 ( .A(n168), .B(n562), .C(n164), .D(n563), .Y(n798) );
  INVX1 U1109 ( .A(\opcode[0][1] ), .Y(n164) );
  INVX1 U1110 ( .A(\opcode[1][1] ), .Y(n168) );
  AOI22X1 U1111 ( .A(n564), .B(\opcode[4][1] ), .C(n565), .D(\opcode[5][1] ), 
        .Y(n796) );
  AOI22X1 U1112 ( .A(n566), .B(\opcode[6][1] ), .C(n567), .D(\opcode[7][1] ), 
        .Y(n795) );
  NAND3X1 U1113 ( .A(n800), .B(n801), .C(n802), .Y(n793) );
  NOR2X1 U1114 ( .A(n803), .B(n804), .Y(n802) );
  OAI22X1 U1115 ( .A(n469), .B(n573), .C(n472), .D(n574), .Y(n804) );
  INVX1 U1116 ( .A(\opcode[9][1] ), .Y(n472) );
  INVX1 U1117 ( .A(\opcode[8][1] ), .Y(n469) );
  OAI22X1 U1118 ( .A(n475), .B(n575), .C(n479), .D(n576), .Y(n803) );
  INVX1 U1119 ( .A(\opcode[11][1] ), .Y(n479) );
  INVX1 U1120 ( .A(\opcode[10][1] ), .Y(n475) );
  AOI22X1 U1121 ( .A(n577), .B(\opcode[15][1] ), .C(n578), .D(\opcode[14][1] ), 
        .Y(n801) );
  AOI22X1 U1122 ( .A(n579), .B(\opcode[13][1] ), .C(n580), .D(\opcode[12][1] ), 
        .Y(n800) );
  INVX1 U1123 ( .A(n805), .Y(n1331) );
  MUX2X1 U1124 ( .B(n806), .A(OUT_OPCODE[0]), .S(n522), .Y(n805) );
  NAND3X1 U1125 ( .A(N195), .B(n98), .C(n84), .Y(n522) );
  NAND2X1 U1126 ( .A(n807), .B(n808), .Y(n806) );
  NOR2X1 U1127 ( .A(n809), .B(n810), .Y(n808) );
  NAND3X1 U1128 ( .A(n811), .B(n812), .C(n813), .Y(n810) );
  NOR2X1 U1129 ( .A(n814), .B(n815), .Y(n813) );
  OAI22X1 U1130 ( .A(n486), .B(n532), .C(n489), .D(n533), .Y(n815) );
  NAND2X1 U1131 ( .A(n816), .B(n817), .Y(n533) );
  INVX1 U1132 ( .A(\opcode[17][0] ), .Y(n489) );
  NAND2X1 U1133 ( .A(n818), .B(n817), .Y(n532) );
  INVX1 U1134 ( .A(\opcode[16][0] ), .Y(n486) );
  OAI22X1 U1135 ( .A(n492), .B(n534), .C(n495), .D(n535), .Y(n814) );
  NAND2X1 U1136 ( .A(n816), .B(n819), .Y(n535) );
  INVX1 U1137 ( .A(\opcode[19][0] ), .Y(n495) );
  NAND2X1 U1138 ( .A(n818), .B(n819), .Y(n534) );
  INVX1 U1139 ( .A(\opcode[18][0] ), .Y(n492) );
  AOI22X1 U1140 ( .A(n536), .B(\opcode[23][0] ), .C(n537), .D(\opcode[22][0] ), 
        .Y(n812) );
  AOI22X1 U1141 ( .A(n538), .B(\opcode[21][0] ), .C(n539), .D(\opcode[20][0] ), 
        .Y(n811) );
  INVX1 U1142 ( .A(n822), .Y(n818) );
  NAND3X1 U1143 ( .A(n823), .B(n824), .C(readptr[4]), .Y(n822) );
  INVX1 U1144 ( .A(n825), .Y(n816) );
  NAND3X1 U1145 ( .A(readptr[0]), .B(n824), .C(readptr[4]), .Y(n825) );
  NAND3X1 U1146 ( .A(n826), .B(n827), .C(n828), .Y(n809) );
  NOR2X1 U1147 ( .A(n829), .B(n830), .Y(n828) );
  OAI22X1 U1148 ( .A(n122), .B(n545), .C(n117), .D(n546), .Y(n830) );
  NAND2X1 U1149 ( .A(n817), .B(n831), .Y(n546) );
  INVX1 U1150 ( .A(\opcode[25][0] ), .Y(n117) );
  NAND2X1 U1151 ( .A(n817), .B(n832), .Y(n545) );
  INVX1 U1152 ( .A(\opcode[24][0] ), .Y(n122) );
  OAI22X1 U1153 ( .A(n112), .B(n547), .C(n107), .D(n548), .Y(n829) );
  NAND2X1 U1154 ( .A(n819), .B(n831), .Y(n548) );
  INVX1 U1155 ( .A(\opcode[27][0] ), .Y(n107) );
  NAND2X1 U1156 ( .A(n819), .B(n832), .Y(n547) );
  INVX1 U1157 ( .A(\opcode[26][0] ), .Y(n112) );
  AOI22X1 U1158 ( .A(n549), .B(\opcode[31][0] ), .C(n550), .D(\opcode[30][0] ), 
        .Y(n827) );
  AOI22X1 U1159 ( .A(n551), .B(\opcode[29][0] ), .C(n552), .D(\opcode[28][0] ), 
        .Y(n826) );
  INVX1 U1160 ( .A(n833), .Y(n832) );
  NAND3X1 U1161 ( .A(readptr[3]), .B(n823), .C(readptr[4]), .Y(n833) );
  INVX1 U1162 ( .A(n834), .Y(n831) );
  NAND3X1 U1163 ( .A(readptr[3]), .B(readptr[0]), .C(readptr[4]), .Y(n834) );
  NOR2X1 U1164 ( .A(n835), .B(n836), .Y(n807) );
  NAND3X1 U1165 ( .A(n837), .B(n838), .C(n839), .Y(n836) );
  NOR2X1 U1166 ( .A(n840), .B(n841), .Y(n839) );
  OAI22X1 U1167 ( .A(n172), .B(n560), .C(n169), .D(n561), .Y(n841) );
  NAND2X1 U1168 ( .A(n842), .B(n819), .Y(n561) );
  INVX1 U1169 ( .A(\opcode[2][0] ), .Y(n169) );
  NAND2X1 U1170 ( .A(n843), .B(n819), .Y(n560) );
  INVX1 U1171 ( .A(\opcode[3][0] ), .Y(n172) );
  OAI22X1 U1172 ( .A(n166), .B(n562), .C(n162), .D(n563), .Y(n840) );
  NAND2X1 U1173 ( .A(n842), .B(n817), .Y(n563) );
  INVX1 U1174 ( .A(\opcode[0][0] ), .Y(n162) );
  NAND2X1 U1175 ( .A(n843), .B(n817), .Y(n562) );
  INVX1 U1176 ( .A(\opcode[1][0] ), .Y(n166) );
  AOI22X1 U1177 ( .A(n564), .B(\opcode[4][0] ), .C(n565), .D(\opcode[5][0] ), 
        .Y(n838) );
  AOI22X1 U1178 ( .A(n566), .B(\opcode[6][0] ), .C(n567), .D(\opcode[7][0] ), 
        .Y(n837) );
  INVX1 U1179 ( .A(n844), .Y(n843) );
  NAND3X1 U1180 ( .A(n824), .B(n845), .C(readptr[0]), .Y(n844) );
  INVX1 U1181 ( .A(n846), .Y(n842) );
  NAND3X1 U1182 ( .A(n824), .B(n845), .C(n823), .Y(n846) );
  INVX1 U1183 ( .A(readptr[3]), .Y(n824) );
  NAND3X1 U1184 ( .A(n847), .B(n848), .C(n849), .Y(n835) );
  NOR2X1 U1185 ( .A(n850), .B(n851), .Y(n849) );
  OAI22X1 U1186 ( .A(n471), .B(n573), .C(n474), .D(n574), .Y(n851) );
  NAND2X1 U1187 ( .A(n852), .B(n817), .Y(n574) );
  INVX1 U1188 ( .A(\opcode[9][0] ), .Y(n474) );
  NAND2X1 U1189 ( .A(n853), .B(n817), .Y(n573) );
  NOR2X1 U1190 ( .A(readptr[1]), .B(readptr[2]), .Y(n817) );
  INVX1 U1191 ( .A(\opcode[8][0] ), .Y(n471) );
  OAI22X1 U1192 ( .A(n477), .B(n575), .C(n481), .D(n576), .Y(n850) );
  NAND2X1 U1193 ( .A(n852), .B(n819), .Y(n576) );
  INVX1 U1194 ( .A(\opcode[11][0] ), .Y(n481) );
  NAND2X1 U1195 ( .A(n853), .B(n819), .Y(n575) );
  NOR2X1 U1196 ( .A(n517), .B(readptr[2]), .Y(n819) );
  INVX1 U1197 ( .A(\opcode[10][0] ), .Y(n477) );
  AOI22X1 U1198 ( .A(n577), .B(\opcode[15][0] ), .C(n578), .D(\opcode[14][0] ), 
        .Y(n848) );
  NOR2X1 U1199 ( .A(n517), .B(n855), .Y(n820) );
  AOI22X1 U1200 ( .A(n579), .B(\opcode[13][0] ), .C(n580), .D(\opcode[12][0] ), 
        .Y(n847) );
  INVX1 U1201 ( .A(n857), .Y(n853) );
  NAND3X1 U1202 ( .A(n823), .B(n845), .C(readptr[3]), .Y(n857) );
  INVX1 U1203 ( .A(readptr[0]), .Y(n823) );
  NOR2X1 U1204 ( .A(n855), .B(readptr[1]), .Y(n821) );
  INVX1 U1205 ( .A(readptr[2]), .Y(n855) );
  INVX1 U1207 ( .A(n859), .Y(n852) );
  NAND3X1 U1208 ( .A(readptr[0]), .B(n845), .C(readptr[3]), .Y(n859) );
  INVX1 U1209 ( .A(readptr[4]), .Y(n845) );
  AND2X1 U1210 ( .A(N337), .B(n84), .Y(N347) );
  AND2X1 U1211 ( .A(N336), .B(n84), .Y(N346) );
  AND2X1 U1212 ( .A(N335), .B(n84), .Y(N345) );
  AND2X1 U1213 ( .A(N334), .B(n84), .Y(N344) );
  AND2X1 U1214 ( .A(N333), .B(n84), .Y(N343) );
  AND2X1 U1215 ( .A(N193), .B(n84), .Y(N342) );
  AND2X1 U1216 ( .A(N192), .B(n84), .Y(N341) );
  AND2X1 U1217 ( .A(N191), .B(n84), .Y(N340) );
  AND2X1 U1218 ( .A(N190), .B(n84), .Y(N339) );
  AND2X1 U1219 ( .A(N189), .B(n84), .Y(N338) );
  AND2X1 U1220 ( .A(R_ENABLE), .B(n313), .Y(N195) );
  NAND3X1 U1221 ( .A(n861), .B(n863), .C(n864), .Y(n313) );
  NOR2X1 U1222 ( .A(n865), .B(n866), .Y(n864) );
  XOR2X1 U1223 ( .A(writeptr[4]), .B(readptr[4]), .Y(n866) );
  XOR2X1 U1224 ( .A(n83), .B(readptr[3]), .Y(n865) );
  XOR2X1 U1225 ( .A(n517), .B(n78), .Y(n863) );
  INVX1 U1226 ( .A(readptr[1]), .Y(n517) );
  NOR2X1 U1227 ( .A(n867), .B(n909), .Y(n861) );
  XOR2X1 U1228 ( .A(n81), .B(readptr[0]), .Y(n909) );
  XOR2X1 U1229 ( .A(n76), .B(readptr[2]), .Y(n867) );
endmodule


module memoryblock_0 ( CLK, NEXT_BYTE, RCV_DATA, RCV_OPCODE, RST, W_ENABLE, 
        EOP, EMPTY, FULL, B_READY, PRGA_IN, PRGA_OPCODE );
  input [7:0] RCV_DATA;
  input [1:0] RCV_OPCODE;
  output [7:0] PRGA_IN;
  output [1:0] PRGA_OPCODE;
  input CLK, NEXT_BYTE, RST, W_ENABLE, EOP;
  output EMPTY, FULL, B_READY;
  wire   R_ENABLE;
  wire   [4:0] BYTE_COUNT;
  wire   [7:0] DATA;
  wire   [1:0] OUT_OPCODE;

  RBUFFER_0 U_0 ( .CLK(CLK), .RST(RST), .NEXT_BYTE(NEXT_BYTE), .DATA(DATA), 
        .OPCODE(OUT_OPCODE), .BYTE_COUNT(BYTE_COUNT), .EOP(EOP), .B_READY(
        B_READY), .R_ENABLE(R_ENABLE), .PRGA_IN(PRGA_IN), .PRGA_OPCODE(
        PRGA_OPCODE) );
  RFIFO_0 U_1 ( .CLK(CLK), .RST(RST), .W_ENABLE(W_ENABLE), .R_ENABLE(R_ENABLE), 
        .RCV_DATA(RCV_DATA), .RCV_OPCODE(RCV_OPCODE), .DATA(DATA), 
        .OUT_OPCODE(OUT_OPCODE), .BYTE_COUNT(BYTE_COUNT), .EMPTY(EMPTY), 
        .FULL(FULL) );
endmodule


module rx_CRC_CALC_0 ( CLK, RST, W_ENABLE, OPCODE, RCV_DATA, RX_CRC );
  input [1:0] OPCODE;
  input [7:0] RCV_DATA;
  output [15:0] RX_CRC;
  input CLK, RST, W_ENABLE;
  wire   n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n56, n60, n79, n80, n81, n82, n100, n102, n104,
         n106, n108, n110, n112, n114, n116, n118, n120, n122, n124, n126,
         n128, n130, n131, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246;
  wire   [15:0] current_crc;
  wire   [15:0] cache_1;

  DFFPOSX1 \cache_1_reg[0]  ( .D(n173), .CLK(CLK), .Q(cache_1[0]) );
  DFFPOSX1 \cache_1_reg[8]  ( .D(n174), .CLK(CLK), .Q(cache_1[8]) );
  DFFPOSX1 \cache_1_reg[15]  ( .D(n175), .CLK(CLK), .Q(cache_1[15]) );
  DFFPOSX1 \cache_1_reg[1]  ( .D(n176), .CLK(CLK), .Q(cache_1[1]) );
  DFFPOSX1 \cache_1_reg[9]  ( .D(n177), .CLK(CLK), .Q(cache_1[9]) );
  DFFPOSX1 \cache_1_reg[2]  ( .D(n178), .CLK(CLK), .Q(cache_1[2]) );
  DFFPOSX1 \cache_1_reg[10]  ( .D(n179), .CLK(CLK), .Q(cache_1[10]) );
  DFFPOSX1 \cache_1_reg[3]  ( .D(n180), .CLK(CLK), .Q(cache_1[3]) );
  DFFPOSX1 \cache_1_reg[11]  ( .D(n181), .CLK(CLK), .Q(cache_1[11]) );
  DFFPOSX1 \cache_1_reg[4]  ( .D(n182), .CLK(CLK), .Q(cache_1[4]) );
  DFFPOSX1 \cache_1_reg[12]  ( .D(n183), .CLK(CLK), .Q(cache_1[12]) );
  DFFPOSX1 \cache_1_reg[5]  ( .D(n184), .CLK(CLK), .Q(cache_1[5]) );
  DFFPOSX1 \cache_1_reg[13]  ( .D(n185), .CLK(CLK), .Q(cache_1[13]) );
  DFFPOSX1 \cache_1_reg[6]  ( .D(n186), .CLK(CLK), .Q(cache_1[6]) );
  DFFPOSX1 \cache_1_reg[14]  ( .D(n187), .CLK(CLK), .Q(cache_1[14]) );
  DFFPOSX1 \cache_1_reg[7]  ( .D(n188), .CLK(CLK), .Q(cache_1[7]) );
  DFFPOSX1 \cache_2_reg[15]  ( .D(n189), .CLK(CLK), .Q(RX_CRC[15]) );
  DFFPOSX1 \cache_2_reg[14]  ( .D(n190), .CLK(CLK), .Q(RX_CRC[14]) );
  DFFPOSX1 \cache_2_reg[13]  ( .D(n191), .CLK(CLK), .Q(RX_CRC[13]) );
  DFFPOSX1 \cache_2_reg[12]  ( .D(n192), .CLK(CLK), .Q(RX_CRC[12]) );
  DFFPOSX1 \cache_2_reg[11]  ( .D(n193), .CLK(CLK), .Q(RX_CRC[11]) );
  DFFPOSX1 \cache_2_reg[10]  ( .D(n194), .CLK(CLK), .Q(RX_CRC[10]) );
  DFFPOSX1 \cache_2_reg[9]  ( .D(n195), .CLK(CLK), .Q(RX_CRC[9]) );
  DFFPOSX1 \cache_2_reg[8]  ( .D(n196), .CLK(CLK), .Q(RX_CRC[8]) );
  DFFPOSX1 \cache_2_reg[7]  ( .D(n197), .CLK(CLK), .Q(RX_CRC[7]) );
  DFFPOSX1 \cache_2_reg[6]  ( .D(n198), .CLK(CLK), .Q(RX_CRC[6]) );
  DFFPOSX1 \cache_2_reg[5]  ( .D(n199), .CLK(CLK), .Q(RX_CRC[5]) );
  DFFPOSX1 \cache_2_reg[4]  ( .D(n200), .CLK(CLK), .Q(RX_CRC[4]) );
  DFFPOSX1 \cache_2_reg[3]  ( .D(n201), .CLK(CLK), .Q(RX_CRC[3]) );
  DFFPOSX1 \cache_2_reg[2]  ( .D(n202), .CLK(CLK), .Q(RX_CRC[2]) );
  DFFPOSX1 \cache_2_reg[1]  ( .D(n203), .CLK(CLK), .Q(RX_CRC[1]) );
  DFFPOSX1 \cache_2_reg[0]  ( .D(n204), .CLK(CLK), .Q(RX_CRC[0]) );
  OAI21X1 U3 ( .A(n42), .B(n60), .C(n246), .Y(n204) );
  NAND2X1 U4 ( .A(RX_CRC[0]), .B(n43), .Y(n246) );
  OAI21X1 U5 ( .A(n41), .B(n102), .C(n245), .Y(n203) );
  NAND2X1 U6 ( .A(RX_CRC[1]), .B(n43), .Y(n245) );
  OAI21X1 U7 ( .A(n41), .B(n110), .C(n244), .Y(n202) );
  NAND2X1 U8 ( .A(RX_CRC[2]), .B(n43), .Y(n244) );
  OAI21X1 U9 ( .A(n41), .B(n118), .C(n243), .Y(n201) );
  NAND2X1 U10 ( .A(RX_CRC[3]), .B(n43), .Y(n243) );
  OAI21X1 U11 ( .A(n41), .B(n126), .C(n242), .Y(n200) );
  NAND2X1 U12 ( .A(RX_CRC[4]), .B(n43), .Y(n242) );
  OAI21X1 U13 ( .A(n41), .B(n148), .C(n241), .Y(n199) );
  NAND2X1 U14 ( .A(RX_CRC[5]), .B(n42), .Y(n241) );
  OAI21X1 U15 ( .A(n41), .B(n152), .C(n240), .Y(n198) );
  NAND2X1 U16 ( .A(RX_CRC[6]), .B(n42), .Y(n240) );
  OAI21X1 U17 ( .A(n41), .B(n156), .C(n239), .Y(n197) );
  NAND2X1 U18 ( .A(RX_CRC[7]), .B(n42), .Y(n239) );
  OAI21X1 U19 ( .A(n41), .B(n80), .C(n238), .Y(n196) );
  NAND2X1 U20 ( .A(RX_CRC[8]), .B(n42), .Y(n238) );
  OAI21X1 U21 ( .A(n41), .B(n106), .C(n237), .Y(n195) );
  NAND2X1 U22 ( .A(RX_CRC[9]), .B(n42), .Y(n237) );
  OAI21X1 U23 ( .A(n42), .B(n114), .C(n236), .Y(n194) );
  NAND2X1 U24 ( .A(RX_CRC[10]), .B(n42), .Y(n236) );
  OAI21X1 U25 ( .A(n42), .B(n122), .C(n235), .Y(n193) );
  NAND2X1 U26 ( .A(RX_CRC[11]), .B(n42), .Y(n235) );
  OAI21X1 U27 ( .A(n42), .B(n130), .C(n234), .Y(n192) );
  NAND2X1 U28 ( .A(RX_CRC[12]), .B(n42), .Y(n234) );
  OAI21X1 U29 ( .A(n42), .B(n150), .C(n233), .Y(n191) );
  NAND2X1 U30 ( .A(RX_CRC[13]), .B(n43), .Y(n233) );
  OAI21X1 U31 ( .A(n42), .B(n154), .C(n232), .Y(n190) );
  NAND2X1 U32 ( .A(RX_CRC[14]), .B(n43), .Y(n232) );
  OAI21X1 U33 ( .A(n42), .B(n82), .C(n231), .Y(n189) );
  NAND2X1 U34 ( .A(RX_CRC[15]), .B(n43), .Y(n231) );
  OAI22X1 U35 ( .A(n41), .B(n155), .C(n39), .D(n156), .Y(n188) );
  OAI22X1 U37 ( .A(n41), .B(n153), .C(n39), .D(n154), .Y(n187) );
  OAI22X1 U39 ( .A(n41), .B(n151), .C(n39), .D(n152), .Y(n186) );
  OAI22X1 U41 ( .A(n41), .B(n149), .C(n39), .D(n150), .Y(n185) );
  OAI22X1 U43 ( .A(n40), .B(n131), .C(n39), .D(n148), .Y(n184) );
  OAI22X1 U45 ( .A(n40), .B(n128), .C(n39), .D(n130), .Y(n183) );
  OAI22X1 U47 ( .A(n40), .B(n124), .C(n39), .D(n126), .Y(n182) );
  OAI22X1 U49 ( .A(n40), .B(n120), .C(n39), .D(n122), .Y(n181) );
  OAI22X1 U51 ( .A(n40), .B(n116), .C(n39), .D(n118), .Y(n180) );
  OAI22X1 U53 ( .A(n40), .B(n112), .C(n38), .D(n114), .Y(n179) );
  OAI22X1 U55 ( .A(n40), .B(n108), .C(n38), .D(n110), .Y(n178) );
  OAI22X1 U57 ( .A(n40), .B(n104), .C(n38), .D(n106), .Y(n177) );
  OAI22X1 U59 ( .A(n40), .B(n100), .C(n38), .D(n102), .Y(n176) );
  OAI22X1 U61 ( .A(n40), .B(n81), .C(n38), .D(n82), .Y(n175) );
  OAI22X1 U63 ( .A(n40), .B(n79), .C(n38), .D(n80), .Y(n174) );
  OAI22X1 U65 ( .A(n40), .B(n56), .C(n38), .D(n60), .Y(n173) );
  OAI22X1 U70 ( .A(n81), .B(n37), .C(n228), .D(n35), .Y(n172) );
  XOR2X1 U71 ( .A(n227), .B(current_crc[7]), .Y(n228) );
  OAI22X1 U72 ( .A(n35), .B(n151), .C(n153), .D(n37), .Y(n171) );
  OAI22X1 U73 ( .A(n35), .B(n131), .C(n149), .D(n229), .Y(n170) );
  OAI22X1 U74 ( .A(n230), .B(n124), .C(n128), .D(n37), .Y(n169) );
  OAI22X1 U75 ( .A(n35), .B(n116), .C(n120), .D(n229), .Y(n168) );
  OAI22X1 U77 ( .A(n230), .B(n108), .C(n112), .D(n37), .Y(n167) );
  OAI22X1 U78 ( .A(n104), .B(n37), .C(n226), .D(n230), .Y(n166) );
  XOR2X1 U79 ( .A(n100), .B(n45), .Y(n226) );
  OAI22X1 U80 ( .A(n79), .B(n229), .C(n225), .D(n35), .Y(n165) );
  XOR2X1 U81 ( .A(n224), .B(n223), .Y(n225) );
  XOR2X1 U82 ( .A(n56), .B(n45), .Y(n224) );
  OAI22X1 U84 ( .A(n155), .B(n37), .C(n46), .D(n230), .Y(n164) );
  OAI22X1 U86 ( .A(n151), .B(n229), .C(n222), .D(n35), .Y(n163) );
  XOR2X1 U87 ( .A(n221), .B(n220), .Y(n222) );
  OAI22X1 U89 ( .A(n131), .B(n37), .C(n219), .D(n230), .Y(n162) );
  OAI22X1 U91 ( .A(n124), .B(n229), .C(n218), .D(n35), .Y(n161) );
  XOR2X1 U92 ( .A(n217), .B(n216), .Y(n218) );
  OAI22X1 U94 ( .A(n116), .B(n37), .C(n215), .D(n230), .Y(n160) );
  OAI22X1 U96 ( .A(n108), .B(n229), .C(n214), .D(n35), .Y(n159) );
  XOR2X1 U97 ( .A(n213), .B(n212), .Y(n214) );
  OAI22X1 U99 ( .A(n100), .B(n37), .C(n211), .D(n230), .Y(n158) );
  XOR2X1 U100 ( .A(n210), .B(n209), .Y(n211) );
  XOR2X1 U101 ( .A(n208), .B(n207), .Y(n210) );
  OAI22X1 U103 ( .A(n56), .B(n229), .C(n227), .D(n35), .Y(n157) );
  XOR2X1 U104 ( .A(n206), .B(n205), .Y(n227) );
  XOR2X1 U105 ( .A(n45), .B(n212), .Y(n205) );
  XOR2X1 U106 ( .A(current_crc[8]), .B(RCV_DATA[0]), .Y(n212) );
  XOR2X1 U108 ( .A(n81), .B(RCV_DATA[7]), .Y(n208) );
  XOR2X1 U110 ( .A(n46), .B(n207), .Y(n206) );
  XOR2X1 U111 ( .A(n215), .B(n219), .Y(n207) );
  XNOR2X1 U112 ( .A(n220), .B(n216), .Y(n219) );
  XOR2X1 U113 ( .A(current_crc[11]), .B(RCV_DATA[3]), .Y(n216) );
  XNOR2X1 U114 ( .A(n128), .B(RCV_DATA[4]), .Y(n220) );
  XOR2X1 U116 ( .A(n213), .B(n48), .Y(n215) );
  XOR2X1 U118 ( .A(n112), .B(RCV_DATA[2]), .Y(n217) );
  XOR2X1 U120 ( .A(n104), .B(RCV_DATA[1]), .Y(n213) );
  XOR2X1 U123 ( .A(n223), .B(n47), .Y(n209) );
  XOR2X1 U125 ( .A(n149), .B(RCV_DATA[5]), .Y(n221) );
  XNOR2X1 U127 ( .A(n153), .B(RCV_DATA[6]), .Y(n223) );
  OAI21X1 U129 ( .A(n50), .B(n49), .C(n230), .Y(n229) );
  NAND3X1 U130 ( .A(OPCODE[0]), .B(n49), .C(W_ENABLE), .Y(n230) );
  DFFSR \current_crc_reg[14]  ( .D(n171), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[14]) );
  DFFSR \current_crc_reg[12]  ( .D(n169), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[12]) );
  DFFSR \current_crc_reg[10]  ( .D(n167), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[10]) );
  DFFSR \current_crc_reg[13]  ( .D(n170), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[13]) );
  DFFSR \current_crc_reg[11]  ( .D(n168), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[11]) );
  DFFSR \current_crc_reg[15]  ( .D(n172), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[15]) );
  DFFSR \current_crc_reg[8]  ( .D(n165), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[8]) );
  DFFSR \current_crc_reg[6]  ( .D(n163), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[6]) );
  DFFSR \current_crc_reg[4]  ( .D(n161), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[4]) );
  DFFSR \current_crc_reg[2]  ( .D(n159), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[2]) );
  DFFSR \current_crc_reg[0]  ( .D(n157), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[0]) );
  DFFSR \current_crc_reg[9]  ( .D(n166), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[9]) );
  DFFSR \current_crc_reg[7]  ( .D(n164), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[7]) );
  DFFSR \current_crc_reg[5]  ( .D(n162), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[5]) );
  DFFSR \current_crc_reg[3]  ( .D(n160), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[3]) );
  DFFSR \current_crc_reg[1]  ( .D(n158), .CLK(CLK), .R(n44), .S(1'b1), .Q(
        current_crc[1]) );
  INVX2 U36 ( .A(n32), .Y(n38) );
  INVX2 U68 ( .A(n230), .Y(n34) );
  BUFX2 U69 ( .A(n32), .Y(n43) );
  INVX2 U76 ( .A(n32), .Y(n39) );
  OR2X2 U83 ( .A(n35), .B(RST), .Y(n32) );
  INVX2 U85 ( .A(n34), .Y(n35) );
  INVX2 U88 ( .A(n36), .Y(n37) );
  INVX2 U90 ( .A(n229), .Y(n36) );
  INVX2 U93 ( .A(RST), .Y(n44) );
  INVX1 U95 ( .A(OPCODE[0]), .Y(n50) );
  INVX1 U98 ( .A(OPCODE[1]), .Y(n49) );
  BUFX4 U102 ( .A(n32), .Y(n40) );
  BUFX4 U107 ( .A(n32), .Y(n41) );
  BUFX4 U109 ( .A(n32), .Y(n42) );
  INVX2 U115 ( .A(n208), .Y(n45) );
  INVX2 U117 ( .A(n209), .Y(n46) );
  INVX2 U119 ( .A(n221), .Y(n47) );
  INVX2 U121 ( .A(n217), .Y(n48) );
  INVX2 U122 ( .A(current_crc[0]), .Y(n56) );
  INVX2 U124 ( .A(cache_1[0]), .Y(n60) );
  INVX2 U126 ( .A(current_crc[8]), .Y(n79) );
  INVX2 U128 ( .A(cache_1[8]), .Y(n80) );
  INVX2 U131 ( .A(current_crc[15]), .Y(n81) );
  INVX2 U132 ( .A(cache_1[15]), .Y(n82) );
  INVX2 U133 ( .A(current_crc[1]), .Y(n100) );
  INVX2 U134 ( .A(cache_1[1]), .Y(n102) );
  INVX2 U135 ( .A(current_crc[9]), .Y(n104) );
  INVX2 U136 ( .A(cache_1[9]), .Y(n106) );
  INVX2 U137 ( .A(current_crc[2]), .Y(n108) );
  INVX2 U138 ( .A(cache_1[2]), .Y(n110) );
  INVX2 U139 ( .A(current_crc[10]), .Y(n112) );
  INVX2 U140 ( .A(cache_1[10]), .Y(n114) );
  INVX2 U141 ( .A(current_crc[3]), .Y(n116) );
  INVX2 U142 ( .A(cache_1[3]), .Y(n118) );
  INVX2 U143 ( .A(current_crc[11]), .Y(n120) );
  INVX2 U144 ( .A(cache_1[11]), .Y(n122) );
  INVX2 U145 ( .A(current_crc[4]), .Y(n124) );
  INVX2 U146 ( .A(cache_1[4]), .Y(n126) );
  INVX2 U147 ( .A(current_crc[12]), .Y(n128) );
  INVX2 U148 ( .A(cache_1[12]), .Y(n130) );
  INVX2 U149 ( .A(current_crc[5]), .Y(n131) );
  INVX2 U150 ( .A(cache_1[5]), .Y(n148) );
  INVX2 U151 ( .A(current_crc[13]), .Y(n149) );
  INVX2 U152 ( .A(cache_1[13]), .Y(n150) );
  INVX2 U153 ( .A(current_crc[6]), .Y(n151) );
  INVX2 U154 ( .A(cache_1[6]), .Y(n152) );
  INVX2 U155 ( .A(current_crc[14]), .Y(n153) );
  INVX2 U156 ( .A(cache_1[14]), .Y(n154) );
  INVX2 U157 ( .A(current_crc[7]), .Y(n155) );
  INVX2 U158 ( .A(cache_1[7]), .Y(n156) );
endmodule


module rx_accumulator_0 ( CLK, RST, RCV_DATA, W_ENABLE, rx_CHECK_CRC );
  input [7:0] RCV_DATA;
  output [15:0] rx_CHECK_CRC;
  input CLK, RST, W_ENABLE;
  wire   n40, n42, n44, n46, n48, n50, n52, n54, n56, n57, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91;

  OAI21X1 U2 ( .A(n40), .B(n59), .C(n91), .Y(n75) );
  NAND2X1 U3 ( .A(rx_CHECK_CRC[8]), .B(n40), .Y(n91) );
  OAI21X1 U4 ( .A(n42), .B(n59), .C(n90), .Y(n74) );
  NAND2X1 U5 ( .A(RCV_DATA[0]), .B(n42), .Y(n90) );
  OAI21X1 U7 ( .A(n40), .B(n57), .C(n89), .Y(n73) );
  NAND2X1 U8 ( .A(rx_CHECK_CRC[9]), .B(n40), .Y(n89) );
  OAI21X1 U9 ( .A(n42), .B(n57), .C(n88), .Y(n72) );
  NAND2X1 U10 ( .A(RCV_DATA[1]), .B(n42), .Y(n88) );
  OAI21X1 U12 ( .A(n40), .B(n56), .C(n87), .Y(n71) );
  NAND2X1 U13 ( .A(rx_CHECK_CRC[10]), .B(n40), .Y(n87) );
  OAI21X1 U14 ( .A(n42), .B(n56), .C(n86), .Y(n70) );
  NAND2X1 U15 ( .A(RCV_DATA[2]), .B(n42), .Y(n86) );
  OAI21X1 U17 ( .A(n40), .B(n54), .C(n85), .Y(n69) );
  NAND2X1 U18 ( .A(rx_CHECK_CRC[11]), .B(n40), .Y(n85) );
  OAI21X1 U19 ( .A(n42), .B(n54), .C(n84), .Y(n68) );
  NAND2X1 U20 ( .A(RCV_DATA[3]), .B(n42), .Y(n84) );
  OAI21X1 U22 ( .A(n40), .B(n52), .C(n83), .Y(n67) );
  NAND2X1 U23 ( .A(rx_CHECK_CRC[12]), .B(n40), .Y(n83) );
  OAI21X1 U24 ( .A(n42), .B(n52), .C(n82), .Y(n66) );
  NAND2X1 U25 ( .A(RCV_DATA[4]), .B(n42), .Y(n82) );
  OAI21X1 U27 ( .A(n40), .B(n50), .C(n81), .Y(n65) );
  NAND2X1 U28 ( .A(rx_CHECK_CRC[13]), .B(n40), .Y(n81) );
  OAI21X1 U29 ( .A(n42), .B(n50), .C(n80), .Y(n64) );
  NAND2X1 U30 ( .A(RCV_DATA[5]), .B(n42), .Y(n80) );
  OAI21X1 U32 ( .A(n40), .B(n48), .C(n79), .Y(n63) );
  NAND2X1 U33 ( .A(rx_CHECK_CRC[14]), .B(n40), .Y(n79) );
  OAI21X1 U34 ( .A(n42), .B(n48), .C(n78), .Y(n62) );
  NAND2X1 U35 ( .A(RCV_DATA[6]), .B(n42), .Y(n78) );
  OAI21X1 U37 ( .A(n40), .B(n46), .C(n77), .Y(n61) );
  NAND2X1 U38 ( .A(rx_CHECK_CRC[15]), .B(n40), .Y(n77) );
  OAI21X1 U41 ( .A(n42), .B(n46), .C(n76), .Y(n60) );
  NAND2X1 U42 ( .A(RCV_DATA[7]), .B(n42), .Y(n76) );
  DFFSR \present_CHECK_CRC_reg[7]  ( .D(n60), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[7]) );
  DFFSR \present_CHECK_CRC_reg[6]  ( .D(n62), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[6]) );
  DFFSR \present_CHECK_CRC_reg[5]  ( .D(n64), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[5]) );
  DFFSR \present_CHECK_CRC_reg[4]  ( .D(n66), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[4]) );
  DFFSR \present_CHECK_CRC_reg[3]  ( .D(n68), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[3]) );
  DFFSR \present_CHECK_CRC_reg[2]  ( .D(n70), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[2]) );
  DFFSR \present_CHECK_CRC_reg[1]  ( .D(n72), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[1]) );
  DFFSR \present_CHECK_CRC_reg[0]  ( .D(n74), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[0]) );
  DFFSR \present_CHECK_CRC_reg[15]  ( .D(n61), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[15]) );
  DFFSR \present_CHECK_CRC_reg[14]  ( .D(n63), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[14]) );
  DFFSR \present_CHECK_CRC_reg[13]  ( .D(n65), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[13]) );
  DFFSR \present_CHECK_CRC_reg[12]  ( .D(n67), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[12]) );
  DFFSR \present_CHECK_CRC_reg[11]  ( .D(n69), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[11]) );
  DFFSR \present_CHECK_CRC_reg[10]  ( .D(n71), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[10]) );
  DFFSR \present_CHECK_CRC_reg[9]  ( .D(n73), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[9]) );
  DFFSR \present_CHECK_CRC_reg[8]  ( .D(n75), .CLK(CLK), .R(n44), .S(1'b1), 
        .Q(rx_CHECK_CRC[8]) );
  INVX2 U50 ( .A(n40), .Y(n42) );
  INVX2 U51 ( .A(W_ENABLE), .Y(n40) );
  INVX2 U52 ( .A(RST), .Y(n44) );
  INVX2 U53 ( .A(rx_CHECK_CRC[7]), .Y(n46) );
  INVX2 U54 ( .A(rx_CHECK_CRC[6]), .Y(n48) );
  INVX2 U55 ( .A(rx_CHECK_CRC[5]), .Y(n50) );
  INVX2 U56 ( .A(rx_CHECK_CRC[4]), .Y(n52) );
  INVX2 U57 ( .A(rx_CHECK_CRC[3]), .Y(n54) );
  INVX2 U58 ( .A(rx_CHECK_CRC[2]), .Y(n56) );
  INVX2 U59 ( .A(rx_CHECK_CRC[1]), .Y(n57) );
  INVX2 U60 ( .A(rx_CHECK_CRC[0]), .Y(n59) );
endmodule


module rx_decode_0 ( CLK, RST, DP1_RX, SHIFT_ENABLE, EOP, D_ORIG, BITSTUFF, 
        BS_ERROR );
  input CLK, RST, DP1_RX, SHIFT_ENABLE, EOP;
  output D_ORIG, BITSTUFF, BS_ERROR;
  wire   DP_hold1, DP_hold2, N29, N30, N31, N32, n6, n8, n9, n10, n12, n13,
         n14, n15, n16, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74;
  wire   [3:0] state;

  DFFSR DP_hold2_reg ( .D(n47), .CLK(CLK), .R(1'b1), .S(n6), .Q(DP_hold2) );
  DFFSR DP_hold1_reg ( .D(n48), .CLK(CLK), .R(1'b1), .S(n6), .Q(DP_hold1) );
  OR2X2 U10 ( .A(n8), .B(state[1]), .Y(n55) );
  NAND2X1 U20 ( .A(n74), .B(n73), .Y(n48) );
  AOI22X1 U21 ( .A(DP_hold1), .B(n12), .C(DP1_RX), .D(n72), .Y(n74) );
  NAND2X1 U22 ( .A(n71), .B(n73), .Y(n47) );
  AOI22X1 U23 ( .A(n10), .B(DP_hold1), .C(DP_hold2), .D(n70), .Y(n71) );
  NAND2X1 U24 ( .A(SHIFT_ENABLE), .B(n72), .Y(n70) );
  XNOR2X1 U25 ( .A(DP_hold1), .B(DP_hold2), .Y(D_ORIG) );
  NOR2X1 U26 ( .A(n69), .B(EOP), .Y(N32) );
  AOI21X1 U27 ( .A(n68), .B(BITSTUFF), .C(BS_ERROR), .Y(n69) );
  NAND3X1 U28 ( .A(state[3]), .B(n16), .C(n66), .Y(n67) );
  NOR2X1 U29 ( .A(state[2]), .B(state[1]), .Y(n66) );
  NOR2X1 U30 ( .A(n72), .B(state[3]), .Y(BITSTUFF) );
  NOR2X1 U31 ( .A(n65), .B(n14), .Y(N31) );
  AOI21X1 U32 ( .A(state[2]), .B(n64), .C(n63), .Y(n65) );
  OAI21X1 U33 ( .A(n62), .B(n61), .C(n60), .Y(n63) );
  NAND2X1 U34 ( .A(state[0]), .B(n68), .Y(n61) );
  NAND2X1 U35 ( .A(state[1]), .B(n15), .Y(n62) );
  OAI21X1 U36 ( .A(state[1]), .B(n59), .C(SHIFT_ENABLE), .Y(n64) );
  NOR2X1 U37 ( .A(n58), .B(n14), .Y(N30) );
  AOI21X1 U38 ( .A(state[1]), .B(n57), .C(n56), .Y(n58) );
  OAI21X1 U39 ( .A(n16), .B(n55), .C(n60), .Y(n56) );
  NAND2X1 U40 ( .A(n12), .B(n59), .Y(n60) );
  NAND2X1 U41 ( .A(n13), .B(n16), .Y(n72) );
  OAI21X1 U42 ( .A(n59), .B(n54), .C(SHIFT_ENABLE), .Y(n57) );
  NAND2X1 U43 ( .A(n16), .B(n15), .Y(n54) );
  NOR2X1 U44 ( .A(n53), .B(n14), .Y(N29) );
  NOR2X1 U45 ( .A(EOP), .B(state[3]), .Y(n73) );
  AOI21X1 U46 ( .A(state[0]), .B(n9), .C(n52), .Y(n53) );
  OAI21X1 U47 ( .A(n8), .B(n51), .C(n50), .Y(n52) );
  NAND3X1 U48 ( .A(n13), .B(n59), .C(SHIFT_ENABLE), .Y(n50) );
  NAND2X1 U49 ( .A(n49), .B(n16), .Y(n51) );
  NAND2X1 U50 ( .A(state[2]), .B(state[1]), .Y(n49) );
  NOR2X1 U51 ( .A(n59), .B(n9), .Y(n68) );
  XOR2X1 U52 ( .A(DP1_RX), .B(DP_hold2), .Y(n59) );
  DFFSR \state_reg[3]  ( .D(N32), .CLK(CLK), .R(n6), .S(1'b1), .Q(state[3]) );
  DFFSR \state_reg[0]  ( .D(N29), .CLK(CLK), .R(n6), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[2]  ( .D(N31), .CLK(CLK), .R(n6), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[1]  ( .D(N30), .CLK(CLK), .R(n6), .S(1'b1), .Q(state[1]) );
  INVX2 U8 ( .A(RST), .Y(n6) );
  INVX2 U11 ( .A(n68), .Y(n8) );
  INVX2 U12 ( .A(SHIFT_ENABLE), .Y(n9) );
  INVX2 U13 ( .A(n70), .Y(n10) );
  INVX2 U14 ( .A(n67), .Y(BS_ERROR) );
  INVX2 U15 ( .A(n72), .Y(n12) );
  INVX2 U16 ( .A(n49), .Y(n13) );
  INVX2 U17 ( .A(n73), .Y(n14) );
  INVX2 U18 ( .A(state[2]), .Y(n15) );
  INVX2 U19 ( .A(state[0]), .Y(n16) );
endmodule


module rx_edgedetect_0 ( CLK, RST, DP1_RX, D_EDGE );
  input CLK, RST, DP1_RX;
  output D_EDGE;
  wire   DP_hold1, DP_hold2, n2, n5;

  DFFSR DP_hold1_reg ( .D(DP1_RX), .CLK(CLK), .R(1'b1), .S(n2), .Q(DP_hold1)
         );
  DFFSR DP_hold2_reg ( .D(DP_hold1), .CLK(CLK), .R(1'b1), .S(n2), .Q(DP_hold2)
         );
  NOR2X1 U6 ( .A(RST), .B(n5), .Y(D_EDGE) );
  XNOR2X1 U7 ( .A(DP_hold2), .B(DP_hold1), .Y(n5) );
  INVX2 U4 ( .A(RST), .Y(n2) );
endmodule


module rx_eopdetect_0 ( DP1_RX, DM1_RX, EOP );
  input DP1_RX, DM1_RX;
  output EOP;


  NOR2X1 U1 ( .A(DP1_RX), .B(DM1_RX), .Y(EOP) );
endmodule


module rx_rcu_0 ( CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR, 
        RX_CRC, RX_CHECK_CRC, RCV_DATA, RCVING, W_ENABLE, R_ERROR, CRC_ERROR, 
        OPCODE );
  input [15:0] RX_CRC;
  input [15:0] RX_CHECK_CRC;
  input [7:0] RCV_DATA;
  output [1:0] OPCODE;
  input CLK, RST, D_EDGE, EOP, SHIFT_ENABLE, BITSTUFF, BS_ERROR;
  output RCVING, W_ENABLE, R_ERROR, CRC_ERROR;
  wire   nxtR_ERROR, curR_ERROR, curCRC_ERROR, n1, n2, n18, n19, n23, n24, n25,
         n26, n28, n30, n35, n43, n44, n49, n58, n64, n68, n69, n73, n76, n82,
         n93, n101, n104, n108, n110, n112, n114, n115, n118, n124, n128, n130,
         n131, n132, n135, n141, n143, n148, n149, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297;
  wire   [3:0] state;
  wire   [3:0] count;
  wire   [3:0] nextstate;

  DFFPOSX1 curCRC_ERROR_reg ( .D(n196), .CLK(CLK), .Q(curCRC_ERROR) );
  DFFPOSX1 curR_ERROR_reg ( .D(n197), .CLK(CLK), .Q(curR_ERROR) );
  DFFPOSX1 CRC_ERROR_reg ( .D(n172), .CLK(CLK), .Q(CRC_ERROR) );
  OAI21X1 U5 ( .A(EOP), .B(n23), .C(n294), .Y(n295) );
  AOI22X1 U6 ( .A(BS_ERROR), .B(n293), .C(n292), .D(n44), .Y(n294) );
  OAI21X1 U7 ( .A(n192), .B(n26), .C(n291), .Y(n292) );
  AOI22X1 U8 ( .A(n290), .B(D_EDGE), .C(n19), .D(n289), .Y(n291) );
  OAI21X1 U9 ( .A(n183), .B(n190), .C(n184), .Y(n289) );
  NOR2X1 U11 ( .A(n183), .B(n177), .Y(n290) );
  OAI21X1 U12 ( .A(n288), .B(n24), .C(n287), .Y(n293) );
  OAI21X1 U13 ( .A(n2), .B(n286), .C(n285), .Y(n296) );
  NAND2X1 U15 ( .A(n178), .B(n282), .Y(n286) );
  NAND2X1 U16 ( .A(n281), .B(n280), .Y(nextstate[2]) );
  NOR2X1 U17 ( .A(n279), .B(n278), .Y(n280) );
  OAI21X1 U18 ( .A(n26), .B(n277), .C(n283), .Y(n278) );
  OAI21X1 U19 ( .A(n2), .B(n276), .C(n49), .Y(n277) );
  NAND2X1 U20 ( .A(n179), .B(n187), .Y(n276) );
  NAND2X1 U21 ( .A(n275), .B(n274), .Y(n279) );
  NOR2X1 U22 ( .A(n273), .B(n272), .Y(n281) );
  OAI22X1 U23 ( .A(n171), .B(n44), .C(n271), .D(n190), .Y(n272) );
  OAI21X1 U24 ( .A(n49), .B(n270), .C(n269), .Y(n273) );
  OAI21X1 U25 ( .A(n268), .B(n267), .C(n266), .Y(n269) );
  AOI22X1 U26 ( .A(n265), .B(n264), .C(n282), .D(n192), .Y(n270) );
  NOR2X1 U27 ( .A(D_EDGE), .B(n183), .Y(n265) );
  OAI21X1 U28 ( .A(n170), .B(n192), .C(n263), .Y(nextstate[1]) );
  OAI21X1 U30 ( .A(n260), .B(n259), .C(n190), .Y(n262) );
  OAI21X1 U31 ( .A(n287), .B(n180), .C(n258), .Y(n259) );
  OAI21X1 U33 ( .A(n23), .B(n256), .C(n175), .Y(n260) );
  NAND2X1 U34 ( .A(n181), .B(n192), .Y(n256) );
  OAI22X1 U35 ( .A(n255), .B(n254), .C(n44), .D(n253), .Y(nextstate[0]) );
  OAI21X1 U36 ( .A(n183), .B(n28), .C(n252), .Y(n253) );
  NAND3X1 U37 ( .A(n190), .B(n183), .C(n251), .Y(n252) );
  OAI21X1 U38 ( .A(n25), .B(n192), .C(n250), .Y(n251) );
  AOI22X1 U39 ( .A(n257), .B(n249), .C(n248), .D(n247), .Y(n250) );
  OAI22X1 U42 ( .A(state[0]), .B(n184), .C(n246), .D(n183), .Y(n254) );
  AOI22X1 U43 ( .A(EOP), .B(n249), .C(D_EDGE), .D(n174), .Y(n246) );
  OAI21X1 U45 ( .A(n35), .B(n244), .C(n243), .Y(n255) );
  NOR2X1 U46 ( .A(n49), .B(n282), .Y(n243) );
  AOI22X1 U47 ( .A(n242), .B(n257), .C(D_EDGE), .D(n249), .Y(n244) );
  NOR2X1 U48 ( .A(n181), .B(EOP), .Y(n257) );
  NOR2X1 U50 ( .A(BS_ERROR), .B(n25), .Y(n242) );
  AOI21X1 U52 ( .A(CRC_ERROR), .B(RST), .C(n240), .Y(n241) );
  OAI21X1 U53 ( .A(n239), .B(n238), .C(n237), .Y(n240) );
  NAND2X1 U54 ( .A(curCRC_ERROR), .B(n236), .Y(n238) );
  NAND2X1 U55 ( .A(n58), .B(n44), .Y(n239) );
  OAI21X1 U56 ( .A(n58), .B(n189), .C(n235), .Y(n197) );
  AOI21X1 U57 ( .A(n297), .B(n58), .C(n173), .Y(n235) );
  NAND3X1 U59 ( .A(n233), .B(n44), .C(curR_ERROR), .Y(n234) );
  OAI21X1 U60 ( .A(n19), .B(n183), .C(n232), .Y(n233) );
  OAI21X1 U61 ( .A(n178), .B(n26), .C(n231), .Y(n297) );
  OAI21X1 U64 ( .A(n19), .B(n247), .C(n177), .Y(n229) );
  OAI21X1 U65 ( .A(n267), .B(n176), .C(EOP), .Y(n230) );
  OAI21X1 U69 ( .A(n227), .B(n188), .C(n237), .Y(n196) );
  NAND3X1 U70 ( .A(n2), .B(n58), .C(n226), .Y(n237) );
  NOR2X1 U71 ( .A(n26), .B(n228), .Y(n226) );
  NAND3X1 U72 ( .A(n49), .B(n187), .C(n179), .Y(n228) );
  AOI21X1 U76 ( .A(n236), .B(n44), .C(RST), .Y(n227) );
  OAI21X1 U77 ( .A(n183), .B(n25), .C(n232), .Y(n236) );
  NAND2X1 U78 ( .A(n288), .B(n245), .Y(n232) );
  NOR2X1 U79 ( .A(D_EDGE), .B(n35), .Y(n245) );
  OAI21X1 U81 ( .A(n224), .B(n185), .C(n223), .Y(n195) );
  NAND3X1 U82 ( .A(n165), .B(n185), .C(count[0]), .Y(n223) );
  AOI21X1 U83 ( .A(n222), .B(n182), .C(n221), .Y(n224) );
  OAI21X1 U84 ( .A(n159), .B(n186), .C(n220), .Y(n194) );
  NAND3X1 U85 ( .A(n219), .B(n186), .C(n160), .Y(n220) );
  OAI21X1 U87 ( .A(n217), .B(n187), .C(n216), .Y(n193) );
  NAND3X1 U88 ( .A(n219), .B(n187), .C(n215), .Y(n216) );
  NOR2X1 U89 ( .A(n214), .B(n186), .Y(n215) );
  AOI21X1 U90 ( .A(n222), .B(n186), .C(n218), .Y(n217) );
  OAI21X1 U91 ( .A(n160), .B(n168), .C(n274), .Y(n218) );
  NAND3X1 U93 ( .A(count[1]), .B(count[0]), .C(n213), .Y(n214) );
  AOI22X1 U95 ( .A(n221), .B(count[0]), .C(n182), .D(n165), .Y(n212) );
  NAND3X1 U97 ( .A(n219), .B(n191), .C(SHIFT_ENABLE), .Y(n211) );
  OAI21X1 U100 ( .A(n213), .B(n168), .C(n274), .Y(n221) );
  NAND2X1 U101 ( .A(EOP), .B(n210), .Y(n274) );
  NOR2X1 U103 ( .A(n266), .B(n169), .Y(n222) );
  NOR2X1 U104 ( .A(n187), .B(n225), .Y(n266) );
  NAND3X1 U105 ( .A(n185), .B(n186), .C(n182), .Y(n225) );
  NOR2X1 U110 ( .A(BITSTUFF), .B(n164), .Y(n213) );
  NAND3X1 U115 ( .A(n208), .B(n166), .C(n248), .Y(n284) );
  NAND3X1 U117 ( .A(n207), .B(n206), .C(n205), .Y(n247) );
  NOR2X1 U119 ( .A(RCV_DATA[6]), .B(RCV_DATA[5]), .Y(n203) );
  NOR2X1 U120 ( .A(RCV_DATA[4]), .B(RCV_DATA[3]), .Y(n204) );
  NOR2X1 U121 ( .A(RCV_DATA[2]), .B(RCV_DATA[1]), .Y(n206) );
  NOR2X1 U122 ( .A(RCV_DATA[0]), .B(n167), .Y(n207) );
  NAND3X1 U124 ( .A(n170), .B(n261), .C(n271), .Y(RCVING) );
  NOR2X1 U125 ( .A(n210), .B(n202), .Y(n271) );
  OAI21X1 U126 ( .A(n24), .B(n43), .C(n209), .Y(n202) );
  NAND3X1 U127 ( .A(n35), .B(n44), .C(n288), .Y(n209) );
  OAI21X1 U129 ( .A(n49), .B(n26), .C(n283), .Y(n201) );
  NAND3X1 U130 ( .A(n35), .B(n44), .C(n249), .Y(n283) );
  NAND3X1 U131 ( .A(n200), .B(n199), .C(n169), .Y(OPCODE[1]) );
  NAND3X1 U133 ( .A(n23), .B(n287), .C(n175), .Y(n210) );
  NOR2X1 U135 ( .A(n25), .B(n24), .Y(n268) );
  NOR2X1 U141 ( .A(n44), .B(state[2]), .Y(n208) );
  OAI21X1 U144 ( .A(n183), .B(n171), .C(n44), .Y(n199) );
  NOR2X1 U146 ( .A(n174), .B(state[0]), .Y(n288) );
  OAI21X1 U148 ( .A(n198), .B(n19), .C(n49), .Y(n200) );
  NOR2X1 U149 ( .A(state[0]), .B(n183), .Y(n198) );
  OAI21X1 U150 ( .A(n44), .B(n26), .C(n261), .Y(OPCODE[0]) );
  NAND3X1 U151 ( .A(n49), .B(n35), .C(n264), .Y(n261) );
  NOR2X1 U155 ( .A(n43), .B(n183), .Y(n282) );
  OR2X2 U3 ( .A(n297), .B(n173), .Y(nxtR_ERROR) );
  OR2X2 U4 ( .A(n296), .B(n295), .Y(nextstate[3]) );
  AND2X2 U14 ( .A(n284), .B(n283), .Y(n285) );
  AND2X2 U29 ( .A(n262), .B(n261), .Y(n263) );
  AND2X2 U62 ( .A(n230), .B(n275), .Y(n231) );
  OR2X2 U63 ( .A(n24), .B(n229), .Y(n275) );
  AND2X2 U99 ( .A(n222), .B(n274), .Y(n219) );
  AND2X2 U114 ( .A(n284), .B(n209), .Y(n258) );
  AND2X2 U118 ( .A(n204), .B(n203), .Y(n205) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(CLK), .R(n58), .S(1'b1), .Q(
        state[1]) );
  DFFSR R_ERROR_reg ( .D(nxtR_ERROR), .CLK(CLK), .R(n58), .S(1'b1), .Q(R_ERROR) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(CLK), .R(n58), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(CLK), .R(n58), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(CLK), .R(n58), .S(1'b1), .Q(
        state[3]) );
  DFFSR \count_reg[0]  ( .D(n158), .CLK(CLK), .R(n58), .S(1'b1), .Q(count[0])
         );
  DFFSR \count_reg[1]  ( .D(n195), .CLK(CLK), .R(n58), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n194), .CLK(CLK), .R(n58), .S(1'b1), .Q(count[2])
         );
  DFFSR \count_reg[3]  ( .D(n193), .CLK(CLK), .R(n58), .S(1'b1), .Q(count[3])
         );
  AND2X2 U10 ( .A(n183), .B(n44), .Y(n1) );
  NAND2X1 U32 ( .A(n154), .B(n153), .Y(n2) );
  INVX2 U73 ( .A(state[3]), .Y(n18) );
  INVX2 U74 ( .A(n18), .Y(n19) );
  OR2X2 U75 ( .A(n28), .B(n24), .Y(n23) );
  INVX2 U80 ( .A(n23), .Y(n267) );
  NAND2X1 U86 ( .A(n264), .B(n1), .Y(n287) );
  INVX2 U92 ( .A(state[2]), .Y(n183) );
  INVX2 U94 ( .A(n25), .Y(n264) );
  INVX1 U96 ( .A(n287), .Y(n176) );
  OR2X2 U98 ( .A(n44), .B(state[2]), .Y(n24) );
  OR2X2 U102 ( .A(n177), .B(n19), .Y(n25) );
  OR2X2 U106 ( .A(n43), .B(n183), .Y(n26) );
  OR2X1 U107 ( .A(state[0]), .B(n19), .Y(n43) );
  OR2X2 U108 ( .A(n177), .B(n174), .Y(n28) );
  INVX1 U109 ( .A(n28), .Y(n249) );
  INVX2 U111 ( .A(n258), .Y(n30) );
  OR2X2 U112 ( .A(n30), .B(OPCODE[0]), .Y(W_ENABLE) );
  INVX2 U113 ( .A(RST), .Y(n58) );
  INVX1 U116 ( .A(n183), .Y(n35) );
  INVX1 U123 ( .A(n43), .Y(n248) );
  INVX2 U128 ( .A(state[1]), .Y(n44) );
  INVX1 U132 ( .A(n44), .Y(n49) );
  XNOR2X1 U134 ( .A(RX_CHECK_CRC[10]), .B(RX_CRC[10]), .Y(n76) );
  XNOR2X1 U136 ( .A(RX_CHECK_CRC[9]), .B(RX_CRC[9]), .Y(n73) );
  XOR2X1 U137 ( .A(RX_CHECK_CRC[7]), .B(RX_CRC[7]), .Y(n68) );
  XOR2X1 U138 ( .A(RX_CHECK_CRC[8]), .B(RX_CRC[8]), .Y(n64) );
  NOR2X1 U139 ( .A(n68), .B(n64), .Y(n69) );
  NAND3X1 U140 ( .A(n76), .B(n73), .C(n69), .Y(n112) );
  XNOR2X1 U142 ( .A(RX_CHECK_CRC[14]), .B(RX_CRC[14]), .Y(n108) );
  XNOR2X1 U143 ( .A(RX_CHECK_CRC[13]), .B(RX_CRC[13]), .Y(n104) );
  XOR2X1 U145 ( .A(RX_CHECK_CRC[11]), .B(RX_CRC[11]), .Y(n93) );
  XOR2X1 U147 ( .A(RX_CHECK_CRC[12]), .B(RX_CRC[12]), .Y(n82) );
  NOR2X1 U152 ( .A(n93), .B(n82), .Y(n101) );
  NAND3X1 U153 ( .A(n108), .B(n104), .C(n101), .Y(n110) );
  NOR2X1 U154 ( .A(n112), .B(n110), .Y(n154) );
  NOR2X1 U156 ( .A(n155), .B(RX_CHECK_CRC[0]), .Y(n114) );
  OAI22X1 U157 ( .A(RX_CRC[1]), .B(n114), .C(n114), .D(n157), .Y(n131) );
  AND2X1 U158 ( .A(RX_CHECK_CRC[0]), .B(n155), .Y(n115) );
  OAI22X1 U159 ( .A(n115), .B(n156), .C(RX_CHECK_CRC[1]), .D(n115), .Y(n130)
         );
  XOR2X1 U160 ( .A(RX_CHECK_CRC[15]), .B(RX_CRC[15]), .Y(n124) );
  XOR2X1 U161 ( .A(RX_CHECK_CRC[2]), .B(RX_CRC[2]), .Y(n118) );
  NOR2X1 U162 ( .A(n124), .B(n118), .Y(n128) );
  NAND3X1 U163 ( .A(n131), .B(n130), .C(n128), .Y(n152) );
  XNOR2X1 U164 ( .A(RX_CHECK_CRC[6]), .B(RX_CRC[6]), .Y(n148) );
  XNOR2X1 U165 ( .A(RX_CHECK_CRC[5]), .B(RX_CRC[5]), .Y(n143) );
  XOR2X1 U166 ( .A(RX_CHECK_CRC[3]), .B(RX_CRC[3]), .Y(n135) );
  XOR2X1 U167 ( .A(RX_CHECK_CRC[4]), .B(RX_CRC[4]), .Y(n132) );
  NOR2X1 U168 ( .A(n135), .B(n132), .Y(n141) );
  NAND3X1 U169 ( .A(n148), .B(n143), .C(n141), .Y(n149) );
  NOR2X1 U170 ( .A(n152), .B(n149), .Y(n153) );
  INVX2 U171 ( .A(RX_CRC[0]), .Y(n155) );
  INVX2 U172 ( .A(RX_CRC[1]), .Y(n156) );
  INVX2 U173 ( .A(RX_CHECK_CRC[1]), .Y(n157) );
  INVX2 U174 ( .A(n212), .Y(n158) );
  INVX2 U175 ( .A(n218), .Y(n159) );
  INVX2 U176 ( .A(n214), .Y(n160) );
  INVX2 U177 ( .A(SHIFT_ENABLE), .Y(n164) );
  INVX2 U178 ( .A(n211), .Y(n165) );
  INVX2 U179 ( .A(n247), .Y(n166) );
  INVX2 U180 ( .A(RCV_DATA[7]), .Y(n167) );
  INVX2 U181 ( .A(n222), .Y(n168) );
  INVX2 U182 ( .A(n210), .Y(n169) );
  INVX2 U183 ( .A(n201), .Y(n170) );
  INVX2 U184 ( .A(n288), .Y(n171) );
  INVX2 U185 ( .A(n241), .Y(n172) );
  INVX2 U186 ( .A(n234), .Y(n173) );
  INVX2 U187 ( .A(n19), .Y(n174) );
  INVX2 U188 ( .A(n268), .Y(n175) );
  INVX2 U189 ( .A(state[0]), .Y(n177) );
  INVX2 U190 ( .A(n228), .Y(n178) );
  INVX2 U191 ( .A(n225), .Y(n179) );
  INVX2 U192 ( .A(n257), .Y(n180) );
  INVX2 U193 ( .A(n266), .Y(n181) );
  INVX2 U194 ( .A(count[0]), .Y(n182) );
  INVX2 U195 ( .A(n245), .Y(n184) );
  INVX2 U196 ( .A(count[1]), .Y(n185) );
  INVX2 U197 ( .A(count[2]), .Y(n186) );
  INVX2 U198 ( .A(count[3]), .Y(n187) );
  INVX2 U199 ( .A(curCRC_ERROR), .Y(n188) );
  INVX2 U200 ( .A(curR_ERROR), .Y(n189) );
  INVX2 U201 ( .A(BS_ERROR), .Y(n190) );
  INVX2 U202 ( .A(BITSTUFF), .Y(n191) );
  INVX2 U203 ( .A(EOP), .Y(n192) );
endmodule


module rx_shift_reg_0 ( CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF, RCV_DATA );
  output [7:0] RCV_DATA;
  input CLK, RST, SHIFT_ENABLE, D_ORIG, BITSTUFF;
  wire   n17, n20, n22, n25, n28, n31, n34, n37, n40, n43, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71;
  wire   [7:0] present_val;

  DFFPOSX1 \RCV_DATA_reg[7]  ( .D(n47), .CLK(CLK), .Q(RCV_DATA[7]) );
  DFFPOSX1 \RCV_DATA_reg[6]  ( .D(n49), .CLK(CLK), .Q(RCV_DATA[6]) );
  DFFPOSX1 \RCV_DATA_reg[5]  ( .D(n51), .CLK(CLK), .Q(RCV_DATA[5]) );
  DFFPOSX1 \RCV_DATA_reg[4]  ( .D(n53), .CLK(CLK), .Q(RCV_DATA[4]) );
  DFFPOSX1 \RCV_DATA_reg[3]  ( .D(n55), .CLK(CLK), .Q(RCV_DATA[3]) );
  DFFPOSX1 \RCV_DATA_reg[2]  ( .D(n57), .CLK(CLK), .Q(RCV_DATA[2]) );
  DFFPOSX1 \RCV_DATA_reg[1]  ( .D(n59), .CLK(CLK), .Q(RCV_DATA[1]) );
  DFFPOSX1 \RCV_DATA_reg[0]  ( .D(n61), .CLK(CLK), .Q(RCV_DATA[0]) );
  OAI21X1 U2 ( .A(RST), .B(n43), .C(n71), .Y(n61) );
  NAND2X1 U3 ( .A(RCV_DATA[0]), .B(RST), .Y(n71) );
  OAI22X1 U4 ( .A(n20), .B(n43), .C(n70), .D(n40), .Y(n60) );
  OAI21X1 U6 ( .A(RST), .B(n40), .C(n69), .Y(n59) );
  NAND2X1 U7 ( .A(RCV_DATA[1]), .B(RST), .Y(n69) );
  OAI22X1 U8 ( .A(n20), .B(n40), .C(n70), .D(n37), .Y(n58) );
  OAI21X1 U10 ( .A(RST), .B(n37), .C(n68), .Y(n57) );
  NAND2X1 U11 ( .A(RCV_DATA[2]), .B(RST), .Y(n68) );
  OAI22X1 U12 ( .A(n20), .B(n37), .C(n70), .D(n34), .Y(n56) );
  OAI21X1 U14 ( .A(RST), .B(n34), .C(n67), .Y(n55) );
  NAND2X1 U15 ( .A(RCV_DATA[3]), .B(RST), .Y(n67) );
  OAI22X1 U16 ( .A(n20), .B(n34), .C(n70), .D(n31), .Y(n54) );
  OAI21X1 U18 ( .A(RST), .B(n31), .C(n66), .Y(n53) );
  NAND2X1 U19 ( .A(RCV_DATA[4]), .B(RST), .Y(n66) );
  OAI22X1 U20 ( .A(n20), .B(n31), .C(n70), .D(n28), .Y(n52) );
  OAI21X1 U22 ( .A(RST), .B(n28), .C(n65), .Y(n51) );
  NAND2X1 U23 ( .A(RCV_DATA[5]), .B(RST), .Y(n65) );
  OAI22X1 U24 ( .A(n20), .B(n28), .C(n70), .D(n25), .Y(n50) );
  OAI21X1 U26 ( .A(RST), .B(n25), .C(n64), .Y(n49) );
  NAND2X1 U27 ( .A(RCV_DATA[6]), .B(RST), .Y(n64) );
  OAI22X1 U28 ( .A(n20), .B(n25), .C(n70), .D(n22), .Y(n48) );
  OAI21X1 U30 ( .A(RST), .B(n22), .C(n63), .Y(n47) );
  NAND2X1 U31 ( .A(RCV_DATA[7]), .B(RST), .Y(n63) );
  OAI21X1 U32 ( .A(n20), .B(n22), .C(n62), .Y(n46) );
  NAND2X1 U33 ( .A(D_ORIG), .B(n20), .Y(n62) );
  NAND2X1 U36 ( .A(SHIFT_ENABLE), .B(n45), .Y(n70) );
  DFFSR \present_val_reg[7]  ( .D(n46), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[7]) );
  DFFSR \present_val_reg[6]  ( .D(n48), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[6]) );
  DFFSR \present_val_reg[5]  ( .D(n50), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[5]) );
  DFFSR \present_val_reg[4]  ( .D(n52), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[4]) );
  DFFSR \present_val_reg[3]  ( .D(n54), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[3]) );
  DFFSR \present_val_reg[2]  ( .D(n56), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[2]) );
  DFFSR \present_val_reg[1]  ( .D(n58), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[1]) );
  DFFSR \present_val_reg[0]  ( .D(n60), .CLK(CLK), .R(n17), .S(1'b1), .Q(
        present_val[0]) );
  INVX2 U5 ( .A(n70), .Y(n20) );
  INVX2 U37 ( .A(RST), .Y(n17) );
  INVX2 U38 ( .A(present_val[7]), .Y(n22) );
  INVX2 U39 ( .A(present_val[6]), .Y(n25) );
  INVX2 U40 ( .A(present_val[5]), .Y(n28) );
  INVX2 U41 ( .A(present_val[4]), .Y(n31) );
  INVX2 U42 ( .A(present_val[3]), .Y(n34) );
  INVX2 U43 ( .A(present_val[2]), .Y(n37) );
  INVX2 U44 ( .A(present_val[1]), .Y(n40) );
  INVX2 U45 ( .A(present_val[0]), .Y(n43) );
  INVX2 U46 ( .A(BITSTUFF), .Y(n45) );
endmodule


module rx_timer_0 ( CLK, RST, D_EDGE, RCVING, SHIFT_ENABLE );
  input CLK, RST, D_EDGE, RCVING;
  output SHIFT_ENABLE;
  wire   state, n6, n7, n8, n9, n10, n11, n12, n19, n20, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34;
  wire   [3:0] count;
  wire   [3:0] nextcount;

  NOR2X1 U17 ( .A(n34), .B(n33), .Y(nextcount[3]) );
  AOI22X1 U18 ( .A(n32), .B(n31), .C(n30), .D(count[3]), .Y(n34) );
  XOR2X1 U19 ( .A(n29), .B(n31), .Y(n30) );
  NOR2X1 U20 ( .A(count[3]), .B(n20), .Y(n32) );
  NOR2X1 U23 ( .A(n27), .B(n33), .Y(nextcount[1]) );
  NAND2X1 U24 ( .A(state), .B(n26), .Y(nextcount[0]) );
  OAI21X1 U25 ( .A(D_EDGE), .B(n19), .C(RCVING), .Y(n26) );
  NAND3X1 U28 ( .A(RCVING), .B(n25), .C(state), .Y(n33) );
  OAI21X1 U29 ( .A(n27), .B(n24), .C(n28), .Y(n29) );
  NAND2X1 U30 ( .A(count[0]), .B(count[1]), .Y(n28) );
  XOR2X1 U31 ( .A(n24), .B(n27), .Y(n31) );
  XNOR2X1 U32 ( .A(count[0]), .B(count[1]), .Y(n27) );
  DFFSR state_reg ( .D(RCVING), .CLK(CLK), .R(n11), .S(1'b1), .Q(state) );
  DFFSR \count_reg[2]  ( .D(nextcount[2]), .CLK(CLK), .R(n11), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[0]  ( .D(nextcount[0]), .CLK(CLK), .R(n11), .S(1'b1), .Q(
        count[0]) );
  DFFSR \count_reg[3]  ( .D(nextcount[3]), .CLK(CLK), .R(n11), .S(1'b1), .Q(
        count[3]) );
  DFFSR \count_reg[1]  ( .D(nextcount[1]), .CLK(CLK), .R(n11), .S(1'b1), .Q(
        count[1]) );
  AND2X1 U8 ( .A(n12), .B(count[3]), .Y(n7) );
  INVX2 U9 ( .A(n8), .Y(nextcount[2]) );
  INVX2 U10 ( .A(RST), .Y(n11) );
  AND2X2 U11 ( .A(n6), .B(n7), .Y(SHIFT_ENABLE) );
  NOR2X1 U12 ( .A(n31), .B(n29), .Y(n6) );
  OAI21X1 U13 ( .A(n9), .B(n10), .C(RCVING), .Y(n8) );
  NAND2X1 U14 ( .A(n25), .B(state), .Y(n9) );
  XNOR2X1 U15 ( .A(n28), .B(count[2]), .Y(n10) );
  INVX2 U16 ( .A(n33), .Y(n12) );
  INVX2 U21 ( .A(count[0]), .Y(n19) );
  INVX2 U22 ( .A(n29), .Y(n20) );
  INVX2 U26 ( .A(count[2]), .Y(n24) );
  INVX2 U27 ( .A(D_EDGE), .Y(n25) );
endmodule


module receiver_block_rewire_0 ( CLK, DM1_RX, DP1_RX, RST, BS_ERROR, CRC_ERROR, 
        EOP_external, OPCODE, RCV_DATA, R_ERROR, W_ENABLE );
  output [1:0] OPCODE;
  output [7:0] RCV_DATA;
  input CLK, DM1_RX, DP1_RX, RST;
  output BS_ERROR, CRC_ERROR, EOP_external, R_ERROR, W_ENABLE;
  wire   SHIFT_ENABLE, BITSTUFF, D_ORIG, D_EDGE, RCVING, n1, n2;
  wire   [15:0] RX_CRC;
  wire   [15:0] rx_CHECK_CRC;

  rx_CRC_CALC_0 U_2 ( .CLK(CLK), .RST(n1), .W_ENABLE(W_ENABLE), .OPCODE(OPCODE), .RCV_DATA(RCV_DATA), .RX_CRC(RX_CRC) );
  rx_accumulator_0 U_3 ( .CLK(CLK), .RST(n1), .RCV_DATA(RCV_DATA), .W_ENABLE(
        W_ENABLE), .rx_CHECK_CRC(rx_CHECK_CRC) );
  rx_decode_0 U_1 ( .CLK(CLK), .RST(n1), .DP1_RX(DP1_RX), .SHIFT_ENABLE(
        SHIFT_ENABLE), .EOP(EOP_external), .D_ORIG(D_ORIG), .BITSTUFF(BITSTUFF), .BS_ERROR(BS_ERROR) );
  rx_edgedetect_0 U_0 ( .CLK(CLK), .RST(n1), .DP1_RX(DP1_RX), .D_EDGE(D_EDGE)
         );
  rx_eopdetect_0 U_4 ( .DP1_RX(DP1_RX), .DM1_RX(DM1_RX), .EOP(EOP_external) );
  rx_rcu_0 U_5 ( .CLK(CLK), .RST(n1), .D_EDGE(D_EDGE), .EOP(EOP_external), 
        .SHIFT_ENABLE(SHIFT_ENABLE), .BITSTUFF(BITSTUFF), .BS_ERROR(BS_ERROR), 
        .RX_CRC(RX_CRC), .RX_CHECK_CRC(rx_CHECK_CRC), .RCV_DATA(RCV_DATA), 
        .RCVING(RCVING), .W_ENABLE(W_ENABLE), .R_ERROR(R_ERROR), .CRC_ERROR(
        CRC_ERROR), .OPCODE(OPCODE) );
  rx_shift_reg_0 U_6 ( .CLK(CLK), .RST(n1), .SHIFT_ENABLE(SHIFT_ENABLE), 
        .D_ORIG(D_ORIG), .BITSTUFF(BITSTUFF), .RCV_DATA(RCV_DATA) );
  rx_timer_0 U_7 ( .CLK(CLK), .RST(n1), .D_EDGE(D_EDGE), .RCVING(RCVING), 
        .SHIFT_ENABLE(SHIFT_ENABLE) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module tx_CRC_CALC_0 ( CLK, RST, EOP, T_STROBE, PRGA_OPCODE, PRGA_OUT, TX_CRC
 );
  input [1:0] PRGA_OPCODE;
  input [7:0] PRGA_OUT;
  output [15:0] TX_CRC;
  input CLK, RST, EOP, T_STROBE;
  wire   n1, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122;

  OAI22X1 U39 ( .A(n25), .B(n20), .C(n122), .D(n19), .Y(n97) );
  XNOR2X1 U40 ( .A(n120), .B(n80), .Y(n122) );
  OAI22X1 U41 ( .A(n79), .B(n20), .C(n19), .D(n37), .Y(n96) );
  OAI22X1 U42 ( .A(n36), .B(n20), .C(n19), .D(n35), .Y(n95) );
  OAI22X1 U43 ( .A(n34), .B(n20), .C(n19), .D(n33), .Y(n94) );
  OAI22X1 U44 ( .A(n32), .B(n20), .C(n19), .D(n31), .Y(n93) );
  OAI22X1 U45 ( .A(n29), .B(n20), .C(n19), .D(n28), .Y(n92) );
  OAI22X1 U46 ( .A(n27), .B(n20), .C(n119), .D(n19), .Y(n91) );
  XNOR2X1 U47 ( .A(TX_CRC[1]), .B(n118), .Y(n119) );
  OAI22X1 U48 ( .A(n24), .B(n20), .C(n117), .D(n19), .Y(n90) );
  XOR2X1 U49 ( .A(n116), .B(n115), .Y(n117) );
  XNOR2X1 U50 ( .A(TX_CRC[0]), .B(n118), .Y(n116) );
  OAI22X1 U51 ( .A(n80), .B(n20), .C(n114), .D(n19), .Y(n89) );
  OAI22X1 U52 ( .A(n20), .B(n37), .C(n113), .D(n19), .Y(n88) );
  XNOR2X1 U53 ( .A(n112), .B(n111), .Y(n113) );
  OAI22X1 U54 ( .A(n20), .B(n35), .C(n110), .D(n121), .Y(n87) );
  OAI22X1 U55 ( .A(n20), .B(n33), .C(n109), .D(n121), .Y(n86) );
  XNOR2X1 U56 ( .A(n108), .B(n107), .Y(n109) );
  OAI22X1 U57 ( .A(n20), .B(n31), .C(n106), .D(n121), .Y(n85) );
  OAI22X1 U58 ( .A(n20), .B(n28), .C(n105), .D(n121), .Y(n84) );
  XOR2X1 U59 ( .A(n104), .B(n103), .Y(n105) );
  OAI22X1 U60 ( .A(n20), .B(n26), .C(n102), .D(n121), .Y(n83) );
  XOR2X1 U61 ( .A(n101), .B(n100), .Y(n102) );
  XOR2X1 U62 ( .A(n118), .B(n114), .Y(n101) );
  OAI22X1 U63 ( .A(n20), .B(n23), .C(n120), .D(n121), .Y(n82) );
  XOR2X1 U64 ( .A(n99), .B(n98), .Y(n120) );
  XOR2X1 U65 ( .A(n103), .B(n118), .Y(n98) );
  XNOR2X1 U66 ( .A(n25), .B(PRGA_OUT[7]), .Y(n118) );
  XNOR2X1 U67 ( .A(n24), .B(PRGA_OUT[0]), .Y(n103) );
  XOR2X1 U68 ( .A(n114), .B(n100), .Y(n99) );
  XOR2X1 U69 ( .A(n106), .B(n110), .Y(n100) );
  XNOR2X1 U70 ( .A(n107), .B(n112), .Y(n110) );
  XOR2X1 U71 ( .A(TX_CRC[12]), .B(PRGA_OUT[4]), .Y(n112) );
  XOR2X1 U72 ( .A(TX_CRC[11]), .B(PRGA_OUT[3]), .Y(n107) );
  XNOR2X1 U73 ( .A(n104), .B(n30), .Y(n106) );
  XOR2X1 U74 ( .A(TX_CRC[10]), .B(PRGA_OUT[2]), .Y(n108) );
  XNOR2X1 U75 ( .A(TX_CRC[9]), .B(PRGA_OUT[1]), .Y(n104) );
  XNOR2X1 U76 ( .A(n111), .B(n115), .Y(n114) );
  XNOR2X1 U77 ( .A(n79), .B(PRGA_OUT[6]), .Y(n115) );
  XOR2X1 U78 ( .A(TX_CRC[13]), .B(PRGA_OUT[5]), .Y(n111) );
  NAND3X1 U80 ( .A(PRGA_OPCODE[0]), .B(n81), .C(T_STROBE), .Y(n121) );
  DFFSR \current_crc_reg[6]  ( .D(n88), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[6]) );
  DFFSR \current_crc_reg[5]  ( .D(n87), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[5]) );
  DFFSR \current_crc_reg[4]  ( .D(n86), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[4]) );
  DFFSR \current_crc_reg[3]  ( .D(n85), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[3]) );
  DFFSR \current_crc_reg[2]  ( .D(n84), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[2]) );
  DFFSR \current_crc_reg[1]  ( .D(n83), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[1]) );
  DFFSR \current_crc_reg[0]  ( .D(n82), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[0]) );
  DFFSR \current_crc_reg[15]  ( .D(n97), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[15]) );
  DFFSR \current_crc_reg[14]  ( .D(n96), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[14]) );
  DFFSR \current_crc_reg[13]  ( .D(n95), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[13]) );
  DFFSR \current_crc_reg[12]  ( .D(n94), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[12]) );
  DFFSR \current_crc_reg[11]  ( .D(n93), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[11]) );
  DFFSR \current_crc_reg[10]  ( .D(n92), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[10]) );
  DFFSR \current_crc_reg[9]  ( .D(n91), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[9]) );
  DFFSR \current_crc_reg[8]  ( .D(n90), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[8]) );
  DFFSR \current_crc_reg[7]  ( .D(n89), .CLK(CLK), .R(n21), .S(1'b1), .Q(
        TX_CRC[7]) );
  AND2X2 U3 ( .A(n19), .B(n22), .Y(n1) );
  INVX2 U20 ( .A(n1), .Y(n20) );
  INVX2 U21 ( .A(RST), .Y(n21) );
  INVX2 U22 ( .A(n18), .Y(n19) );
  INVX2 U23 ( .A(n121), .Y(n18) );
  INVX2 U24 ( .A(EOP), .Y(n22) );
  INVX2 U25 ( .A(TX_CRC[0]), .Y(n23) );
  INVX2 U26 ( .A(TX_CRC[8]), .Y(n24) );
  INVX2 U27 ( .A(TX_CRC[15]), .Y(n25) );
  INVX2 U28 ( .A(TX_CRC[1]), .Y(n26) );
  INVX2 U29 ( .A(TX_CRC[9]), .Y(n27) );
  INVX2 U30 ( .A(TX_CRC[2]), .Y(n28) );
  INVX2 U31 ( .A(TX_CRC[10]), .Y(n29) );
  INVX2 U32 ( .A(n108), .Y(n30) );
  INVX2 U33 ( .A(TX_CRC[3]), .Y(n31) );
  INVX2 U34 ( .A(TX_CRC[11]), .Y(n32) );
  INVX2 U35 ( .A(TX_CRC[4]), .Y(n33) );
  INVX2 U36 ( .A(TX_CRC[12]), .Y(n34) );
  INVX2 U37 ( .A(TX_CRC[5]), .Y(n35) );
  INVX2 U38 ( .A(TX_CRC[13]), .Y(n36) );
  INVX2 U79 ( .A(TX_CRC[6]), .Y(n37) );
  INVX2 U81 ( .A(TX_CRC[14]), .Y(n79) );
  INVX2 U82 ( .A(TX_CRC[7]), .Y(n80) );
  INVX2 U83 ( .A(PRGA_OPCODE[1]), .Y(n81) );
endmodule


module tx_encode_0 ( clk, rst, SHIFT_ENABLE_E, d_encode, EOP, t_bitstuff, 
        dp_tx_out, dm_tx_out );
  input clk, rst, SHIFT_ENABLE_E, d_encode, EOP;
  output t_bitstuff, dp_tx_out, dm_tx_out;
  wire   DE_holdout, DE_holdout_BS, DE_holdout_last, DE_holdout_nxt, dm_tx_nxt,
         n16, n17, n21, n25, n28, n29, n30, n31, n34, n35, n42, n53, n54, n56,
         n57, n58, n59, n60, n63, n66, n68, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104;
  wire   [3:0] state;
  wire   [3:0] nextstate;

  DFFSR DE_holdout_reg ( .D(DE_holdout_nxt), .CLK(clk), .R(1'b1), .S(n16), .Q(
        DE_holdout) );
  DFFPOSX1 DE_holdout_last_reg ( .D(n68), .CLK(clk), .Q(DE_holdout_last) );
  DFFSR dp_tx_out_reg ( .D(DE_holdout_nxt), .CLK(clk), .R(1'b1), .S(n16), .Q(
        dp_tx_out) );
  AOI21X1 U3 ( .A(state[3]), .B(n104), .C(n30), .Y(nextstate[3]) );
  OAI21X1 U4 ( .A(n103), .B(n60), .C(n102), .Y(nextstate[2]) );
  AOI21X1 U5 ( .A(n101), .B(n17), .C(n34), .Y(n102) );
  NOR2X1 U7 ( .A(state[2]), .B(n59), .Y(n101) );
  AOI21X1 U8 ( .A(n35), .B(n59), .C(n99), .Y(n103) );
  OAI21X1 U9 ( .A(state[1]), .B(n100), .C(n98), .Y(nextstate[1]) );
  AOI21X1 U10 ( .A(state[1]), .B(n97), .C(n34), .Y(n98) );
  OAI21X1 U11 ( .A(state[0]), .B(n96), .C(n21), .Y(n97) );
  NAND3X1 U12 ( .A(SHIFT_ENABLE_E), .B(n35), .C(state[0]), .Y(n100) );
  OAI21X1 U14 ( .A(n58), .B(n21), .C(n95), .Y(nextstate[0]) );
  OAI21X1 U15 ( .A(n94), .B(n93), .C(SHIFT_ENABLE_E), .Y(n95) );
  OAI21X1 U16 ( .A(n31), .B(n92), .C(n91), .Y(n93) );
  NAND2X1 U17 ( .A(n90), .B(n42), .Y(n92) );
  NOR2X1 U18 ( .A(state[0]), .B(n96), .Y(n94) );
  NAND3X1 U19 ( .A(d_encode), .B(n89), .C(n88), .Y(n96) );
  XNOR2X1 U20 ( .A(n54), .B(n53), .Y(n88) );
  NOR2X1 U22 ( .A(n31), .B(SHIFT_ENABLE_E), .Y(n99) );
  OAI22X1 U23 ( .A(n16), .B(n54), .C(rst), .D(n53), .Y(n68) );
  OAI22X1 U26 ( .A(n25), .B(n63), .C(n53), .D(n87), .Y(n66) );
  NAND2X1 U28 ( .A(n34), .B(SHIFT_ENABLE_E), .Y(n87) );
  NAND3X1 U30 ( .A(n90), .B(n58), .C(n89), .Y(n91) );
  NOR2X1 U31 ( .A(state[3]), .B(n86), .Y(t_bitstuff) );
  OAI21X1 U32 ( .A(n57), .B(n56), .C(n85), .Y(dm_tx_nxt) );
  AOI22X1 U33 ( .A(n84), .B(n90), .C(n83), .D(n82), .Y(n85) );
  NOR2X1 U34 ( .A(n90), .B(n31), .Y(n83) );
  NOR2X1 U36 ( .A(EOP), .B(state[3]), .Y(n89) );
  NOR2X1 U37 ( .A(EOP), .B(n81), .Y(n84) );
  AOI22X1 U38 ( .A(state[0]), .B(n80), .C(n28), .D(n58), .Y(n81) );
  XNOR2X1 U40 ( .A(DE_holdout_BS), .B(n78), .Y(n80) );
  OAI21X1 U41 ( .A(n57), .B(n56), .C(n77), .Y(DE_holdout_nxt) );
  OAI21X1 U42 ( .A(n76), .B(n75), .C(n30), .Y(n77) );
  OAI21X1 U44 ( .A(n90), .B(n82), .C(n74), .Y(n75) );
  NAND3X1 U45 ( .A(n79), .B(n58), .C(n90), .Y(n74) );
  XOR2X1 U46 ( .A(DE_holdout), .B(SHIFT_ENABLE_E), .Y(n79) );
  XNOR2X1 U47 ( .A(n73), .B(n53), .Y(n82) );
  NAND2X1 U49 ( .A(SHIFT_ENABLE_E), .B(n42), .Y(n73) );
  OAI21X1 U51 ( .A(n86), .B(n72), .C(n71), .Y(n76) );
  AOI21X1 U52 ( .A(n70), .B(n29), .C(state[3]), .Y(n71) );
  NOR2X1 U54 ( .A(n63), .B(n86), .Y(n70) );
  NAND2X1 U55 ( .A(n78), .B(n63), .Y(n72) );
  NAND2X1 U57 ( .A(SHIFT_ENABLE_E), .B(d_encode), .Y(n78) );
  NAND2X1 U58 ( .A(state[0]), .B(n90), .Y(n86) );
  NOR2X1 U59 ( .A(n60), .B(n59), .Y(n90) );
  NAND3X1 U62 ( .A(n59), .B(n60), .C(n58), .Y(n104) );
  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(clk), .R(n16), .S(1'b1), .Q(
        state[3]) );
  DFFSR dm_tx_out_reg ( .D(dm_tx_nxt), .CLK(clk), .R(n16), .S(1'b1), .Q(
        dm_tx_out) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n16), .S(1'b1), .Q(
        state[0]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n16), .S(1'b1), .Q(
        state[1]) );
  DFFSR DE_holdout_BS_reg ( .D(n66), .CLK(clk), .R(n16), .S(1'b1), .Q(
        DE_holdout_BS) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n16), .S(1'b1), .Q(
        state[2]) );
  INVX2 U29 ( .A(rst), .Y(n16) );
  INVX2 U35 ( .A(n100), .Y(n17) );
  INVX2 U39 ( .A(n99), .Y(n21) );
  INVX2 U43 ( .A(n87), .Y(n25) );
  INVX2 U48 ( .A(n79), .Y(n28) );
  INVX2 U50 ( .A(n78), .Y(n29) );
  INVX2 U53 ( .A(EOP), .Y(n30) );
  INVX2 U56 ( .A(n89), .Y(n31) );
  INVX2 U60 ( .A(n91), .Y(n34) );
  INVX2 U61 ( .A(n96), .Y(n35) );
  INVX2 U63 ( .A(d_encode), .Y(n42) );
  INVX2 U64 ( .A(DE_holdout), .Y(n53) );
  INVX2 U65 ( .A(DE_holdout_last), .Y(n54) );
  INVX2 U66 ( .A(state[3]), .Y(n56) );
  INVX2 U68 ( .A(n104), .Y(n57) );
  INVX2 U69 ( .A(state[0]), .Y(n58) );
  INVX2 U70 ( .A(state[1]), .Y(n59) );
  INVX2 U71 ( .A(state[2]), .Y(n60) );
  INVX2 U72 ( .A(DE_holdout_BS), .Y(n63) );
endmodule


module tx_shiftreg_0 ( clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe, 
        send_data, d_encode );
  input [7:0] send_data;
  input clk, rst, SHIFT_ENABLE_R, t_bitstuff, t_strobe;
  output d_encode;
  wire   n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80;
  wire   [7:1] present_val;
  wire   [2:0] count;

  DFFSR \count_reg[0]  ( .D(n55), .CLK(clk), .R(1'b1), .S(n14), .Q(count[0])
         );
  DFFSR \count_reg[1]  ( .D(n57), .CLK(clk), .R(1'b1), .S(n14), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n56), .CLK(clk), .R(1'b1), .S(n14), .Q(count[2])
         );
  OAI21X1 U30 ( .A(n13), .B(n54), .C(n79), .Y(n65) );
  AOI22X1 U31 ( .A(send_data[0]), .B(n17), .C(present_val[1]), .D(n15), .Y(n79) );
  OAI21X1 U32 ( .A(n13), .B(n21), .C(n78), .Y(n64) );
  NAND2X1 U33 ( .A(send_data[7]), .B(n17), .Y(n78) );
  OAI21X1 U34 ( .A(n13), .B(n22), .C(n77), .Y(n63) );
  AOI22X1 U35 ( .A(send_data[6]), .B(n17), .C(present_val[7]), .D(n15), .Y(n77) );
  OAI21X1 U36 ( .A(n13), .B(n23), .C(n76), .Y(n62) );
  AOI22X1 U37 ( .A(send_data[5]), .B(n17), .C(present_val[6]), .D(n15), .Y(n76) );
  OAI21X1 U38 ( .A(n13), .B(n24), .C(n75), .Y(n61) );
  AOI22X1 U39 ( .A(send_data[4]), .B(n17), .C(present_val[5]), .D(n15), .Y(n75) );
  OAI21X1 U40 ( .A(n13), .B(n25), .C(n74), .Y(n60) );
  AOI22X1 U41 ( .A(send_data[3]), .B(n17), .C(present_val[4]), .D(n15), .Y(n74) );
  OAI21X1 U42 ( .A(n13), .B(n26), .C(n73), .Y(n59) );
  AOI22X1 U43 ( .A(send_data[2]), .B(n17), .C(present_val[3]), .D(n15), .Y(n73) );
  OAI21X1 U44 ( .A(n27), .B(n13), .C(n72), .Y(n58) );
  AOI22X1 U45 ( .A(send_data[1]), .B(n17), .C(present_val[2]), .D(n15), .Y(n72) );
  OAI21X1 U46 ( .A(n71), .B(n70), .C(n69), .Y(n57) );
  OAI21X1 U47 ( .A(n18), .B(n11), .C(count[1]), .Y(n69) );
  NAND2X1 U48 ( .A(count[0]), .B(n19), .Y(n70) );
  OAI21X1 U49 ( .A(n17), .B(n20), .C(n68), .Y(n56) );
  NAND3X1 U50 ( .A(count[1]), .B(count[0]), .C(n15), .Y(n68) );
  OAI22X1 U51 ( .A(n18), .B(n13), .C(count[0]), .D(n71), .Y(n55) );
  NAND2X1 U52 ( .A(n13), .B(n67), .Y(n71) );
  OAI21X1 U53 ( .A(t_bitstuff), .B(n16), .C(n67), .Y(n80) );
  NAND3X1 U54 ( .A(SHIFT_ENABLE_R), .B(count[0]), .C(n66), .Y(n67) );
  NOR2X1 U55 ( .A(n19), .B(n20), .Y(n66) );
  DFFSR \present_val_reg[7]  ( .D(n64), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[7]) );
  DFFSR \present_val_reg[1]  ( .D(n58), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[1]) );
  DFFSR \present_val_reg[6]  ( .D(n63), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[6]) );
  DFFSR \present_val_reg[5]  ( .D(n62), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[5]) );
  DFFSR \present_val_reg[4]  ( .D(n61), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[4]) );
  DFFSR \present_val_reg[3]  ( .D(n60), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[3]) );
  DFFSR \present_val_reg[2]  ( .D(n59), .CLK(clk), .R(n14), .S(1'b1), .Q(
        present_val[2]) );
  DFFSR \present_val_reg[0]  ( .D(n65), .CLK(clk), .R(n14), .S(1'b1), .Q(
        d_encode) );
  INVX4 U3 ( .A(n11), .Y(n13) );
  INVX2 U15 ( .A(rst), .Y(n14) );
  INVX2 U16 ( .A(n67), .Y(n17) );
  INVX2 U17 ( .A(n80), .Y(n11) );
  INVX2 U18 ( .A(n71), .Y(n15) );
  INVX2 U19 ( .A(SHIFT_ENABLE_R), .Y(n16) );
  INVX2 U20 ( .A(count[0]), .Y(n18) );
  INVX2 U21 ( .A(count[1]), .Y(n19) );
  INVX2 U22 ( .A(count[2]), .Y(n20) );
  INVX2 U23 ( .A(present_val[7]), .Y(n21) );
  INVX2 U24 ( .A(present_val[6]), .Y(n22) );
  INVX2 U25 ( .A(present_val[5]), .Y(n23) );
  INVX2 U26 ( .A(present_val[4]), .Y(n24) );
  INVX2 U27 ( .A(present_val[3]), .Y(n25) );
  INVX2 U28 ( .A(present_val[2]), .Y(n26) );
  INVX2 U29 ( .A(present_val[1]), .Y(n27) );
  INVX2 U56 ( .A(d_encode), .Y(n54) );
endmodule


module tx_tcu_0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module tx_tcu_0 ( clk, rst, p_ready, t_bitstuff, PRGA_OUT, prga_opcode, t_crc, 
        sending, EOP, next_byte, send_data, t_strobe );
  input [7:0] PRGA_OUT;
  input [1:0] prga_opcode;
  input [15:0] t_crc;
  output [7:0] send_data;
  input clk, rst, p_ready, t_bitstuff;
  output sending, EOP, next_byte, t_strobe;
  wire   N59, N60, N61, N62, N63, N64, N65, N84, N85, N86, N87, N88, N89, N90,
         N188, \r81/carry[6] , \r81/carry[5] , \r81/carry[4] , \r81/carry[3] ,
         \r81/carry[2] , \r81/carry[1] , \r81/B[0] , n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198;
  wire   [2:0] state;
  wire   [6:0] count;
  wire   [2:0] nextstate;
  wire   [7:0] flop_data;
  wire   [7:0] current_send_data;

  DFFPOSX1 \flop_data_reg[7]  ( .D(n152), .CLK(clk), .Q(flop_data[7]) );
  DFFPOSX1 \current_send_data_reg[7]  ( .D(n183), .CLK(clk), .Q(
        current_send_data[7]) );
  DFFPOSX1 \flop_data_reg[6]  ( .D(n153), .CLK(clk), .Q(flop_data[6]) );
  DFFPOSX1 \current_send_data_reg[6]  ( .D(n184), .CLK(clk), .Q(
        current_send_data[6]) );
  DFFPOSX1 \flop_data_reg[5]  ( .D(n154), .CLK(clk), .Q(flop_data[5]) );
  DFFPOSX1 \current_send_data_reg[5]  ( .D(n185), .CLK(clk), .Q(
        current_send_data[5]) );
  DFFPOSX1 \flop_data_reg[4]  ( .D(n155), .CLK(clk), .Q(flop_data[4]) );
  DFFPOSX1 \current_send_data_reg[4]  ( .D(n186), .CLK(clk), .Q(
        current_send_data[4]) );
  DFFPOSX1 \flop_data_reg[3]  ( .D(n156), .CLK(clk), .Q(flop_data[3]) );
  DFFPOSX1 \current_send_data_reg[3]  ( .D(n187), .CLK(clk), .Q(
        current_send_data[3]) );
  DFFPOSX1 \flop_data_reg[2]  ( .D(n157), .CLK(clk), .Q(flop_data[2]) );
  DFFPOSX1 \current_send_data_reg[2]  ( .D(n188), .CLK(clk), .Q(
        current_send_data[2]) );
  DFFPOSX1 \flop_data_reg[1]  ( .D(n174), .CLK(clk), .Q(flop_data[1]) );
  DFFPOSX1 \current_send_data_reg[1]  ( .D(n189), .CLK(clk), .Q(
        current_send_data[1]) );
  DFFPOSX1 \flop_data_reg[0]  ( .D(n175), .CLK(clk), .Q(flop_data[0]) );
  DFFPOSX1 \current_send_data_reg[0]  ( .D(n190), .CLK(clk), .Q(
        current_send_data[0]) );
  DFFPOSX1 \send_data_reg[7]  ( .D(n191), .CLK(clk), .Q(send_data[7]) );
  DFFPOSX1 \send_data_reg[6]  ( .D(n192), .CLK(clk), .Q(send_data[6]) );
  DFFPOSX1 \send_data_reg[5]  ( .D(n193), .CLK(clk), .Q(send_data[5]) );
  DFFPOSX1 \send_data_reg[4]  ( .D(n194), .CLK(clk), .Q(send_data[4]) );
  DFFPOSX1 \send_data_reg[3]  ( .D(n195), .CLK(clk), .Q(send_data[3]) );
  DFFPOSX1 \send_data_reg[2]  ( .D(n196), .CLK(clk), .Q(send_data[2]) );
  DFFPOSX1 \send_data_reg[1]  ( .D(n197), .CLK(clk), .Q(send_data[1]) );
  DFFPOSX1 \send_data_reg[0]  ( .D(n198), .CLK(clk), .Q(send_data[0]) );
  tx_tcu_0_DW01_inc_0 r80 ( .A({N188, count[5:0]}), .SUM({N65, N64, N63, N62, 
        N61, N60, N59}) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n15), .S(1'b1), .Q(
        state[2]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n15), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n15), .S(1'b1), .Q(
        state[0]) );
  DFFSR \count_reg[3]  ( .D(n180), .CLK(clk), .R(n15), .S(1'b1), .Q(count[3])
         );
  DFFSR \count_reg[2]  ( .D(n181), .CLK(clk), .R(n15), .S(1'b1), .Q(count[2])
         );
  DFFSR \count_reg[1]  ( .D(n182), .CLK(clk), .R(n15), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[0]  ( .D(n176), .CLK(clk), .R(n15), .S(1'b1), .Q(count[0])
         );
  DFFSR \count_reg[4]  ( .D(n179), .CLK(clk), .R(n15), .S(1'b1), .Q(count[4])
         );
  DFFSR \count_reg[5]  ( .D(n178), .CLK(clk), .R(n15), .S(1'b1), .Q(count[5])
         );
  DFFSR \count_reg[6]  ( .D(n177), .CLK(clk), .R(n15), .S(1'b1), .Q(N188) );
  INVX2 U13 ( .A(n12), .Y(n15) );
  BUFX2 U14 ( .A(rst), .Y(n13) );
  BUFX2 U15 ( .A(rst), .Y(n12) );
  BUFX2 U16 ( .A(rst), .Y(n14) );
  INVX2 U17 ( .A(N188), .Y(n11) );
  XOR2X1 U18 ( .A(N188), .B(\r81/carry[6] ), .Y(N90) );
  AND2X1 U19 ( .A(count[5]), .B(\r81/carry[5] ), .Y(\r81/carry[6] ) );
  XOR2X1 U20 ( .A(\r81/carry[5] ), .B(count[5]), .Y(N89) );
  AND2X1 U21 ( .A(count[4]), .B(\r81/carry[4] ), .Y(\r81/carry[5] ) );
  XOR2X1 U22 ( .A(\r81/carry[4] ), .B(count[4]), .Y(N88) );
  AND2X1 U23 ( .A(count[3]), .B(\r81/carry[3] ), .Y(\r81/carry[4] ) );
  XOR2X1 U24 ( .A(\r81/carry[3] ), .B(count[3]), .Y(N87) );
  AND2X1 U25 ( .A(count[2]), .B(\r81/carry[2] ), .Y(\r81/carry[3] ) );
  XOR2X1 U26 ( .A(\r81/carry[2] ), .B(count[2]), .Y(N86) );
  AND2X1 U27 ( .A(count[1]), .B(\r81/carry[1] ), .Y(\r81/carry[2] ) );
  XOR2X1 U28 ( .A(\r81/carry[1] ), .B(count[1]), .Y(N85) );
  AND2X1 U29 ( .A(count[0]), .B(\r81/B[0] ), .Y(\r81/carry[1] ) );
  XOR2X1 U30 ( .A(\r81/B[0] ), .B(count[0]), .Y(N84) );
  NOR2X1 U31 ( .A(n16), .B(n17), .Y(t_strobe) );
  NAND2X1 U32 ( .A(n18), .B(n19), .Y(n17) );
  NAND2X1 U33 ( .A(n11), .B(n20), .Y(n16) );
  OR2X1 U34 ( .A(n21), .B(n22), .Y(sending) );
  OAI21X1 U35 ( .A(N188), .B(n23), .C(n24), .Y(n22) );
  NAND3X1 U36 ( .A(n25), .B(n26), .C(n27), .Y(n21) );
  NAND3X1 U37 ( .A(n28), .B(n27), .C(n29), .Y(nextstate[2]) );
  AOI22X1 U38 ( .A(n30), .B(p_ready), .C(n31), .D(n32), .Y(n29) );
  NOR2X1 U39 ( .A(state[1]), .B(state[0]), .Y(n30) );
  NAND3X1 U40 ( .A(n33), .B(n34), .C(n35), .Y(nextstate[1]) );
  AOI22X1 U41 ( .A(n36), .B(n18), .C(n31), .D(n37), .Y(n35) );
  INVX1 U42 ( .A(n38), .Y(n36) );
  NAND3X1 U43 ( .A(n39), .B(n40), .C(p_ready), .Y(n33) );
  NAND3X1 U44 ( .A(n41), .B(n28), .C(n42), .Y(nextstate[0]) );
  AOI21X1 U45 ( .A(n18), .B(n38), .C(n43), .Y(n42) );
  OAI21X1 U46 ( .A(n44), .B(n27), .C(n45), .Y(n43) );
  NAND3X1 U47 ( .A(p_ready), .B(n37), .C(n31), .Y(n45) );
  AND2X1 U48 ( .A(n46), .B(n47), .Y(n31) );
  INVX1 U49 ( .A(n48), .Y(n44) );
  NAND3X1 U50 ( .A(n19), .B(n11), .C(count[0]), .Y(n38) );
  INVX1 U51 ( .A(n49), .Y(n28) );
  AND2X1 U52 ( .A(n26), .B(n25), .Y(n41) );
  OAI21X1 U53 ( .A(n50), .B(n51), .C(n52), .Y(next_byte) );
  MUX2X1 U54 ( .B(n53), .A(n54), .S(n55), .Y(n152) );
  INVX1 U55 ( .A(n56), .Y(n153) );
  MUX2X1 U56 ( .B(PRGA_OUT[6]), .A(flop_data[6]), .S(n55), .Y(n56) );
  INVX1 U57 ( .A(n57), .Y(n154) );
  MUX2X1 U58 ( .B(PRGA_OUT[5]), .A(flop_data[5]), .S(n55), .Y(n57) );
  INVX1 U59 ( .A(n58), .Y(n155) );
  MUX2X1 U60 ( .B(PRGA_OUT[4]), .A(flop_data[4]), .S(n55), .Y(n58) );
  INVX1 U61 ( .A(n59), .Y(n156) );
  MUX2X1 U62 ( .B(PRGA_OUT[3]), .A(flop_data[3]), .S(n55), .Y(n59) );
  INVX1 U63 ( .A(n60), .Y(n157) );
  MUX2X1 U64 ( .B(PRGA_OUT[2]), .A(flop_data[2]), .S(n55), .Y(n60) );
  INVX1 U65 ( .A(n61), .Y(n174) );
  MUX2X1 U66 ( .B(PRGA_OUT[1]), .A(flop_data[1]), .S(n55), .Y(n61) );
  INVX1 U67 ( .A(n62), .Y(n175) );
  MUX2X1 U68 ( .B(PRGA_OUT[0]), .A(flop_data[0]), .S(n55), .Y(n62) );
  NAND3X1 U69 ( .A(n63), .B(n23), .C(n64), .Y(n55) );
  AND2X1 U70 ( .A(n24), .B(n52), .Y(n64) );
  MUX2X1 U71 ( .B(n65), .A(n66), .S(n40), .Y(n52) );
  NOR2X1 U72 ( .A(p_ready), .B(n67), .Y(n66) );
  NOR2X1 U73 ( .A(n14), .B(n65), .Y(n63) );
  INVX1 U74 ( .A(t_bitstuff), .Y(\r81/B[0] ) );
  OAI21X1 U75 ( .A(n20), .B(n68), .C(n69), .Y(n176) );
  AOI22X1 U76 ( .A(N59), .B(n70), .C(N84), .D(n71), .Y(n69) );
  OAI21X1 U77 ( .A(n11), .B(n68), .C(n72), .Y(n177) );
  AOI22X1 U78 ( .A(N65), .B(n70), .C(N90), .D(n71), .Y(n72) );
  OAI21X1 U79 ( .A(n73), .B(n68), .C(n74), .Y(n178) );
  AOI22X1 U80 ( .A(N64), .B(n70), .C(N89), .D(n71), .Y(n74) );
  OAI21X1 U81 ( .A(n75), .B(n68), .C(n76), .Y(n179) );
  AOI22X1 U82 ( .A(N63), .B(n70), .C(N88), .D(n71), .Y(n76) );
  OAI21X1 U83 ( .A(n77), .B(n68), .C(n78), .Y(n180) );
  AOI22X1 U84 ( .A(N62), .B(n70), .C(N87), .D(n71), .Y(n78) );
  OAI21X1 U85 ( .A(n79), .B(n68), .C(n80), .Y(n181) );
  AOI22X1 U86 ( .A(N61), .B(n70), .C(N86), .D(n71), .Y(n80) );
  OAI21X1 U87 ( .A(n81), .B(n68), .C(n82), .Y(n182) );
  AOI22X1 U88 ( .A(N60), .B(n70), .C(N85), .D(n71), .Y(n82) );
  OAI21X1 U89 ( .A(n32), .B(n51), .C(n34), .Y(n71) );
  OR2X1 U90 ( .A(n25), .B(n48), .Y(n34) );
  NAND3X1 U91 ( .A(state[0]), .B(n83), .C(state[1]), .Y(n25) );
  INVX1 U92 ( .A(n37), .Y(n32) );
  NAND2X1 U93 ( .A(n48), .B(n50), .Y(n37) );
  AND2X1 U94 ( .A(prga_opcode[1]), .B(prga_opcode[0]), .Y(n50) );
  AND2X1 U95 ( .A(n68), .B(n84), .Y(n70) );
  OAI21X1 U96 ( .A(n48), .B(n27), .C(n85), .Y(n84) );
  NOR2X1 U97 ( .A(n18), .B(n49), .Y(n85) );
  NOR2X1 U98 ( .A(n86), .B(n87), .Y(n48) );
  NAND3X1 U99 ( .A(count[4]), .B(count[1]), .C(count[5]), .Y(n87) );
  NAND3X1 U100 ( .A(count[0]), .B(count[3]), .C(n88), .Y(n86) );
  NOR2X1 U101 ( .A(N188), .B(n79), .Y(n88) );
  NAND2X1 U102 ( .A(n18), .B(t_bitstuff), .Y(n68) );
  INVX1 U103 ( .A(count[1]), .Y(n81) );
  OAI21X1 U104 ( .A(n89), .B(n90), .C(n91), .Y(n183) );
  INVX1 U105 ( .A(current_send_data[7]), .Y(n90) );
  OAI21X1 U106 ( .A(n89), .B(n92), .C(n93), .Y(n184) );
  INVX1 U107 ( .A(current_send_data[6]), .Y(n92) );
  OAI21X1 U108 ( .A(n89), .B(n94), .C(n95), .Y(n185) );
  INVX1 U109 ( .A(current_send_data[5]), .Y(n94) );
  OAI21X1 U110 ( .A(n89), .B(n96), .C(n97), .Y(n186) );
  INVX1 U111 ( .A(current_send_data[4]), .Y(n96) );
  OAI21X1 U112 ( .A(n89), .B(n98), .C(n99), .Y(n187) );
  INVX1 U113 ( .A(current_send_data[3]), .Y(n98) );
  OAI21X1 U114 ( .A(n89), .B(n100), .C(n101), .Y(n188) );
  INVX1 U115 ( .A(current_send_data[2]), .Y(n100) );
  OAI21X1 U116 ( .A(n89), .B(n102), .C(n103), .Y(n189) );
  INVX1 U117 ( .A(current_send_data[1]), .Y(n102) );
  OAI21X1 U118 ( .A(n89), .B(n104), .C(n105), .Y(n190) );
  INVX1 U119 ( .A(current_send_data[0]), .Y(n104) );
  AOI21X1 U120 ( .A(state[0]), .B(state[1]), .C(n13), .Y(n89) );
  NAND2X1 U121 ( .A(n106), .B(n91), .Y(n191) );
  NOR2X1 U122 ( .A(n107), .B(n108), .Y(n91) );
  OAI21X1 U123 ( .A(n53), .B(n109), .C(n110), .Y(n108) );
  NAND2X1 U124 ( .A(t_crc[15]), .B(n111), .Y(n110) );
  INVX1 U125 ( .A(n112), .Y(n109) );
  INVX1 U126 ( .A(PRGA_OUT[7]), .Y(n53) );
  OAI22X1 U127 ( .A(n54), .B(n113), .C(n114), .D(n115), .Y(n107) );
  NAND2X1 U128 ( .A(n116), .B(state[0]), .Y(n115) );
  OAI21X1 U129 ( .A(N188), .B(t_crc[7]), .C(n15), .Y(n114) );
  INVX1 U130 ( .A(n117), .Y(n113) );
  INVX1 U131 ( .A(flop_data[7]), .Y(n54) );
  AOI22X1 U132 ( .A(n118), .B(current_send_data[7]), .C(send_data[7]), .D(n12), 
        .Y(n106) );
  NAND2X1 U133 ( .A(n119), .B(n93), .Y(n192) );
  AND2X1 U134 ( .A(n120), .B(n121), .Y(n93) );
  AOI22X1 U135 ( .A(t_crc[6]), .B(n122), .C(n117), .D(flop_data[6]), .Y(n121)
         );
  AOI22X1 U136 ( .A(t_crc[14]), .B(n111), .C(n112), .D(PRGA_OUT[6]), .Y(n120)
         );
  AOI22X1 U137 ( .A(n118), .B(current_send_data[6]), .C(send_data[6]), .D(n12), 
        .Y(n119) );
  NAND2X1 U138 ( .A(n123), .B(n95), .Y(n193) );
  AND2X1 U139 ( .A(n124), .B(n125), .Y(n95) );
  AOI22X1 U140 ( .A(t_crc[5]), .B(n122), .C(n117), .D(flop_data[5]), .Y(n125)
         );
  AOI22X1 U141 ( .A(t_crc[13]), .B(n111), .C(n112), .D(PRGA_OUT[5]), .Y(n124)
         );
  AOI22X1 U142 ( .A(n118), .B(current_send_data[5]), .C(send_data[5]), .D(n13), 
        .Y(n123) );
  NAND2X1 U143 ( .A(n126), .B(n97), .Y(n194) );
  AND2X1 U144 ( .A(n127), .B(n128), .Y(n97) );
  AOI22X1 U145 ( .A(t_crc[4]), .B(n122), .C(n117), .D(flop_data[4]), .Y(n128)
         );
  AOI22X1 U146 ( .A(t_crc[12]), .B(n111), .C(n112), .D(PRGA_OUT[4]), .Y(n127)
         );
  AOI22X1 U147 ( .A(n118), .B(current_send_data[4]), .C(send_data[4]), .D(n13), 
        .Y(n126) );
  NAND2X1 U148 ( .A(n129), .B(n99), .Y(n195) );
  AND2X1 U149 ( .A(n130), .B(n131), .Y(n99) );
  AOI22X1 U150 ( .A(t_crc[3]), .B(n122), .C(n117), .D(flop_data[3]), .Y(n131)
         );
  AOI22X1 U151 ( .A(t_crc[11]), .B(n111), .C(n112), .D(PRGA_OUT[3]), .Y(n130)
         );
  AOI22X1 U152 ( .A(n118), .B(current_send_data[3]), .C(send_data[3]), .D(n13), 
        .Y(n129) );
  NAND2X1 U153 ( .A(n132), .B(n101), .Y(n196) );
  AND2X1 U154 ( .A(n133), .B(n134), .Y(n101) );
  AOI22X1 U155 ( .A(t_crc[2]), .B(n122), .C(n117), .D(flop_data[2]), .Y(n134)
         );
  AOI22X1 U156 ( .A(t_crc[10]), .B(n111), .C(n112), .D(PRGA_OUT[2]), .Y(n133)
         );
  AOI22X1 U157 ( .A(n118), .B(current_send_data[2]), .C(send_data[2]), .D(n13), 
        .Y(n132) );
  NAND2X1 U158 ( .A(n135), .B(n103), .Y(n197) );
  AND2X1 U159 ( .A(n136), .B(n137), .Y(n103) );
  AOI22X1 U160 ( .A(t_crc[1]), .B(n122), .C(n117), .D(flop_data[1]), .Y(n137)
         );
  AOI22X1 U161 ( .A(t_crc[9]), .B(n111), .C(n112), .D(PRGA_OUT[1]), .Y(n136)
         );
  AOI22X1 U162 ( .A(n118), .B(current_send_data[1]), .C(send_data[1]), .D(n13), 
        .Y(n135) );
  NAND2X1 U163 ( .A(n138), .B(n105), .Y(n198) );
  AND2X1 U164 ( .A(n139), .B(n140), .Y(n105) );
  AOI22X1 U165 ( .A(t_crc[0]), .B(n122), .C(n117), .D(flop_data[0]), .Y(n140)
         );
  NOR2X1 U166 ( .A(n24), .B(n13), .Y(n117) );
  NOR2X1 U167 ( .A(n46), .B(n18), .Y(n24) );
  NOR2X1 U168 ( .A(n40), .B(n67), .Y(n18) );
  INVX1 U169 ( .A(n39), .Y(n67) );
  NOR2X1 U170 ( .A(state[1]), .B(state[2]), .Y(n39) );
  INVX1 U171 ( .A(n51), .Y(n46) );
  INVX1 U172 ( .A(n141), .Y(n122) );
  NAND3X1 U173 ( .A(n116), .B(state[0]), .C(n142), .Y(n141) );
  NOR2X1 U174 ( .A(n14), .B(N188), .Y(n142) );
  AOI22X1 U175 ( .A(t_crc[8]), .B(n111), .C(n112), .D(PRGA_OUT[0]), .Y(n139)
         );
  NOR2X1 U176 ( .A(n26), .B(n13), .Y(n112) );
  NAND2X1 U177 ( .A(n65), .B(n40), .Y(n26) );
  NOR2X1 U178 ( .A(n83), .B(n143), .Y(n65) );
  INVX1 U179 ( .A(state[1]), .Y(n143) );
  NOR2X1 U180 ( .A(n27), .B(n14), .Y(n111) );
  NAND2X1 U181 ( .A(n116), .B(n40), .Y(n27) );
  AOI22X1 U182 ( .A(n118), .B(current_send_data[0]), .C(send_data[0]), .D(n12), 
        .Y(n138) );
  INVX1 U183 ( .A(n144), .Y(n118) );
  NAND3X1 U184 ( .A(state[0]), .B(n15), .C(state[1]), .Y(n144) );
  OAI21X1 U185 ( .A(n51), .B(n47), .C(n145), .Y(EOP) );
  NAND3X1 U186 ( .A(N188), .B(n146), .C(n49), .Y(n145) );
  NOR2X1 U187 ( .A(n23), .B(n147), .Y(n49) );
  OAI21X1 U188 ( .A(n148), .B(n149), .C(state[0]), .Y(n147) );
  NAND3X1 U189 ( .A(count[2]), .B(N188), .C(count[3]), .Y(n149) );
  NAND3X1 U190 ( .A(n75), .B(n73), .C(n150), .Y(n148) );
  NOR2X1 U191 ( .A(count[1]), .B(count[0]), .Y(n150) );
  INVX1 U192 ( .A(count[5]), .Y(n73) );
  INVX1 U193 ( .A(count[4]), .Y(n75) );
  INVX1 U194 ( .A(n116), .Y(n23) );
  NOR2X1 U195 ( .A(n83), .B(state[1]), .Y(n116) );
  NAND3X1 U196 ( .A(n19), .B(n20), .C(N188), .Y(n47) );
  INVX1 U197 ( .A(count[0]), .Y(n20) );
  NOR2X1 U198 ( .A(n146), .B(count[1]), .Y(n19) );
  NAND3X1 U199 ( .A(n79), .B(n77), .C(n151), .Y(n146) );
  NOR2X1 U200 ( .A(count[5]), .B(count[4]), .Y(n151) );
  INVX1 U201 ( .A(count[3]), .Y(n77) );
  INVX1 U202 ( .A(count[2]), .Y(n79) );
  NAND3X1 U203 ( .A(n40), .B(n83), .C(state[1]), .Y(n51) );
  INVX1 U204 ( .A(state[2]), .Y(n83) );
  INVX1 U205 ( .A(state[0]), .Y(n40) );
endmodule


module tx_timer_0 ( CLK, RST, SENDING, SHIFT_ENABLE_R, SHIFT_ENABLE_E );
  input CLK, RST, SENDING;
  output SHIFT_ENABLE_R, SHIFT_ENABLE_E;
  wire   state, nxt_SHIFT_ENABLE_E, n7, n8, n9, n10, n11, n20, n21, n22, n23,
         n24, n25, n26, n27;
  wire   [3:0] count;
  wire   [3:0] nextcount;
  assign SHIFT_ENABLE_R = nxt_SHIFT_ENABLE_E;

  NOR2X1 U14 ( .A(n27), .B(n26), .Y(nextcount[3]) );
  XNOR2X1 U15 ( .A(count[3]), .B(n25), .Y(n27) );
  NOR2X1 U16 ( .A(n24), .B(n9), .Y(n25) );
  AOI21X1 U17 ( .A(n23), .B(state), .C(n11), .Y(nextcount[2]) );
  XNOR2X1 U18 ( .A(n24), .B(n9), .Y(n23) );
  NAND2X1 U19 ( .A(count[1]), .B(count[0]), .Y(n24) );
  NOR2X1 U20 ( .A(n22), .B(n26), .Y(nextcount[1]) );
  NAND3X1 U21 ( .A(SENDING), .B(n21), .C(state), .Y(n26) );
  XNOR2X1 U22 ( .A(count[0]), .B(count[1]), .Y(n22) );
  OAI21X1 U23 ( .A(count[0]), .B(n11), .C(state), .Y(nextcount[0]) );
  NOR2X1 U24 ( .A(n21), .B(n20), .Y(nxt_SHIFT_ENABLE_E) );
  NAND3X1 U25 ( .A(count[3]), .B(SENDING), .C(state), .Y(n20) );
  NAND3X1 U26 ( .A(n10), .B(n9), .C(n8), .Y(n21) );
  DFFSR state_reg ( .D(SENDING), .CLK(CLK), .R(n7), .S(1'b1), .Q(state) );
  DFFSR \count_reg[2]  ( .D(nextcount[2]), .CLK(CLK), .R(n7), .S(1'b1), .Q(
        count[2]) );
  DFFSR \count_reg[0]  ( .D(nextcount[0]), .CLK(CLK), .R(n7), .S(1'b1), .Q(
        count[0]) );
  DFFSR \count_reg[3]  ( .D(nextcount[3]), .CLK(CLK), .R(n7), .S(1'b1), .Q(
        count[3]) );
  DFFSR \count_reg[1]  ( .D(nextcount[1]), .CLK(CLK), .R(n7), .S(1'b1), .Q(
        count[1]) );
  DFFSR SHIFT_ENABLE_E_reg ( .D(nxt_SHIFT_ENABLE_E), .CLK(CLK), .R(n7), .S(
        1'b1), .Q(SHIFT_ENABLE_E) );
  INVX2 U9 ( .A(RST), .Y(n7) );
  INVX2 U10 ( .A(count[0]), .Y(n8) );
  INVX2 U11 ( .A(count[2]), .Y(n9) );
  INVX2 U12 ( .A(count[1]), .Y(n10) );
  INVX2 U13 ( .A(SENDING), .Y(n11) );
endmodule


module transmitter_block_0 ( PRGA_OUT, clk, p_ready, prga_opcode, rst, SENDING, 
        dm_tx_out, dp_tx_out, NEXT_BYTE );
  input [7:0] PRGA_OUT;
  input [1:0] prga_opcode;
  input clk, p_ready, rst;
  output SENDING, dm_tx_out, dp_tx_out, NEXT_BYTE;
  wire   t_strobe, EOP, SHIFT_ENABLE_E, d_encode, t_bitstuff, SHIFT_ENABLE_R;
  wire   [15:0] TX_CRC;
  wire   [7:0] send_data;

  tx_CRC_CALC_0 U_1 ( .CLK(clk), .RST(rst), .EOP(EOP), .T_STROBE(t_strobe), 
        .PRGA_OPCODE(prga_opcode), .PRGA_OUT(PRGA_OUT), .TX_CRC(TX_CRC) );
  tx_encode_0 U_0 ( .clk(clk), .rst(rst), .SHIFT_ENABLE_E(SHIFT_ENABLE_E), 
        .d_encode(d_encode), .EOP(EOP), .t_bitstuff(t_bitstuff), .dp_tx_out(
        dp_tx_out), .dm_tx_out(dm_tx_out) );
  tx_shiftreg_0 U_2 ( .clk(clk), .rst(rst), .SHIFT_ENABLE_R(SHIFT_ENABLE_R), 
        .t_bitstuff(t_bitstuff), .t_strobe(t_strobe), .send_data(send_data), 
        .d_encode(d_encode) );
  tx_tcu_0 U_3 ( .clk(clk), .rst(rst), .p_ready(p_ready), .t_bitstuff(
        t_bitstuff), .PRGA_OUT(PRGA_OUT), .prga_opcode(prga_opcode), .t_crc(
        TX_CRC), .sending(SENDING), .EOP(EOP), .next_byte(NEXT_BYTE), 
        .send_data(send_data), .t_strobe(t_strobe) );
  tx_timer_0 U_4 ( .CLK(clk), .RST(rst), .SENDING(SENDING), .SHIFT_ENABLE_R(
        SHIFT_ENABLE_R), .SHIFT_ENABLE_E(SHIFT_ENABLE_E) );
endmodule


module RMEDT_REWIRE_0 ( CLK, DM1_RX, DP1_RX, RST, SERIAL_IN, DATA_IN, BS_ERROR, 
        CRC_ERROR, EMPTY, FULL, KEY_ERROR, PROG_ERROR, PARITY_ERROR, RBUF_FULL, 
        R_ERROR, SENDING, dm_tx_out, dp_tx_out, W_ENABLE_R, R_ENABLE, DATA, 
        ADDR );
  input [7:0] DATA_IN;
  output [7:0] DATA;
  output [7:0] ADDR;
  input CLK, DM1_RX, DP1_RX, RST, SERIAL_IN;
  output BS_ERROR, CRC_ERROR, EMPTY, FULL, KEY_ERROR, PROG_ERROR, PARITY_ERROR,
         RBUF_FULL, R_ERROR, SENDING, dm_tx_out, dp_tx_out, W_ENABLE_R,
         R_ENABLE;
  wire   B_READY, PDATA_READY, EOP_external, NEXT_BYTE, W_ENABLE, n1, n2;
  wire   [7:0] PRGA_IN;
  wire   [1:0] PRGA_OPCODE;
  wire   [7:0] PROCESSED_DATA;
  wire   [7:0] RCV_DATA;
  wire   [1:0] OPCODE;

  EDBlock_0 U_0 ( .BYTE(PRGA_IN), .BYTE_READY(B_READY), .CLK(CLK), .OPCODE(
        PRGA_OPCODE), .RST(n1), .SERIAL_IN(SERIAL_IN), .DATA_IN(DATA_IN), 
        .KEY_ERROR(KEY_ERROR), .PARITY_ERROR(PARITY_ERROR), .PDATA_READY(
        PDATA_READY), .PROCESSED_DATA(PROCESSED_DATA), .PROG_ERROR(PROG_ERROR), 
        .RBUF_FULL(RBUF_FULL), .W_ENABLE(W_ENABLE_R), .R_ENABLE(R_ENABLE), 
        .DATA(DATA), .ADDR(ADDR) );
  memoryblock_0 U_1 ( .CLK(CLK), .NEXT_BYTE(NEXT_BYTE), .RCV_DATA(RCV_DATA), 
        .RCV_OPCODE(OPCODE), .RST(n1), .W_ENABLE(W_ENABLE), .EOP(EOP_external), 
        .EMPTY(EMPTY), .FULL(FULL), .B_READY(B_READY), .PRGA_IN(PRGA_IN), 
        .PRGA_OPCODE(PRGA_OPCODE) );
  receiver_block_rewire_0 U_2 ( .CLK(CLK), .DM1_RX(DM1_RX), .DP1_RX(DP1_RX), 
        .RST(n1), .BS_ERROR(BS_ERROR), .CRC_ERROR(CRC_ERROR), .EOP_external(
        EOP_external), .OPCODE(OPCODE), .RCV_DATA(RCV_DATA), .R_ERROR(R_ERROR), 
        .W_ENABLE(W_ENABLE) );
  transmitter_block_0 U_3 ( .PRGA_OUT(PROCESSED_DATA), .clk(CLK), .p_ready(
        PDATA_READY), .prga_opcode(PRGA_OPCODE), .rst(n1), .SENDING(SENDING), 
        .dm_tx_out(dm_tx_out), .dp_tx_out(dp_tx_out), .NEXT_BYTE(NEXT_BYTE) );
  INVX2 U1 ( .A(n2), .Y(n1) );
  INVX2 U2 ( .A(RST), .Y(n2) );
endmodule


module rmedt_square_t ( CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN, DATA_IN_H, 
        DATA_IN_S, BSE_H, BSE_S, CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, 
        EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, 
        c_parity_error, c_prog_error, host_is_sending, slave_is_sending, 
        W_ENABLE_H, W_ENABLE_S, R_ENABLE_H, R_ENABLE_S, DATA_H, DATA_S, ADDR_H, 
        ADDR_S );
  input [7:0] DATA_IN_H;
  input [7:0] DATA_IN_S;
  output [7:0] DATA_H;
  output [7:0] DATA_S;
  output [7:0] ADDR_H;
  output [7:0] ADDR_S;
  input CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN;
  output BSE_H, BSE_S, CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, EMPTY_H,
         EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, c_parity_error,
         c_prog_error, host_is_sending, slave_is_sending, W_ENABLE_H,
         W_ENABLE_S, R_ENABLE_H, R_ENABLE_S;
  wire   KEY_ERROR, KEY_ERROR1, PARITY_ERROR, PARITY_ERROR1, PROG_ERROR,
         PROG_ERROR1;

  OR2X2 U1 ( .A(PROG_ERROR), .B(PROG_ERROR1), .Y(c_prog_error) );
  OR2X2 U2 ( .A(PARITY_ERROR), .B(PARITY_ERROR1), .Y(c_parity_error) );
  OR2X2 U3 ( .A(KEY_ERROR), .B(KEY_ERROR1), .Y(c_key_error) );
  RMEDT_REWIRE_1 U_0 ( .CLK(CLK), .DM1_RX(DMRH), .DP1_RX(DPRH), .RST(RST), 
        .SERIAL_IN(SERIAL_IN), .DATA_IN(DATA_IN_H), .BS_ERROR(BSE_H), 
        .CRC_ERROR(CRCE_H), .EMPTY(EMPTY_H), .FULL(FULL_H), .KEY_ERROR(
        KEY_ERROR), .PROG_ERROR(PROG_ERROR), .PARITY_ERROR(PARITY_ERROR), 
        .R_ERROR(RE_H), .SENDING(host_is_sending), .dm_tx_out(DMTS), 
        .dp_tx_out(DPTS), .W_ENABLE_R(W_ENABLE_H), .R_ENABLE(R_ENABLE_H), 
        .DATA(DATA_H), .ADDR(ADDR_H) );
  RMEDT_REWIRE_0 U_1 ( .CLK(CLK), .DM1_RX(DMRS), .DP1_RX(DPRS), .RST(RST), 
        .SERIAL_IN(SERIAL_IN), .DATA_IN(DATA_IN_S), .BS_ERROR(BSE_S), 
        .CRC_ERROR(CRCE_S), .EMPTY(EMPTY_S), .FULL(FULL_S), .KEY_ERROR(
        KEY_ERROR1), .PROG_ERROR(PROG_ERROR1), .PARITY_ERROR(PARITY_ERROR1), 
        .R_ERROR(RE_S), .SENDING(slave_is_sending), .dm_tx_out(DMTH), 
        .dp_tx_out(DPTH), .W_ENABLE_R(W_ENABLE_S), .R_ENABLE(R_ENABLE_S), 
        .DATA(DATA_S), .ADDR(ADDR_S) );
endmodule

module  rmedt_square ( CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN, BSE_H, BSE_S, 
	CRCE_H, CRCE_S, DMTH, DMTS, DPTH, DPTS, DPHS, DMHS, DPSS, DMSS, EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, 
	RE_S, c_key_error, c_parity_error, c_prog_error, host_is_sending, slave_is_sending );

input   CLK, DMRH, DMRS, DPRH, DPRS, RST, SERIAL_IN;
output  BSE_H, BSE_S, CRCE_H, CRCE_S, EMPTY_H, EMPTY_S, FULL_H, FULL_S, RE_H, RE_S, c_key_error, c_parity_error, c_prog_error, DMTH, DMTS, DPTH, DPTS, slave_is_sending, host_is_sending;
inout   DPHS, DMHS, DPSS, DMSS;
wire	nCLK, nDMRH, nDMRS, nDPRH, nDPRS, nRST, nSERIAL_IN, nBSE_H, nBSE_S, nCRCE_H, nCRCE_S, nDMTH, nDMTS, nDPTH, nDPTS, nEMPTY_H, nEMPTY_S, nFULL_H, nFULL_S, nRE_H, nRE_S, nc_key_error, nc_parity_error, nc_prog_error, nhost_is_sending, nslave_is_sending;

        rmedt_square_t I0 ( .CLK(nCLK), .DMRH(nDMRH), .DMRS(nDMRS), .DPRH(nDPRH), 
	.DPRS(nDPRS), .RST(nRST), .SERIAL_IN(nSERIAL_IN), .BSE_H(nBSE_H), .BSE_S(nBSE_S), 
	.CRCE_H(nCRCE_H), .CRCE_S(nCRCE_S), .DMTH(nDMTH), .DMTS(nDMTS), 
	.DPTH(nDPTH), .DPTS(nDPTS), .EMPTY_H(nEMPTY_H), .EMPTY_S(nSERIAL_IN), 
	.FULL_H(nFULL_H), .FULL_S(nFULL_S), .RE_H(nRE_H), .RE_S(nRE_S), 
	.c_key_error(nc_key_error), .c_parity_error(nc_parity_error), .c_prog_error(nc_prog_error), .host_is_sending(nhost_is_sending), 
	.slave_is_sending(nslave_is_sending));

PADVDD U1 (  );
PADGND U2 (  );
PADINC U3 ( .DI(nCLK), .YPAD(CLK) );
PADINC U8 ( .DI(nRST), .YPAD(RST) );
PADINC U9 ( .DI(nSERIAL_IN), .YPAD(SERIAL_IN) );
PADINOUT UIO1 ( .DI(nDPRH), .DO(nDPTH), .OEN(nslave_is_sending), .YPAD(DPHS));
PADINOUT UIO2 ( .DI(nDMRH), .DO(nDMTH), .OEN(nslave_is_sending), .YPAD(DMHS));
PADINOUT UIO3 ( .DI(nDPRS), .DO(nDPTS), .OEN(nhost_is_sending), .YPAD(DPSS));
PADINOUT UIO4 ( .DI(nDMRS), .DO(nDMTS), .OEN(nhost_is_sending), .YPAD(DMSS));
PADOUT UOUT1 ( .DO(BSE_H), .YPAD(nBSE_H) );
PADOUT UOUT2 ( .DO(BSE_S), .YPAD(nBSE_S) );
PADOUT UOUT3 ( .DO(CRCE_H), .YPAD(nCRCE_H) );
PADOUT UOUT4 ( .DO(CRCE_S), .YPAD(nCRCE_S) );
PADOUT UOUT5 ( .DO(EMPTY_H), .YPAD(nEMPTY_H) );
PADOUT UOUT6 ( .DO(EMPTY_S), .YPAD(nEMPTY_S) );
PADOUT UOUT7 ( .DO(FULL_H), .YPAD(nFULL_H) );
PADOUT UOUT8 ( .DO(FULL_S), .YPAD(nFULL_S) );
PADOUT UOUT9 ( .DO(RE_H), .YPAD(nRE_H) );
PADOUT UOUT10 ( .DO(RE_S), .YPAD(nRE_S) );
PADOUT UOUT11 ( .DO(c_key_error), .YPAD(nc_key_error) );
PADOUT UOUT12 ( .DO(c_parity_error), .YPAD(nc_parity_error) );
PADOUT UOUT13 ( .DO(c_prog_error), .YPAD(nc_prog_error) );

endmodule

